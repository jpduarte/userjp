*script to generate hspice simulation using cmdp, Juan Duarte 
*Date: 07/31/2016, time: 19:06:43

.option abstol=1e-6 reltol=1e-6 post ingold 
.option ABSV=1e-2 
.option measform=1 
.temp 27 

.hdl "/users/jpduarte/research/userjp/ncfet/models/fecm.va" 
.include "/users/jpduarte/research/userjp/ncfet/modelcards/modelcard_fe.fe" 

.PARAM Vp_value = 0 
.PARAM Vn_value = 0 
.PARAM r_value = 1 
.PARAM a0_value = -1 
.PARAM b0_value = 0.1 

Vp Vp 0.0 dc = Vp_value 
Vn Vn 0.0 dc = Vn_value 

X1 Vp Vn nmos1 r = 'r_value' a0 = 'a0_value' b0 = 'b0_value'

.DATA datadc Vp_value Vn_value r_value a0_value b0_value 
0.0 0 1 -1 0.1 
0.204081632653 0 1 -1 0.1 
0.408163265306 0 1 -1 0.1 
0.612244897959 0 1 -1 0.1 
0.816326530612 0 1 -1 0.1 
1.02040816327 0 1 -1 0.1 
1.22448979592 0 1 -1 0.1 
1.42857142857 0 1 -1 0.1 
1.63265306122 0 1 -1 0.1 
1.83673469388 0 1 -1 0.1 
2.04081632653 0 1 -1 0.1 
2.24489795918 0 1 -1 0.1 
2.44897959184 0 1 -1 0.1 
2.65306122449 0 1 -1 0.1 
2.85714285714 0 1 -1 0.1 
3.0612244898 0 1 -1 0.1 
3.26530612245 0 1 -1 0.1 
3.4693877551 0 1 -1 0.1 
3.67346938776 0 1 -1 0.1 
3.87755102041 0 1 -1 0.1 
4.08163265306 0 1 -1 0.1 
4.28571428571 0 1 -1 0.1 
4.48979591837 0 1 -1 0.1 
4.69387755102 0 1 -1 0.1 
4.89795918367 0 1 -1 0.1 
5.10204081633 0 1 -1 0.1 
5.30612244898 0 1 -1 0.1 
5.51020408163 0 1 -1 0.1 
5.71428571429 0 1 -1 0.1 
5.91836734694 0 1 -1 0.1 
6.12244897959 0 1 -1 0.1 
6.32653061224 0 1 -1 0.1 
6.5306122449 0 1 -1 0.1 
6.73469387755 0 1 -1 0.1 
6.9387755102 0 1 -1 0.1 
7.14285714286 0 1 -1 0.1 
7.34693877551 0 1 -1 0.1 
7.55102040816 0 1 -1 0.1 
7.75510204082 0 1 -1 0.1 
7.95918367347 0 1 -1 0.1 
8.16326530612 0 1 -1 0.1 
8.36734693878 0 1 -1 0.1 
8.57142857143 0 1 -1 0.1 
8.77551020408 0 1 -1 0.1 
8.97959183673 0 1 -1 0.1 
9.18367346939 0 1 -1 0.1 
9.38775510204 0 1 -1 0.1 
9.59183673469 0 1 -1 0.1 
9.79591836735 0 1 -1 0.1 
10.0 0 1 -1 0.1 
10.0 0 1 -1 0.1 
9.59183673469 0 1 -1 0.1 
9.18367346939 0 1 -1 0.1 
8.77551020408 0 1 -1 0.1 
8.36734693878 0 1 -1 0.1 
7.95918367347 0 1 -1 0.1 
7.55102040816 0 1 -1 0.1 
7.14285714286 0 1 -1 0.1 
6.73469387755 0 1 -1 0.1 
6.32653061224 0 1 -1 0.1 
5.91836734694 0 1 -1 0.1 
5.51020408163 0 1 -1 0.1 
5.10204081633 0 1 -1 0.1 
4.69387755102 0 1 -1 0.1 
4.28571428571 0 1 -1 0.1 
3.87755102041 0 1 -1 0.1 
3.4693877551 0 1 -1 0.1 
3.0612244898 0 1 -1 0.1 
2.65306122449 0 1 -1 0.1 
2.24489795918 0 1 -1 0.1 
1.83673469388 0 1 -1 0.1 
1.42857142857 0 1 -1 0.1 
1.02040816327 0 1 -1 0.1 
0.612244897959 0 1 -1 0.1 
0.204081632653 0 1 -1 0.1 
-0.204081632653 0 1 -1 0.1 
-0.612244897959 0 1 -1 0.1 
-1.02040816327 0 1 -1 0.1 
-1.42857142857 0 1 -1 0.1 
-1.83673469388 0 1 -1 0.1 
-2.24489795918 0 1 -1 0.1 
-2.65306122449 0 1 -1 0.1 
-3.0612244898 0 1 -1 0.1 
-3.4693877551 0 1 -1 0.1 
-3.87755102041 0 1 -1 0.1 
-4.28571428571 0 1 -1 0.1 
-4.69387755102 0 1 -1 0.1 
-5.10204081633 0 1 -1 0.1 
-5.51020408163 0 1 -1 0.1 
-5.91836734694 0 1 -1 0.1 
-6.32653061224 0 1 -1 0.1 
-6.73469387755 0 1 -1 0.1 
-7.14285714286 0 1 -1 0.1 
-7.55102040816 0 1 -1 0.1 
-7.95918367347 0 1 -1 0.1 
-8.36734693878 0 1 -1 0.1 
-8.77551020408 0 1 -1 0.1 
-9.18367346939 0 1 -1 0.1 
-9.59183673469 0 1 -1 0.1 
-10.0 0 1 -1 0.1 
-10.0 0 1 -1 0.1 
-9.59183673469 0 1 -1 0.1 
-9.18367346939 0 1 -1 0.1 
-8.77551020408 0 1 -1 0.1 
-8.36734693878 0 1 -1 0.1 
-7.95918367347 0 1 -1 0.1 
-7.55102040816 0 1 -1 0.1 
-7.14285714286 0 1 -1 0.1 
-6.73469387755 0 1 -1 0.1 
-6.32653061224 0 1 -1 0.1 
-5.91836734694 0 1 -1 0.1 
-5.51020408163 0 1 -1 0.1 
-5.10204081633 0 1 -1 0.1 
-4.69387755102 0 1 -1 0.1 
-4.28571428571 0 1 -1 0.1 
-3.87755102041 0 1 -1 0.1 
-3.4693877551 0 1 -1 0.1 
-3.0612244898 0 1 -1 0.1 
-2.65306122449 0 1 -1 0.1 
-2.24489795918 0 1 -1 0.1 
-1.83673469388 0 1 -1 0.1 
-1.42857142857 0 1 -1 0.1 
-1.02040816327 0 1 -1 0.1 
-0.612244897959 0 1 -1 0.1 
-0.204081632653 0 1 -1 0.1 
0.204081632653 0 1 -1 0.1 
0.612244897959 0 1 -1 0.1 
1.02040816327 0 1 -1 0.1 
1.42857142857 0 1 -1 0.1 
1.83673469388 0 1 -1 0.1 
2.24489795918 0 1 -1 0.1 
2.65306122449 0 1 -1 0.1 
3.0612244898 0 1 -1 0.1 
3.4693877551 0 1 -1 0.1 
3.87755102041 0 1 -1 0.1 
4.28571428571 0 1 -1 0.1 
4.69387755102 0 1 -1 0.1 
5.10204081633 0 1 -1 0.1 
5.51020408163 0 1 -1 0.1 
5.91836734694 0 1 -1 0.1 
6.32653061224 0 1 -1 0.1 
6.73469387755 0 1 -1 0.1 
7.14285714286 0 1 -1 0.1 
7.55102040816 0 1 -1 0.1 
7.95918367347 0 1 -1 0.1 
8.36734693878 0 1 -1 0.1 
8.77551020408 0 1 -1 0.1 
9.18367346939 0 1 -1 0.1 
9.59183673469 0 1 -1 0.1 
10.0 0 1 -1 0.1 
.ENDDATA 
.dc sweep DATA = datadc 
.print dc X1:qfe X1:vfe 
.end