*script to generate hspice simulation using cmdp, Juan Duarte 
*Date: 02/08/2016, time: 19:43:23

.option abstol=1e-6 reltol=1e-6 post ingold 
.option measform=1 
.temp 27 

.hdl "/users/jpduarte/research/BSIMIMG/code/bsimimg.va" 
.include "/users/jpduarte/research/userjp/project4/modelcards/modelcardsimple.nmos" 

.PARAM Vd_value = 0 
.PARAM Vgf_value = 0 
.PARAM Vs_value = 0 
.PARAM Vgb_value = 0 
.PARAM L_value = 1e-06 

Vd Vd 0.0 dc = Vd_value 
Vgf Vgf 0.0 dc = Vgf_value 
Vs Vs 0.0 dc = Vs_value 
Vgb Vgb 0.0 dc = Vgb_value 

X1 Vd Vgf Vs Vgb nmos1 L = 'L_value'

.DATA datadc Vd_value Vgf_value Vs_value Vgb_value L_value 
0.05 0.0 0 -3.0 1e-06 
3.0 0.0 0 -3.0 1e-06 
0.05 0.001 0 -3.0 1e-06 
3.0 0.001 0 -3.0 1e-06 
0.05 0.002 0 -3.0 1e-06 
3.0 0.002 0 -3.0 1e-06 
0.05 0.003 0 -3.0 1e-06 
3.0 0.003 0 -3.0 1e-06 
0.05 0.004 0 -3.0 1e-06 
3.0 0.004 0 -3.0 1e-06 
0.05 0.005 0 -3.0 1e-06 
3.0 0.005 0 -3.0 1e-06 
0.05 0.006 0 -3.0 1e-06 
3.0 0.006 0 -3.0 1e-06 
0.05 0.007 0 -3.0 1e-06 
3.0 0.007 0 -3.0 1e-06 
0.05 0.008 0 -3.0 1e-06 
3.0 0.008 0 -3.0 1e-06 
0.05 0.009 0 -3.0 1e-06 
3.0 0.009 0 -3.0 1e-06 
0.05 0.01 0 -3.0 1e-06 
3.0 0.01 0 -3.0 1e-06 
0.05 0.011 0 -3.0 1e-06 
3.0 0.011 0 -3.0 1e-06 
0.05 0.012 0 -3.0 1e-06 
3.0 0.012 0 -3.0 1e-06 
0.05 0.013 0 -3.0 1e-06 
3.0 0.013 0 -3.0 1e-06 
0.05 0.014 0 -3.0 1e-06 
3.0 0.014 0 -3.0 1e-06 
0.05 0.015 0 -3.0 1e-06 
3.0 0.015 0 -3.0 1e-06 
0.05 0.016 0 -3.0 1e-06 
3.0 0.016 0 -3.0 1e-06 
0.05 0.017 0 -3.0 1e-06 
3.0 0.017 0 -3.0 1e-06 
0.05 0.018 0 -3.0 1e-06 
3.0 0.018 0 -3.0 1e-06 
0.05 0.019 0 -3.0 1e-06 
3.0 0.019 0 -3.0 1e-06 
0.05 0.02 0 -3.0 1e-06 
3.0 0.02 0 -3.0 1e-06 
0.05 0.021 0 -3.0 1e-06 
3.0 0.021 0 -3.0 1e-06 
0.05 0.022 0 -3.0 1e-06 
3.0 0.022 0 -3.0 1e-06 
0.05 0.023 0 -3.0 1e-06 
3.0 0.023 0 -3.0 1e-06 
0.05 0.024 0 -3.0 1e-06 
3.0 0.024 0 -3.0 1e-06 
0.05 0.025 0 -3.0 1e-06 
3.0 0.025 0 -3.0 1e-06 
0.05 0.026 0 -3.0 1e-06 
3.0 0.026 0 -3.0 1e-06 
0.05 0.027 0 -3.0 1e-06 
3.0 0.027 0 -3.0 1e-06 
0.05 0.028 0 -3.0 1e-06 
3.0 0.028 0 -3.0 1e-06 
0.05 0.029 0 -3.0 1e-06 
3.0 0.029 0 -3.0 1e-06 
0.05 0.03 0 -3.0 1e-06 
3.0 0.03 0 -3.0 1e-06 
0.05 0.031 0 -3.0 1e-06 
3.0 0.031 0 -3.0 1e-06 
0.05 0.032 0 -3.0 1e-06 
3.0 0.032 0 -3.0 1e-06 
0.05 0.033 0 -3.0 1e-06 
3.0 0.033 0 -3.0 1e-06 
0.05 0.034 0 -3.0 1e-06 
3.0 0.034 0 -3.0 1e-06 
0.05 0.035 0 -3.0 1e-06 
3.0 0.035 0 -3.0 1e-06 
0.05 0.036 0 -3.0 1e-06 
3.0 0.036 0 -3.0 1e-06 
0.05 0.037 0 -3.0 1e-06 
3.0 0.037 0 -3.0 1e-06 
0.05 0.038 0 -3.0 1e-06 
3.0 0.038 0 -3.0 1e-06 
0.05 0.039 0 -3.0 1e-06 
3.0 0.039 0 -3.0 1e-06 
0.05 0.04 0 -3.0 1e-06 
3.0 0.04 0 -3.0 1e-06 
0.05 0.041 0 -3.0 1e-06 
3.0 0.041 0 -3.0 1e-06 
0.05 0.042 0 -3.0 1e-06 
3.0 0.042 0 -3.0 1e-06 
0.05 0.043 0 -3.0 1e-06 
3.0 0.043 0 -3.0 1e-06 
0.05 0.044 0 -3.0 1e-06 
3.0 0.044 0 -3.0 1e-06 
0.05 0.045 0 -3.0 1e-06 
3.0 0.045 0 -3.0 1e-06 
0.05 0.046 0 -3.0 1e-06 
3.0 0.046 0 -3.0 1e-06 
0.05 0.047 0 -3.0 1e-06 
3.0 0.047 0 -3.0 1e-06 
0.05 0.048 0 -3.0 1e-06 
3.0 0.048 0 -3.0 1e-06 
0.05 0.049 0 -3.0 1e-06 
3.0 0.049 0 -3.0 1e-06 
0.05 0.05 0 -3.0 1e-06 
3.0 0.05 0 -3.0 1e-06 
0.05 0.051 0 -3.0 1e-06 
3.0 0.051 0 -3.0 1e-06 
0.05 0.052 0 -3.0 1e-06 
3.0 0.052 0 -3.0 1e-06 
0.05 0.053 0 -3.0 1e-06 
3.0 0.053 0 -3.0 1e-06 
0.05 0.054 0 -3.0 1e-06 
3.0 0.054 0 -3.0 1e-06 
0.05 0.055 0 -3.0 1e-06 
3.0 0.055 0 -3.0 1e-06 
0.05 0.056 0 -3.0 1e-06 
3.0 0.056 0 -3.0 1e-06 
0.05 0.057 0 -3.0 1e-06 
3.0 0.057 0 -3.0 1e-06 
0.05 0.058 0 -3.0 1e-06 
3.0 0.058 0 -3.0 1e-06 
0.05 0.059 0 -3.0 1e-06 
3.0 0.059 0 -3.0 1e-06 
0.05 0.06 0 -3.0 1e-06 
3.0 0.06 0 -3.0 1e-06 
0.05 0.061 0 -3.0 1e-06 
3.0 0.061 0 -3.0 1e-06 
0.05 0.062 0 -3.0 1e-06 
3.0 0.062 0 -3.0 1e-06 
0.05 0.063 0 -3.0 1e-06 
3.0 0.063 0 -3.0 1e-06 
0.05 0.064 0 -3.0 1e-06 
3.0 0.064 0 -3.0 1e-06 
0.05 0.065 0 -3.0 1e-06 
3.0 0.065 0 -3.0 1e-06 
0.05 0.066 0 -3.0 1e-06 
3.0 0.066 0 -3.0 1e-06 
0.05 0.067 0 -3.0 1e-06 
3.0 0.067 0 -3.0 1e-06 
0.05 0.068 0 -3.0 1e-06 
3.0 0.068 0 -3.0 1e-06 
0.05 0.069 0 -3.0 1e-06 
3.0 0.069 0 -3.0 1e-06 
0.05 0.07 0 -3.0 1e-06 
3.0 0.07 0 -3.0 1e-06 
0.05 0.071 0 -3.0 1e-06 
3.0 0.071 0 -3.0 1e-06 
0.05 0.072 0 -3.0 1e-06 
3.0 0.072 0 -3.0 1e-06 
0.05 0.073 0 -3.0 1e-06 
3.0 0.073 0 -3.0 1e-06 
0.05 0.074 0 -3.0 1e-06 
3.0 0.074 0 -3.0 1e-06 
0.05 0.075 0 -3.0 1e-06 
3.0 0.075 0 -3.0 1e-06 
0.05 0.076 0 -3.0 1e-06 
3.0 0.076 0 -3.0 1e-06 
0.05 0.077 0 -3.0 1e-06 
3.0 0.077 0 -3.0 1e-06 
0.05 0.078 0 -3.0 1e-06 
3.0 0.078 0 -3.0 1e-06 
0.05 0.079 0 -3.0 1e-06 
3.0 0.079 0 -3.0 1e-06 
0.05 0.08 0 -3.0 1e-06 
3.0 0.08 0 -3.0 1e-06 
0.05 0.081 0 -3.0 1e-06 
3.0 0.081 0 -3.0 1e-06 
0.05 0.082 0 -3.0 1e-06 
3.0 0.082 0 -3.0 1e-06 
0.05 0.083 0 -3.0 1e-06 
3.0 0.083 0 -3.0 1e-06 
0.05 0.084 0 -3.0 1e-06 
3.0 0.084 0 -3.0 1e-06 
0.05 0.085 0 -3.0 1e-06 
3.0 0.085 0 -3.0 1e-06 
0.05 0.086 0 -3.0 1e-06 
3.0 0.086 0 -3.0 1e-06 
0.05 0.087 0 -3.0 1e-06 
3.0 0.087 0 -3.0 1e-06 
0.05 0.088 0 -3.0 1e-06 
3.0 0.088 0 -3.0 1e-06 
0.05 0.089 0 -3.0 1e-06 
3.0 0.089 0 -3.0 1e-06 
0.05 0.09 0 -3.0 1e-06 
3.0 0.09 0 -3.0 1e-06 
0.05 0.091 0 -3.0 1e-06 
3.0 0.091 0 -3.0 1e-06 
0.05 0.092 0 -3.0 1e-06 
3.0 0.092 0 -3.0 1e-06 
0.05 0.093 0 -3.0 1e-06 
3.0 0.093 0 -3.0 1e-06 
0.05 0.094 0 -3.0 1e-06 
3.0 0.094 0 -3.0 1e-06 
0.05 0.095 0 -3.0 1e-06 
3.0 0.095 0 -3.0 1e-06 
0.05 0.096 0 -3.0 1e-06 
3.0 0.096 0 -3.0 1e-06 
0.05 0.097 0 -3.0 1e-06 
3.0 0.097 0 -3.0 1e-06 
0.05 0.098 0 -3.0 1e-06 
3.0 0.098 0 -3.0 1e-06 
0.05 0.099 0 -3.0 1e-06 
3.0 0.099 0 -3.0 1e-06 
0.05 0.1 0 -3.0 1e-06 
3.0 0.1 0 -3.0 1e-06 
0.05 0.101 0 -3.0 1e-06 
3.0 0.101 0 -3.0 1e-06 
0.05 0.102 0 -3.0 1e-06 
3.0 0.102 0 -3.0 1e-06 
0.05 0.103 0 -3.0 1e-06 
3.0 0.103 0 -3.0 1e-06 
0.05 0.104 0 -3.0 1e-06 
3.0 0.104 0 -3.0 1e-06 
0.05 0.105 0 -3.0 1e-06 
3.0 0.105 0 -3.0 1e-06 
0.05 0.106 0 -3.0 1e-06 
3.0 0.106 0 -3.0 1e-06 
0.05 0.107 0 -3.0 1e-06 
3.0 0.107 0 -3.0 1e-06 
0.05 0.108 0 -3.0 1e-06 
3.0 0.108 0 -3.0 1e-06 
0.05 0.109 0 -3.0 1e-06 
3.0 0.109 0 -3.0 1e-06 
0.05 0.11 0 -3.0 1e-06 
3.0 0.11 0 -3.0 1e-06 
0.05 0.111 0 -3.0 1e-06 
3.0 0.111 0 -3.0 1e-06 
0.05 0.112 0 -3.0 1e-06 
3.0 0.112 0 -3.0 1e-06 
0.05 0.113 0 -3.0 1e-06 
3.0 0.113 0 -3.0 1e-06 
0.05 0.114 0 -3.0 1e-06 
3.0 0.114 0 -3.0 1e-06 
0.05 0.115 0 -3.0 1e-06 
3.0 0.115 0 -3.0 1e-06 
0.05 0.116 0 -3.0 1e-06 
3.0 0.116 0 -3.0 1e-06 
0.05 0.117 0 -3.0 1e-06 
3.0 0.117 0 -3.0 1e-06 
0.05 0.118 0 -3.0 1e-06 
3.0 0.118 0 -3.0 1e-06 
0.05 0.119 0 -3.0 1e-06 
3.0 0.119 0 -3.0 1e-06 
0.05 0.12 0 -3.0 1e-06 
3.0 0.12 0 -3.0 1e-06 
0.05 0.121 0 -3.0 1e-06 
3.0 0.121 0 -3.0 1e-06 
0.05 0.122 0 -3.0 1e-06 
3.0 0.122 0 -3.0 1e-06 
0.05 0.123 0 -3.0 1e-06 
3.0 0.123 0 -3.0 1e-06 
0.05 0.124 0 -3.0 1e-06 
3.0 0.124 0 -3.0 1e-06 
0.05 0.125 0 -3.0 1e-06 
3.0 0.125 0 -3.0 1e-06 
0.05 0.126 0 -3.0 1e-06 
3.0 0.126 0 -3.0 1e-06 
0.05 0.127 0 -3.0 1e-06 
3.0 0.127 0 -3.0 1e-06 
0.05 0.128 0 -3.0 1e-06 
3.0 0.128 0 -3.0 1e-06 
0.05 0.129 0 -3.0 1e-06 
3.0 0.129 0 -3.0 1e-06 
0.05 0.13 0 -3.0 1e-06 
3.0 0.13 0 -3.0 1e-06 
0.05 0.131 0 -3.0 1e-06 
3.0 0.131 0 -3.0 1e-06 
0.05 0.132 0 -3.0 1e-06 
3.0 0.132 0 -3.0 1e-06 
0.05 0.133 0 -3.0 1e-06 
3.0 0.133 0 -3.0 1e-06 
0.05 0.134 0 -3.0 1e-06 
3.0 0.134 0 -3.0 1e-06 
0.05 0.135 0 -3.0 1e-06 
3.0 0.135 0 -3.0 1e-06 
0.05 0.136 0 -3.0 1e-06 
3.0 0.136 0 -3.0 1e-06 
0.05 0.137 0 -3.0 1e-06 
3.0 0.137 0 -3.0 1e-06 
0.05 0.138 0 -3.0 1e-06 
3.0 0.138 0 -3.0 1e-06 
0.05 0.139 0 -3.0 1e-06 
3.0 0.139 0 -3.0 1e-06 
0.05 0.14 0 -3.0 1e-06 
3.0 0.14 0 -3.0 1e-06 
0.05 0.141 0 -3.0 1e-06 
3.0 0.141 0 -3.0 1e-06 
0.05 0.142 0 -3.0 1e-06 
3.0 0.142 0 -3.0 1e-06 
0.05 0.143 0 -3.0 1e-06 
3.0 0.143 0 -3.0 1e-06 
0.05 0.144 0 -3.0 1e-06 
3.0 0.144 0 -3.0 1e-06 
0.05 0.145 0 -3.0 1e-06 
3.0 0.145 0 -3.0 1e-06 
0.05 0.146 0 -3.0 1e-06 
3.0 0.146 0 -3.0 1e-06 
0.05 0.147 0 -3.0 1e-06 
3.0 0.147 0 -3.0 1e-06 
0.05 0.148 0 -3.0 1e-06 
3.0 0.148 0 -3.0 1e-06 
0.05 0.149 0 -3.0 1e-06 
3.0 0.149 0 -3.0 1e-06 
0.05 0.15 0 -3.0 1e-06 
3.0 0.15 0 -3.0 1e-06 
0.05 0.151 0 -3.0 1e-06 
3.0 0.151 0 -3.0 1e-06 
0.05 0.152 0 -3.0 1e-06 
3.0 0.152 0 -3.0 1e-06 
0.05 0.153 0 -3.0 1e-06 
3.0 0.153 0 -3.0 1e-06 
0.05 0.154 0 -3.0 1e-06 
3.0 0.154 0 -3.0 1e-06 
0.05 0.155 0 -3.0 1e-06 
3.0 0.155 0 -3.0 1e-06 
0.05 0.156 0 -3.0 1e-06 
3.0 0.156 0 -3.0 1e-06 
0.05 0.157 0 -3.0 1e-06 
3.0 0.157 0 -3.0 1e-06 
0.05 0.158 0 -3.0 1e-06 
3.0 0.158 0 -3.0 1e-06 
0.05 0.159 0 -3.0 1e-06 
3.0 0.159 0 -3.0 1e-06 
0.05 0.16 0 -3.0 1e-06 
3.0 0.16 0 -3.0 1e-06 
0.05 0.161 0 -3.0 1e-06 
3.0 0.161 0 -3.0 1e-06 
0.05 0.162 0 -3.0 1e-06 
3.0 0.162 0 -3.0 1e-06 
0.05 0.163 0 -3.0 1e-06 
3.0 0.163 0 -3.0 1e-06 
0.05 0.164 0 -3.0 1e-06 
3.0 0.164 0 -3.0 1e-06 
0.05 0.165 0 -3.0 1e-06 
3.0 0.165 0 -3.0 1e-06 
0.05 0.166 0 -3.0 1e-06 
3.0 0.166 0 -3.0 1e-06 
0.05 0.167 0 -3.0 1e-06 
3.0 0.167 0 -3.0 1e-06 
0.05 0.168 0 -3.0 1e-06 
3.0 0.168 0 -3.0 1e-06 
0.05 0.169 0 -3.0 1e-06 
3.0 0.169 0 -3.0 1e-06 
0.05 0.17 0 -3.0 1e-06 
3.0 0.17 0 -3.0 1e-06 
0.05 0.171 0 -3.0 1e-06 
3.0 0.171 0 -3.0 1e-06 
0.05 0.172 0 -3.0 1e-06 
3.0 0.172 0 -3.0 1e-06 
0.05 0.173 0 -3.0 1e-06 
3.0 0.173 0 -3.0 1e-06 
0.05 0.174 0 -3.0 1e-06 
3.0 0.174 0 -3.0 1e-06 
0.05 0.175 0 -3.0 1e-06 
3.0 0.175 0 -3.0 1e-06 
0.05 0.176 0 -3.0 1e-06 
3.0 0.176 0 -3.0 1e-06 
0.05 0.177 0 -3.0 1e-06 
3.0 0.177 0 -3.0 1e-06 
0.05 0.178 0 -3.0 1e-06 
3.0 0.178 0 -3.0 1e-06 
0.05 0.179 0 -3.0 1e-06 
3.0 0.179 0 -3.0 1e-06 
0.05 0.18 0 -3.0 1e-06 
3.0 0.18 0 -3.0 1e-06 
0.05 0.181 0 -3.0 1e-06 
3.0 0.181 0 -3.0 1e-06 
0.05 0.182 0 -3.0 1e-06 
3.0 0.182 0 -3.0 1e-06 
0.05 0.183 0 -3.0 1e-06 
3.0 0.183 0 -3.0 1e-06 
0.05 0.184 0 -3.0 1e-06 
3.0 0.184 0 -3.0 1e-06 
0.05 0.185 0 -3.0 1e-06 
3.0 0.185 0 -3.0 1e-06 
0.05 0.186 0 -3.0 1e-06 
3.0 0.186 0 -3.0 1e-06 
0.05 0.187 0 -3.0 1e-06 
3.0 0.187 0 -3.0 1e-06 
0.05 0.188 0 -3.0 1e-06 
3.0 0.188 0 -3.0 1e-06 
0.05 0.189 0 -3.0 1e-06 
3.0 0.189 0 -3.0 1e-06 
0.05 0.19 0 -3.0 1e-06 
3.0 0.19 0 -3.0 1e-06 
0.05 0.191 0 -3.0 1e-06 
3.0 0.191 0 -3.0 1e-06 
0.05 0.192 0 -3.0 1e-06 
3.0 0.192 0 -3.0 1e-06 
0.05 0.193 0 -3.0 1e-06 
3.0 0.193 0 -3.0 1e-06 
0.05 0.194 0 -3.0 1e-06 
3.0 0.194 0 -3.0 1e-06 
0.05 0.195 0 -3.0 1e-06 
3.0 0.195 0 -3.0 1e-06 
0.05 0.196 0 -3.0 1e-06 
3.0 0.196 0 -3.0 1e-06 
0.05 0.197 0 -3.0 1e-06 
3.0 0.197 0 -3.0 1e-06 
0.05 0.198 0 -3.0 1e-06 
3.0 0.198 0 -3.0 1e-06 
0.05 0.199 0 -3.0 1e-06 
3.0 0.199 0 -3.0 1e-06 
0.05 0.2 0 -3.0 1e-06 
3.0 0.2 0 -3.0 1e-06 
0.05 0.201 0 -3.0 1e-06 
3.0 0.201 0 -3.0 1e-06 
0.05 0.202 0 -3.0 1e-06 
3.0 0.202 0 -3.0 1e-06 
0.05 0.203 0 -3.0 1e-06 
3.0 0.203 0 -3.0 1e-06 
0.05 0.204 0 -3.0 1e-06 
3.0 0.204 0 -3.0 1e-06 
0.05 0.205 0 -3.0 1e-06 
3.0 0.205 0 -3.0 1e-06 
0.05 0.206 0 -3.0 1e-06 
3.0 0.206 0 -3.0 1e-06 
0.05 0.207 0 -3.0 1e-06 
3.0 0.207 0 -3.0 1e-06 
0.05 0.208 0 -3.0 1e-06 
3.0 0.208 0 -3.0 1e-06 
0.05 0.209 0 -3.0 1e-06 
3.0 0.209 0 -3.0 1e-06 
0.05 0.21 0 -3.0 1e-06 
3.0 0.21 0 -3.0 1e-06 
0.05 0.211 0 -3.0 1e-06 
3.0 0.211 0 -3.0 1e-06 
0.05 0.212 0 -3.0 1e-06 
3.0 0.212 0 -3.0 1e-06 
0.05 0.213 0 -3.0 1e-06 
3.0 0.213 0 -3.0 1e-06 
0.05 0.214 0 -3.0 1e-06 
3.0 0.214 0 -3.0 1e-06 
0.05 0.215 0 -3.0 1e-06 
3.0 0.215 0 -3.0 1e-06 
0.05 0.216 0 -3.0 1e-06 
3.0 0.216 0 -3.0 1e-06 
0.05 0.217 0 -3.0 1e-06 
3.0 0.217 0 -3.0 1e-06 
0.05 0.218 0 -3.0 1e-06 
3.0 0.218 0 -3.0 1e-06 
0.05 0.219 0 -3.0 1e-06 
3.0 0.219 0 -3.0 1e-06 
0.05 0.22 0 -3.0 1e-06 
3.0 0.22 0 -3.0 1e-06 
0.05 0.221 0 -3.0 1e-06 
3.0 0.221 0 -3.0 1e-06 
0.05 0.222 0 -3.0 1e-06 
3.0 0.222 0 -3.0 1e-06 
0.05 0.223 0 -3.0 1e-06 
3.0 0.223 0 -3.0 1e-06 
0.05 0.224 0 -3.0 1e-06 
3.0 0.224 0 -3.0 1e-06 
0.05 0.225 0 -3.0 1e-06 
3.0 0.225 0 -3.0 1e-06 
0.05 0.226 0 -3.0 1e-06 
3.0 0.226 0 -3.0 1e-06 
0.05 0.227 0 -3.0 1e-06 
3.0 0.227 0 -3.0 1e-06 
0.05 0.228 0 -3.0 1e-06 
3.0 0.228 0 -3.0 1e-06 
0.05 0.229 0 -3.0 1e-06 
3.0 0.229 0 -3.0 1e-06 
0.05 0.23 0 -3.0 1e-06 
3.0 0.23 0 -3.0 1e-06 
0.05 0.231 0 -3.0 1e-06 
3.0 0.231 0 -3.0 1e-06 
0.05 0.232 0 -3.0 1e-06 
3.0 0.232 0 -3.0 1e-06 
0.05 0.233 0 -3.0 1e-06 
3.0 0.233 0 -3.0 1e-06 
0.05 0.234 0 -3.0 1e-06 
3.0 0.234 0 -3.0 1e-06 
0.05 0.235 0 -3.0 1e-06 
3.0 0.235 0 -3.0 1e-06 
0.05 0.236 0 -3.0 1e-06 
3.0 0.236 0 -3.0 1e-06 
0.05 0.237 0 -3.0 1e-06 
3.0 0.237 0 -3.0 1e-06 
0.05 0.238 0 -3.0 1e-06 
3.0 0.238 0 -3.0 1e-06 
0.05 0.239 0 -3.0 1e-06 
3.0 0.239 0 -3.0 1e-06 
0.05 0.24 0 -3.0 1e-06 
3.0 0.24 0 -3.0 1e-06 
0.05 0.241 0 -3.0 1e-06 
3.0 0.241 0 -3.0 1e-06 
0.05 0.242 0 -3.0 1e-06 
3.0 0.242 0 -3.0 1e-06 
0.05 0.243 0 -3.0 1e-06 
3.0 0.243 0 -3.0 1e-06 
0.05 0.244 0 -3.0 1e-06 
3.0 0.244 0 -3.0 1e-06 
0.05 0.245 0 -3.0 1e-06 
3.0 0.245 0 -3.0 1e-06 
0.05 0.246 0 -3.0 1e-06 
3.0 0.246 0 -3.0 1e-06 
0.05 0.247 0 -3.0 1e-06 
3.0 0.247 0 -3.0 1e-06 
0.05 0.248 0 -3.0 1e-06 
3.0 0.248 0 -3.0 1e-06 
0.05 0.249 0 -3.0 1e-06 
3.0 0.249 0 -3.0 1e-06 
0.05 0.25 0 -3.0 1e-06 
3.0 0.25 0 -3.0 1e-06 
0.05 0.251 0 -3.0 1e-06 
3.0 0.251 0 -3.0 1e-06 
0.05 0.252 0 -3.0 1e-06 
3.0 0.252 0 -3.0 1e-06 
0.05 0.253 0 -3.0 1e-06 
3.0 0.253 0 -3.0 1e-06 
0.05 0.254 0 -3.0 1e-06 
3.0 0.254 0 -3.0 1e-06 
0.05 0.255 0 -3.0 1e-06 
3.0 0.255 0 -3.0 1e-06 
0.05 0.256 0 -3.0 1e-06 
3.0 0.256 0 -3.0 1e-06 
0.05 0.257 0 -3.0 1e-06 
3.0 0.257 0 -3.0 1e-06 
0.05 0.258 0 -3.0 1e-06 
3.0 0.258 0 -3.0 1e-06 
0.05 0.259 0 -3.0 1e-06 
3.0 0.259 0 -3.0 1e-06 
0.05 0.26 0 -3.0 1e-06 
3.0 0.26 0 -3.0 1e-06 
0.05 0.261 0 -3.0 1e-06 
3.0 0.261 0 -3.0 1e-06 
0.05 0.262 0 -3.0 1e-06 
3.0 0.262 0 -3.0 1e-06 
0.05 0.263 0 -3.0 1e-06 
3.0 0.263 0 -3.0 1e-06 
0.05 0.264 0 -3.0 1e-06 
3.0 0.264 0 -3.0 1e-06 
0.05 0.265 0 -3.0 1e-06 
3.0 0.265 0 -3.0 1e-06 
0.05 0.266 0 -3.0 1e-06 
3.0 0.266 0 -3.0 1e-06 
0.05 0.267 0 -3.0 1e-06 
3.0 0.267 0 -3.0 1e-06 
0.05 0.268 0 -3.0 1e-06 
3.0 0.268 0 -3.0 1e-06 
0.05 0.269 0 -3.0 1e-06 
3.0 0.269 0 -3.0 1e-06 
0.05 0.27 0 -3.0 1e-06 
3.0 0.27 0 -3.0 1e-06 
0.05 0.271 0 -3.0 1e-06 
3.0 0.271 0 -3.0 1e-06 
0.05 0.272 0 -3.0 1e-06 
3.0 0.272 0 -3.0 1e-06 
0.05 0.273 0 -3.0 1e-06 
3.0 0.273 0 -3.0 1e-06 
0.05 0.274 0 -3.0 1e-06 
3.0 0.274 0 -3.0 1e-06 
0.05 0.275 0 -3.0 1e-06 
3.0 0.275 0 -3.0 1e-06 
0.05 0.276 0 -3.0 1e-06 
3.0 0.276 0 -3.0 1e-06 
0.05 0.277 0 -3.0 1e-06 
3.0 0.277 0 -3.0 1e-06 
0.05 0.278 0 -3.0 1e-06 
3.0 0.278 0 -3.0 1e-06 
0.05 0.279 0 -3.0 1e-06 
3.0 0.279 0 -3.0 1e-06 
0.05 0.28 0 -3.0 1e-06 
3.0 0.28 0 -3.0 1e-06 
0.05 0.281 0 -3.0 1e-06 
3.0 0.281 0 -3.0 1e-06 
0.05 0.282 0 -3.0 1e-06 
3.0 0.282 0 -3.0 1e-06 
0.05 0.283 0 -3.0 1e-06 
3.0 0.283 0 -3.0 1e-06 
0.05 0.284 0 -3.0 1e-06 
3.0 0.284 0 -3.0 1e-06 
0.05 0.285 0 -3.0 1e-06 
3.0 0.285 0 -3.0 1e-06 
0.05 0.286 0 -3.0 1e-06 
3.0 0.286 0 -3.0 1e-06 
0.05 0.287 0 -3.0 1e-06 
3.0 0.287 0 -3.0 1e-06 
0.05 0.288 0 -3.0 1e-06 
3.0 0.288 0 -3.0 1e-06 
0.05 0.289 0 -3.0 1e-06 
3.0 0.289 0 -3.0 1e-06 
0.05 0.29 0 -3.0 1e-06 
3.0 0.29 0 -3.0 1e-06 
0.05 0.291 0 -3.0 1e-06 
3.0 0.291 0 -3.0 1e-06 
0.05 0.292 0 -3.0 1e-06 
3.0 0.292 0 -3.0 1e-06 
0.05 0.293 0 -3.0 1e-06 
3.0 0.293 0 -3.0 1e-06 
0.05 0.294 0 -3.0 1e-06 
3.0 0.294 0 -3.0 1e-06 
0.05 0.295 0 -3.0 1e-06 
3.0 0.295 0 -3.0 1e-06 
0.05 0.296 0 -3.0 1e-06 
3.0 0.296 0 -3.0 1e-06 
0.05 0.297 0 -3.0 1e-06 
3.0 0.297 0 -3.0 1e-06 
0.05 0.298 0 -3.0 1e-06 
3.0 0.298 0 -3.0 1e-06 
0.05 0.299 0 -3.0 1e-06 
3.0 0.299 0 -3.0 1e-06 
0.05 0.3 0 -3.0 1e-06 
3.0 0.3 0 -3.0 1e-06 
0.05 0.301 0 -3.0 1e-06 
3.0 0.301 0 -3.0 1e-06 
0.05 0.302 0 -3.0 1e-06 
3.0 0.302 0 -3.0 1e-06 
0.05 0.303 0 -3.0 1e-06 
3.0 0.303 0 -3.0 1e-06 
0.05 0.304 0 -3.0 1e-06 
3.0 0.304 0 -3.0 1e-06 
0.05 0.305 0 -3.0 1e-06 
3.0 0.305 0 -3.0 1e-06 
0.05 0.306 0 -3.0 1e-06 
3.0 0.306 0 -3.0 1e-06 
0.05 0.307 0 -3.0 1e-06 
3.0 0.307 0 -3.0 1e-06 
0.05 0.308 0 -3.0 1e-06 
3.0 0.308 0 -3.0 1e-06 
0.05 0.309 0 -3.0 1e-06 
3.0 0.309 0 -3.0 1e-06 
0.05 0.31 0 -3.0 1e-06 
3.0 0.31 0 -3.0 1e-06 
0.05 0.311 0 -3.0 1e-06 
3.0 0.311 0 -3.0 1e-06 
0.05 0.312 0 -3.0 1e-06 
3.0 0.312 0 -3.0 1e-06 
0.05 0.313 0 -3.0 1e-06 
3.0 0.313 0 -3.0 1e-06 
0.05 0.314 0 -3.0 1e-06 
3.0 0.314 0 -3.0 1e-06 
0.05 0.315 0 -3.0 1e-06 
3.0 0.315 0 -3.0 1e-06 
0.05 0.316 0 -3.0 1e-06 
3.0 0.316 0 -3.0 1e-06 
0.05 0.317 0 -3.0 1e-06 
3.0 0.317 0 -3.0 1e-06 
0.05 0.318 0 -3.0 1e-06 
3.0 0.318 0 -3.0 1e-06 
0.05 0.319 0 -3.0 1e-06 
3.0 0.319 0 -3.0 1e-06 
0.05 0.32 0 -3.0 1e-06 
3.0 0.32 0 -3.0 1e-06 
0.05 0.321 0 -3.0 1e-06 
3.0 0.321 0 -3.0 1e-06 
0.05 0.322 0 -3.0 1e-06 
3.0 0.322 0 -3.0 1e-06 
0.05 0.323 0 -3.0 1e-06 
3.0 0.323 0 -3.0 1e-06 
0.05 0.324 0 -3.0 1e-06 
3.0 0.324 0 -3.0 1e-06 
0.05 0.325 0 -3.0 1e-06 
3.0 0.325 0 -3.0 1e-06 
0.05 0.326 0 -3.0 1e-06 
3.0 0.326 0 -3.0 1e-06 
0.05 0.327 0 -3.0 1e-06 
3.0 0.327 0 -3.0 1e-06 
0.05 0.328 0 -3.0 1e-06 
3.0 0.328 0 -3.0 1e-06 
0.05 0.329 0 -3.0 1e-06 
3.0 0.329 0 -3.0 1e-06 
0.05 0.33 0 -3.0 1e-06 
3.0 0.33 0 -3.0 1e-06 
0.05 0.331 0 -3.0 1e-06 
3.0 0.331 0 -3.0 1e-06 
0.05 0.332 0 -3.0 1e-06 
3.0 0.332 0 -3.0 1e-06 
0.05 0.333 0 -3.0 1e-06 
3.0 0.333 0 -3.0 1e-06 
0.05 0.334 0 -3.0 1e-06 
3.0 0.334 0 -3.0 1e-06 
0.05 0.335 0 -3.0 1e-06 
3.0 0.335 0 -3.0 1e-06 
0.05 0.336 0 -3.0 1e-06 
3.0 0.336 0 -3.0 1e-06 
0.05 0.337 0 -3.0 1e-06 
3.0 0.337 0 -3.0 1e-06 
0.05 0.338 0 -3.0 1e-06 
3.0 0.338 0 -3.0 1e-06 
0.05 0.339 0 -3.0 1e-06 
3.0 0.339 0 -3.0 1e-06 
0.05 0.34 0 -3.0 1e-06 
3.0 0.34 0 -3.0 1e-06 
0.05 0.341 0 -3.0 1e-06 
3.0 0.341 0 -3.0 1e-06 
0.05 0.342 0 -3.0 1e-06 
3.0 0.342 0 -3.0 1e-06 
0.05 0.343 0 -3.0 1e-06 
3.0 0.343 0 -3.0 1e-06 
0.05 0.344 0 -3.0 1e-06 
3.0 0.344 0 -3.0 1e-06 
0.05 0.345 0 -3.0 1e-06 
3.0 0.345 0 -3.0 1e-06 
0.05 0.346 0 -3.0 1e-06 
3.0 0.346 0 -3.0 1e-06 
0.05 0.347 0 -3.0 1e-06 
3.0 0.347 0 -3.0 1e-06 
0.05 0.348 0 -3.0 1e-06 
3.0 0.348 0 -3.0 1e-06 
0.05 0.349 0 -3.0 1e-06 
3.0 0.349 0 -3.0 1e-06 
0.05 0.35 0 -3.0 1e-06 
3.0 0.35 0 -3.0 1e-06 
0.05 0.351 0 -3.0 1e-06 
3.0 0.351 0 -3.0 1e-06 
0.05 0.352 0 -3.0 1e-06 
3.0 0.352 0 -3.0 1e-06 
0.05 0.353 0 -3.0 1e-06 
3.0 0.353 0 -3.0 1e-06 
0.05 0.354 0 -3.0 1e-06 
3.0 0.354 0 -3.0 1e-06 
0.05 0.355 0 -3.0 1e-06 
3.0 0.355 0 -3.0 1e-06 
0.05 0.356 0 -3.0 1e-06 
3.0 0.356 0 -3.0 1e-06 
0.05 0.357 0 -3.0 1e-06 
3.0 0.357 0 -3.0 1e-06 
0.05 0.358 0 -3.0 1e-06 
3.0 0.358 0 -3.0 1e-06 
0.05 0.359 0 -3.0 1e-06 
3.0 0.359 0 -3.0 1e-06 
0.05 0.36 0 -3.0 1e-06 
3.0 0.36 0 -3.0 1e-06 
0.05 0.361 0 -3.0 1e-06 
3.0 0.361 0 -3.0 1e-06 
0.05 0.362 0 -3.0 1e-06 
3.0 0.362 0 -3.0 1e-06 
0.05 0.363 0 -3.0 1e-06 
3.0 0.363 0 -3.0 1e-06 
0.05 0.364 0 -3.0 1e-06 
3.0 0.364 0 -3.0 1e-06 
0.05 0.365 0 -3.0 1e-06 
3.0 0.365 0 -3.0 1e-06 
0.05 0.366 0 -3.0 1e-06 
3.0 0.366 0 -3.0 1e-06 
0.05 0.367 0 -3.0 1e-06 
3.0 0.367 0 -3.0 1e-06 
0.05 0.368 0 -3.0 1e-06 
3.0 0.368 0 -3.0 1e-06 
0.05 0.369 0 -3.0 1e-06 
3.0 0.369 0 -3.0 1e-06 
0.05 0.37 0 -3.0 1e-06 
3.0 0.37 0 -3.0 1e-06 
0.05 0.371 0 -3.0 1e-06 
3.0 0.371 0 -3.0 1e-06 
0.05 0.372 0 -3.0 1e-06 
3.0 0.372 0 -3.0 1e-06 
0.05 0.373 0 -3.0 1e-06 
3.0 0.373 0 -3.0 1e-06 
0.05 0.374 0 -3.0 1e-06 
3.0 0.374 0 -3.0 1e-06 
0.05 0.375 0 -3.0 1e-06 
3.0 0.375 0 -3.0 1e-06 
0.05 0.376 0 -3.0 1e-06 
3.0 0.376 0 -3.0 1e-06 
0.05 0.377 0 -3.0 1e-06 
3.0 0.377 0 -3.0 1e-06 
0.05 0.378 0 -3.0 1e-06 
3.0 0.378 0 -3.0 1e-06 
0.05 0.379 0 -3.0 1e-06 
3.0 0.379 0 -3.0 1e-06 
0.05 0.38 0 -3.0 1e-06 
3.0 0.38 0 -3.0 1e-06 
0.05 0.381 0 -3.0 1e-06 
3.0 0.381 0 -3.0 1e-06 
0.05 0.382 0 -3.0 1e-06 
3.0 0.382 0 -3.0 1e-06 
0.05 0.383 0 -3.0 1e-06 
3.0 0.383 0 -3.0 1e-06 
0.05 0.384 0 -3.0 1e-06 
3.0 0.384 0 -3.0 1e-06 
0.05 0.385 0 -3.0 1e-06 
3.0 0.385 0 -3.0 1e-06 
0.05 0.386 0 -3.0 1e-06 
3.0 0.386 0 -3.0 1e-06 
0.05 0.387 0 -3.0 1e-06 
3.0 0.387 0 -3.0 1e-06 
0.05 0.388 0 -3.0 1e-06 
3.0 0.388 0 -3.0 1e-06 
0.05 0.389 0 -3.0 1e-06 
3.0 0.389 0 -3.0 1e-06 
0.05 0.39 0 -3.0 1e-06 
3.0 0.39 0 -3.0 1e-06 
0.05 0.391 0 -3.0 1e-06 
3.0 0.391 0 -3.0 1e-06 
0.05 0.392 0 -3.0 1e-06 
3.0 0.392 0 -3.0 1e-06 
0.05 0.393 0 -3.0 1e-06 
3.0 0.393 0 -3.0 1e-06 
0.05 0.394 0 -3.0 1e-06 
3.0 0.394 0 -3.0 1e-06 
0.05 0.395 0 -3.0 1e-06 
3.0 0.395 0 -3.0 1e-06 
0.05 0.396 0 -3.0 1e-06 
3.0 0.396 0 -3.0 1e-06 
0.05 0.397 0 -3.0 1e-06 
3.0 0.397 0 -3.0 1e-06 
0.05 0.398 0 -3.0 1e-06 
3.0 0.398 0 -3.0 1e-06 
0.05 0.399 0 -3.0 1e-06 
3.0 0.399 0 -3.0 1e-06 
0.05 0.4 0 -3.0 1e-06 
3.0 0.4 0 -3.0 1e-06 
0.05 0.401 0 -3.0 1e-06 
3.0 0.401 0 -3.0 1e-06 
0.05 0.402 0 -3.0 1e-06 
3.0 0.402 0 -3.0 1e-06 
0.05 0.403 0 -3.0 1e-06 
3.0 0.403 0 -3.0 1e-06 
0.05 0.404 0 -3.0 1e-06 
3.0 0.404 0 -3.0 1e-06 
0.05 0.405 0 -3.0 1e-06 
3.0 0.405 0 -3.0 1e-06 
0.05 0.406 0 -3.0 1e-06 
3.0 0.406 0 -3.0 1e-06 
0.05 0.407 0 -3.0 1e-06 
3.0 0.407 0 -3.0 1e-06 
0.05 0.408 0 -3.0 1e-06 
3.0 0.408 0 -3.0 1e-06 
0.05 0.409 0 -3.0 1e-06 
3.0 0.409 0 -3.0 1e-06 
0.05 0.41 0 -3.0 1e-06 
3.0 0.41 0 -3.0 1e-06 
0.05 0.411 0 -3.0 1e-06 
3.0 0.411 0 -3.0 1e-06 
0.05 0.412 0 -3.0 1e-06 
3.0 0.412 0 -3.0 1e-06 
0.05 0.413 0 -3.0 1e-06 
3.0 0.413 0 -3.0 1e-06 
0.05 0.414 0 -3.0 1e-06 
3.0 0.414 0 -3.0 1e-06 
0.05 0.415 0 -3.0 1e-06 
3.0 0.415 0 -3.0 1e-06 
0.05 0.416 0 -3.0 1e-06 
3.0 0.416 0 -3.0 1e-06 
0.05 0.417 0 -3.0 1e-06 
3.0 0.417 0 -3.0 1e-06 
0.05 0.418 0 -3.0 1e-06 
3.0 0.418 0 -3.0 1e-06 
0.05 0.419 0 -3.0 1e-06 
3.0 0.419 0 -3.0 1e-06 
0.05 0.42 0 -3.0 1e-06 
3.0 0.42 0 -3.0 1e-06 
0.05 0.421 0 -3.0 1e-06 
3.0 0.421 0 -3.0 1e-06 
0.05 0.422 0 -3.0 1e-06 
3.0 0.422 0 -3.0 1e-06 
0.05 0.423 0 -3.0 1e-06 
3.0 0.423 0 -3.0 1e-06 
0.05 0.424 0 -3.0 1e-06 
3.0 0.424 0 -3.0 1e-06 
0.05 0.425 0 -3.0 1e-06 
3.0 0.425 0 -3.0 1e-06 
0.05 0.426 0 -3.0 1e-06 
3.0 0.426 0 -3.0 1e-06 
0.05 0.427 0 -3.0 1e-06 
3.0 0.427 0 -3.0 1e-06 
0.05 0.428 0 -3.0 1e-06 
3.0 0.428 0 -3.0 1e-06 
0.05 0.429 0 -3.0 1e-06 
3.0 0.429 0 -3.0 1e-06 
0.05 0.43 0 -3.0 1e-06 
3.0 0.43 0 -3.0 1e-06 
0.05 0.431 0 -3.0 1e-06 
3.0 0.431 0 -3.0 1e-06 
0.05 0.432 0 -3.0 1e-06 
3.0 0.432 0 -3.0 1e-06 
0.05 0.433 0 -3.0 1e-06 
3.0 0.433 0 -3.0 1e-06 
0.05 0.434 0 -3.0 1e-06 
3.0 0.434 0 -3.0 1e-06 
0.05 0.435 0 -3.0 1e-06 
3.0 0.435 0 -3.0 1e-06 
0.05 0.436 0 -3.0 1e-06 
3.0 0.436 0 -3.0 1e-06 
0.05 0.437 0 -3.0 1e-06 
3.0 0.437 0 -3.0 1e-06 
0.05 0.438 0 -3.0 1e-06 
3.0 0.438 0 -3.0 1e-06 
0.05 0.439 0 -3.0 1e-06 
3.0 0.439 0 -3.0 1e-06 
0.05 0.44 0 -3.0 1e-06 
3.0 0.44 0 -3.0 1e-06 
0.05 0.441 0 -3.0 1e-06 
3.0 0.441 0 -3.0 1e-06 
0.05 0.442 0 -3.0 1e-06 
3.0 0.442 0 -3.0 1e-06 
0.05 0.443 0 -3.0 1e-06 
3.0 0.443 0 -3.0 1e-06 
0.05 0.444 0 -3.0 1e-06 
3.0 0.444 0 -3.0 1e-06 
0.05 0.445 0 -3.0 1e-06 
3.0 0.445 0 -3.0 1e-06 
0.05 0.446 0 -3.0 1e-06 
3.0 0.446 0 -3.0 1e-06 
0.05 0.447 0 -3.0 1e-06 
3.0 0.447 0 -3.0 1e-06 
0.05 0.448 0 -3.0 1e-06 
3.0 0.448 0 -3.0 1e-06 
0.05 0.449 0 -3.0 1e-06 
3.0 0.449 0 -3.0 1e-06 
0.05 0.45 0 -3.0 1e-06 
3.0 0.45 0 -3.0 1e-06 
0.05 0.451 0 -3.0 1e-06 
3.0 0.451 0 -3.0 1e-06 
0.05 0.452 0 -3.0 1e-06 
3.0 0.452 0 -3.0 1e-06 
0.05 0.453 0 -3.0 1e-06 
3.0 0.453 0 -3.0 1e-06 
0.05 0.454 0 -3.0 1e-06 
3.0 0.454 0 -3.0 1e-06 
0.05 0.455 0 -3.0 1e-06 
3.0 0.455 0 -3.0 1e-06 
0.05 0.456 0 -3.0 1e-06 
3.0 0.456 0 -3.0 1e-06 
0.05 0.457 0 -3.0 1e-06 
3.0 0.457 0 -3.0 1e-06 
0.05 0.458 0 -3.0 1e-06 
3.0 0.458 0 -3.0 1e-06 
0.05 0.459 0 -3.0 1e-06 
3.0 0.459 0 -3.0 1e-06 
0.05 0.46 0 -3.0 1e-06 
3.0 0.46 0 -3.0 1e-06 
0.05 0.461 0 -3.0 1e-06 
3.0 0.461 0 -3.0 1e-06 
0.05 0.462 0 -3.0 1e-06 
3.0 0.462 0 -3.0 1e-06 
0.05 0.463 0 -3.0 1e-06 
3.0 0.463 0 -3.0 1e-06 
0.05 0.464 0 -3.0 1e-06 
3.0 0.464 0 -3.0 1e-06 
0.05 0.465 0 -3.0 1e-06 
3.0 0.465 0 -3.0 1e-06 
0.05 0.466 0 -3.0 1e-06 
3.0 0.466 0 -3.0 1e-06 
0.05 0.467 0 -3.0 1e-06 
3.0 0.467 0 -3.0 1e-06 
0.05 0.468 0 -3.0 1e-06 
3.0 0.468 0 -3.0 1e-06 
0.05 0.469 0 -3.0 1e-06 
3.0 0.469 0 -3.0 1e-06 
0.05 0.47 0 -3.0 1e-06 
3.0 0.47 0 -3.0 1e-06 
0.05 0.471 0 -3.0 1e-06 
3.0 0.471 0 -3.0 1e-06 
0.05 0.472 0 -3.0 1e-06 
3.0 0.472 0 -3.0 1e-06 
0.05 0.473 0 -3.0 1e-06 
3.0 0.473 0 -3.0 1e-06 
0.05 0.474 0 -3.0 1e-06 
3.0 0.474 0 -3.0 1e-06 
0.05 0.475 0 -3.0 1e-06 
3.0 0.475 0 -3.0 1e-06 
0.05 0.476 0 -3.0 1e-06 
3.0 0.476 0 -3.0 1e-06 
0.05 0.477 0 -3.0 1e-06 
3.0 0.477 0 -3.0 1e-06 
0.05 0.478 0 -3.0 1e-06 
3.0 0.478 0 -3.0 1e-06 
0.05 0.479 0 -3.0 1e-06 
3.0 0.479 0 -3.0 1e-06 
0.05 0.48 0 -3.0 1e-06 
3.0 0.48 0 -3.0 1e-06 
0.05 0.481 0 -3.0 1e-06 
3.0 0.481 0 -3.0 1e-06 
0.05 0.482 0 -3.0 1e-06 
3.0 0.482 0 -3.0 1e-06 
0.05 0.483 0 -3.0 1e-06 
3.0 0.483 0 -3.0 1e-06 
0.05 0.484 0 -3.0 1e-06 
3.0 0.484 0 -3.0 1e-06 
0.05 0.485 0 -3.0 1e-06 
3.0 0.485 0 -3.0 1e-06 
0.05 0.486 0 -3.0 1e-06 
3.0 0.486 0 -3.0 1e-06 
0.05 0.487 0 -3.0 1e-06 
3.0 0.487 0 -3.0 1e-06 
0.05 0.488 0 -3.0 1e-06 
3.0 0.488 0 -3.0 1e-06 
0.05 0.489 0 -3.0 1e-06 
3.0 0.489 0 -3.0 1e-06 
0.05 0.49 0 -3.0 1e-06 
3.0 0.49 0 -3.0 1e-06 
0.05 0.491 0 -3.0 1e-06 
3.0 0.491 0 -3.0 1e-06 
0.05 0.492 0 -3.0 1e-06 
3.0 0.492 0 -3.0 1e-06 
0.05 0.493 0 -3.0 1e-06 
3.0 0.493 0 -3.0 1e-06 
0.05 0.494 0 -3.0 1e-06 
3.0 0.494 0 -3.0 1e-06 
0.05 0.495 0 -3.0 1e-06 
3.0 0.495 0 -3.0 1e-06 
0.05 0.496 0 -3.0 1e-06 
3.0 0.496 0 -3.0 1e-06 
0.05 0.497 0 -3.0 1e-06 
3.0 0.497 0 -3.0 1e-06 
0.05 0.498 0 -3.0 1e-06 
3.0 0.498 0 -3.0 1e-06 
0.05 0.499 0 -3.0 1e-06 
3.0 0.499 0 -3.0 1e-06 
0.05 0.5 0 -3.0 1e-06 
3.0 0.5 0 -3.0 1e-06 
0.05 0.501 0 -3.0 1e-06 
3.0 0.501 0 -3.0 1e-06 
0.05 0.502 0 -3.0 1e-06 
3.0 0.502 0 -3.0 1e-06 
0.05 0.503 0 -3.0 1e-06 
3.0 0.503 0 -3.0 1e-06 
0.05 0.504 0 -3.0 1e-06 
3.0 0.504 0 -3.0 1e-06 
0.05 0.505 0 -3.0 1e-06 
3.0 0.505 0 -3.0 1e-06 
0.05 0.506 0 -3.0 1e-06 
3.0 0.506 0 -3.0 1e-06 
0.05 0.507 0 -3.0 1e-06 
3.0 0.507 0 -3.0 1e-06 
0.05 0.508 0 -3.0 1e-06 
3.0 0.508 0 -3.0 1e-06 
0.05 0.509 0 -3.0 1e-06 
3.0 0.509 0 -3.0 1e-06 
0.05 0.51 0 -3.0 1e-06 
3.0 0.51 0 -3.0 1e-06 
0.05 0.511 0 -3.0 1e-06 
3.0 0.511 0 -3.0 1e-06 
0.05 0.512 0 -3.0 1e-06 
3.0 0.512 0 -3.0 1e-06 
0.05 0.513 0 -3.0 1e-06 
3.0 0.513 0 -3.0 1e-06 
0.05 0.514 0 -3.0 1e-06 
3.0 0.514 0 -3.0 1e-06 
0.05 0.515 0 -3.0 1e-06 
3.0 0.515 0 -3.0 1e-06 
0.05 0.516 0 -3.0 1e-06 
3.0 0.516 0 -3.0 1e-06 
0.05 0.517 0 -3.0 1e-06 
3.0 0.517 0 -3.0 1e-06 
0.05 0.518 0 -3.0 1e-06 
3.0 0.518 0 -3.0 1e-06 
0.05 0.519 0 -3.0 1e-06 
3.0 0.519 0 -3.0 1e-06 
0.05 0.52 0 -3.0 1e-06 
3.0 0.52 0 -3.0 1e-06 
0.05 0.521 0 -3.0 1e-06 
3.0 0.521 0 -3.0 1e-06 
0.05 0.522 0 -3.0 1e-06 
3.0 0.522 0 -3.0 1e-06 
0.05 0.523 0 -3.0 1e-06 
3.0 0.523 0 -3.0 1e-06 
0.05 0.524 0 -3.0 1e-06 
3.0 0.524 0 -3.0 1e-06 
0.05 0.525 0 -3.0 1e-06 
3.0 0.525 0 -3.0 1e-06 
0.05 0.526 0 -3.0 1e-06 
3.0 0.526 0 -3.0 1e-06 
0.05 0.527 0 -3.0 1e-06 
3.0 0.527 0 -3.0 1e-06 
0.05 0.528 0 -3.0 1e-06 
3.0 0.528 0 -3.0 1e-06 
0.05 0.529 0 -3.0 1e-06 
3.0 0.529 0 -3.0 1e-06 
0.05 0.53 0 -3.0 1e-06 
3.0 0.53 0 -3.0 1e-06 
0.05 0.531 0 -3.0 1e-06 
3.0 0.531 0 -3.0 1e-06 
0.05 0.532 0 -3.0 1e-06 
3.0 0.532 0 -3.0 1e-06 
0.05 0.533 0 -3.0 1e-06 
3.0 0.533 0 -3.0 1e-06 
0.05 0.534 0 -3.0 1e-06 
3.0 0.534 0 -3.0 1e-06 
0.05 0.535 0 -3.0 1e-06 
3.0 0.535 0 -3.0 1e-06 
0.05 0.536 0 -3.0 1e-06 
3.0 0.536 0 -3.0 1e-06 
0.05 0.537 0 -3.0 1e-06 
3.0 0.537 0 -3.0 1e-06 
0.05 0.538 0 -3.0 1e-06 
3.0 0.538 0 -3.0 1e-06 
0.05 0.539 0 -3.0 1e-06 
3.0 0.539 0 -3.0 1e-06 
0.05 0.54 0 -3.0 1e-06 
3.0 0.54 0 -3.0 1e-06 
0.05 0.541 0 -3.0 1e-06 
3.0 0.541 0 -3.0 1e-06 
0.05 0.542 0 -3.0 1e-06 
3.0 0.542 0 -3.0 1e-06 
0.05 0.543 0 -3.0 1e-06 
3.0 0.543 0 -3.0 1e-06 
0.05 0.544 0 -3.0 1e-06 
3.0 0.544 0 -3.0 1e-06 
0.05 0.545 0 -3.0 1e-06 
3.0 0.545 0 -3.0 1e-06 
0.05 0.546 0 -3.0 1e-06 
3.0 0.546 0 -3.0 1e-06 
0.05 0.547 0 -3.0 1e-06 
3.0 0.547 0 -3.0 1e-06 
0.05 0.548 0 -3.0 1e-06 
3.0 0.548 0 -3.0 1e-06 
0.05 0.549 0 -3.0 1e-06 
3.0 0.549 0 -3.0 1e-06 
0.05 0.55 0 -3.0 1e-06 
3.0 0.55 0 -3.0 1e-06 
0.05 0.551 0 -3.0 1e-06 
3.0 0.551 0 -3.0 1e-06 
0.05 0.552 0 -3.0 1e-06 
3.0 0.552 0 -3.0 1e-06 
0.05 0.553 0 -3.0 1e-06 
3.0 0.553 0 -3.0 1e-06 
0.05 0.554 0 -3.0 1e-06 
3.0 0.554 0 -3.0 1e-06 
0.05 0.555 0 -3.0 1e-06 
3.0 0.555 0 -3.0 1e-06 
0.05 0.556 0 -3.0 1e-06 
3.0 0.556 0 -3.0 1e-06 
0.05 0.557 0 -3.0 1e-06 
3.0 0.557 0 -3.0 1e-06 
0.05 0.558 0 -3.0 1e-06 
3.0 0.558 0 -3.0 1e-06 
0.05 0.559 0 -3.0 1e-06 
3.0 0.559 0 -3.0 1e-06 
0.05 0.56 0 -3.0 1e-06 
3.0 0.56 0 -3.0 1e-06 
0.05 0.561 0 -3.0 1e-06 
3.0 0.561 0 -3.0 1e-06 
0.05 0.562 0 -3.0 1e-06 
3.0 0.562 0 -3.0 1e-06 
0.05 0.563 0 -3.0 1e-06 
3.0 0.563 0 -3.0 1e-06 
0.05 0.564 0 -3.0 1e-06 
3.0 0.564 0 -3.0 1e-06 
0.05 0.565 0 -3.0 1e-06 
3.0 0.565 0 -3.0 1e-06 
0.05 0.566 0 -3.0 1e-06 
3.0 0.566 0 -3.0 1e-06 
0.05 0.567 0 -3.0 1e-06 
3.0 0.567 0 -3.0 1e-06 
0.05 0.568 0 -3.0 1e-06 
3.0 0.568 0 -3.0 1e-06 
0.05 0.569 0 -3.0 1e-06 
3.0 0.569 0 -3.0 1e-06 
0.05 0.57 0 -3.0 1e-06 
3.0 0.57 0 -3.0 1e-06 
0.05 0.571 0 -3.0 1e-06 
3.0 0.571 0 -3.0 1e-06 
0.05 0.572 0 -3.0 1e-06 
3.0 0.572 0 -3.0 1e-06 
0.05 0.573 0 -3.0 1e-06 
3.0 0.573 0 -3.0 1e-06 
0.05 0.574 0 -3.0 1e-06 
3.0 0.574 0 -3.0 1e-06 
0.05 0.575 0 -3.0 1e-06 
3.0 0.575 0 -3.0 1e-06 
0.05 0.576 0 -3.0 1e-06 
3.0 0.576 0 -3.0 1e-06 
0.05 0.577 0 -3.0 1e-06 
3.0 0.577 0 -3.0 1e-06 
0.05 0.578 0 -3.0 1e-06 
3.0 0.578 0 -3.0 1e-06 
0.05 0.579 0 -3.0 1e-06 
3.0 0.579 0 -3.0 1e-06 
0.05 0.58 0 -3.0 1e-06 
3.0 0.58 0 -3.0 1e-06 
0.05 0.581 0 -3.0 1e-06 
3.0 0.581 0 -3.0 1e-06 
0.05 0.582 0 -3.0 1e-06 
3.0 0.582 0 -3.0 1e-06 
0.05 0.583 0 -3.0 1e-06 
3.0 0.583 0 -3.0 1e-06 
0.05 0.584 0 -3.0 1e-06 
3.0 0.584 0 -3.0 1e-06 
0.05 0.585 0 -3.0 1e-06 
3.0 0.585 0 -3.0 1e-06 
0.05 0.586 0 -3.0 1e-06 
3.0 0.586 0 -3.0 1e-06 
0.05 0.587 0 -3.0 1e-06 
3.0 0.587 0 -3.0 1e-06 
0.05 0.588 0 -3.0 1e-06 
3.0 0.588 0 -3.0 1e-06 
0.05 0.589 0 -3.0 1e-06 
3.0 0.589 0 -3.0 1e-06 
0.05 0.59 0 -3.0 1e-06 
3.0 0.59 0 -3.0 1e-06 
0.05 0.591 0 -3.0 1e-06 
3.0 0.591 0 -3.0 1e-06 
0.05 0.592 0 -3.0 1e-06 
3.0 0.592 0 -3.0 1e-06 
0.05 0.593 0 -3.0 1e-06 
3.0 0.593 0 -3.0 1e-06 
0.05 0.594 0 -3.0 1e-06 
3.0 0.594 0 -3.0 1e-06 
0.05 0.595 0 -3.0 1e-06 
3.0 0.595 0 -3.0 1e-06 
0.05 0.596 0 -3.0 1e-06 
3.0 0.596 0 -3.0 1e-06 
0.05 0.597 0 -3.0 1e-06 
3.0 0.597 0 -3.0 1e-06 
0.05 0.598 0 -3.0 1e-06 
3.0 0.598 0 -3.0 1e-06 
0.05 0.599 0 -3.0 1e-06 
3.0 0.599 0 -3.0 1e-06 
0.05 0.6 0 -3.0 1e-06 
3.0 0.6 0 -3.0 1e-06 
0.05 0.601 0 -3.0 1e-06 
3.0 0.601 0 -3.0 1e-06 
0.05 0.602 0 -3.0 1e-06 
3.0 0.602 0 -3.0 1e-06 
0.05 0.603 0 -3.0 1e-06 
3.0 0.603 0 -3.0 1e-06 
0.05 0.604 0 -3.0 1e-06 
3.0 0.604 0 -3.0 1e-06 
0.05 0.605 0 -3.0 1e-06 
3.0 0.605 0 -3.0 1e-06 
0.05 0.606 0 -3.0 1e-06 
3.0 0.606 0 -3.0 1e-06 
0.05 0.607 0 -3.0 1e-06 
3.0 0.607 0 -3.0 1e-06 
0.05 0.608 0 -3.0 1e-06 
3.0 0.608 0 -3.0 1e-06 
0.05 0.609 0 -3.0 1e-06 
3.0 0.609 0 -3.0 1e-06 
0.05 0.61 0 -3.0 1e-06 
3.0 0.61 0 -3.0 1e-06 
0.05 0.611 0 -3.0 1e-06 
3.0 0.611 0 -3.0 1e-06 
0.05 0.612 0 -3.0 1e-06 
3.0 0.612 0 -3.0 1e-06 
0.05 0.613 0 -3.0 1e-06 
3.0 0.613 0 -3.0 1e-06 
0.05 0.614 0 -3.0 1e-06 
3.0 0.614 0 -3.0 1e-06 
0.05 0.615 0 -3.0 1e-06 
3.0 0.615 0 -3.0 1e-06 
0.05 0.616 0 -3.0 1e-06 
3.0 0.616 0 -3.0 1e-06 
0.05 0.617 0 -3.0 1e-06 
3.0 0.617 0 -3.0 1e-06 
0.05 0.618 0 -3.0 1e-06 
3.0 0.618 0 -3.0 1e-06 
0.05 0.619 0 -3.0 1e-06 
3.0 0.619 0 -3.0 1e-06 
0.05 0.62 0 -3.0 1e-06 
3.0 0.62 0 -3.0 1e-06 
0.05 0.621 0 -3.0 1e-06 
3.0 0.621 0 -3.0 1e-06 
0.05 0.622 0 -3.0 1e-06 
3.0 0.622 0 -3.0 1e-06 
0.05 0.623 0 -3.0 1e-06 
3.0 0.623 0 -3.0 1e-06 
0.05 0.624 0 -3.0 1e-06 
3.0 0.624 0 -3.0 1e-06 
0.05 0.625 0 -3.0 1e-06 
3.0 0.625 0 -3.0 1e-06 
0.05 0.626 0 -3.0 1e-06 
3.0 0.626 0 -3.0 1e-06 
0.05 0.627 0 -3.0 1e-06 
3.0 0.627 0 -3.0 1e-06 
0.05 0.628 0 -3.0 1e-06 
3.0 0.628 0 -3.0 1e-06 
0.05 0.629 0 -3.0 1e-06 
3.0 0.629 0 -3.0 1e-06 
0.05 0.63 0 -3.0 1e-06 
3.0 0.63 0 -3.0 1e-06 
0.05 0.631 0 -3.0 1e-06 
3.0 0.631 0 -3.0 1e-06 
0.05 0.632 0 -3.0 1e-06 
3.0 0.632 0 -3.0 1e-06 
0.05 0.633 0 -3.0 1e-06 
3.0 0.633 0 -3.0 1e-06 
0.05 0.634 0 -3.0 1e-06 
3.0 0.634 0 -3.0 1e-06 
0.05 0.635 0 -3.0 1e-06 
3.0 0.635 0 -3.0 1e-06 
0.05 0.636 0 -3.0 1e-06 
3.0 0.636 0 -3.0 1e-06 
0.05 0.637 0 -3.0 1e-06 
3.0 0.637 0 -3.0 1e-06 
0.05 0.638 0 -3.0 1e-06 
3.0 0.638 0 -3.0 1e-06 
0.05 0.639 0 -3.0 1e-06 
3.0 0.639 0 -3.0 1e-06 
0.05 0.64 0 -3.0 1e-06 
3.0 0.64 0 -3.0 1e-06 
0.05 0.641 0 -3.0 1e-06 
3.0 0.641 0 -3.0 1e-06 
0.05 0.642 0 -3.0 1e-06 
3.0 0.642 0 -3.0 1e-06 
0.05 0.643 0 -3.0 1e-06 
3.0 0.643 0 -3.0 1e-06 
0.05 0.644 0 -3.0 1e-06 
3.0 0.644 0 -3.0 1e-06 
0.05 0.645 0 -3.0 1e-06 
3.0 0.645 0 -3.0 1e-06 
0.05 0.646 0 -3.0 1e-06 
3.0 0.646 0 -3.0 1e-06 
0.05 0.647 0 -3.0 1e-06 
3.0 0.647 0 -3.0 1e-06 
0.05 0.648 0 -3.0 1e-06 
3.0 0.648 0 -3.0 1e-06 
0.05 0.649 0 -3.0 1e-06 
3.0 0.649 0 -3.0 1e-06 
0.05 0.65 0 -3.0 1e-06 
3.0 0.65 0 -3.0 1e-06 
0.05 0.651 0 -3.0 1e-06 
3.0 0.651 0 -3.0 1e-06 
0.05 0.652 0 -3.0 1e-06 
3.0 0.652 0 -3.0 1e-06 
0.05 0.653 0 -3.0 1e-06 
3.0 0.653 0 -3.0 1e-06 
0.05 0.654 0 -3.0 1e-06 
3.0 0.654 0 -3.0 1e-06 
0.05 0.655 0 -3.0 1e-06 
3.0 0.655 0 -3.0 1e-06 
0.05 0.656 0 -3.0 1e-06 
3.0 0.656 0 -3.0 1e-06 
0.05 0.657 0 -3.0 1e-06 
3.0 0.657 0 -3.0 1e-06 
0.05 0.658 0 -3.0 1e-06 
3.0 0.658 0 -3.0 1e-06 
0.05 0.659 0 -3.0 1e-06 
3.0 0.659 0 -3.0 1e-06 
0.05 0.66 0 -3.0 1e-06 
3.0 0.66 0 -3.0 1e-06 
0.05 0.661 0 -3.0 1e-06 
3.0 0.661 0 -3.0 1e-06 
0.05 0.662 0 -3.0 1e-06 
3.0 0.662 0 -3.0 1e-06 
0.05 0.663 0 -3.0 1e-06 
3.0 0.663 0 -3.0 1e-06 
0.05 0.664 0 -3.0 1e-06 
3.0 0.664 0 -3.0 1e-06 
0.05 0.665 0 -3.0 1e-06 
3.0 0.665 0 -3.0 1e-06 
0.05 0.666 0 -3.0 1e-06 
3.0 0.666 0 -3.0 1e-06 
0.05 0.667 0 -3.0 1e-06 
3.0 0.667 0 -3.0 1e-06 
0.05 0.668 0 -3.0 1e-06 
3.0 0.668 0 -3.0 1e-06 
0.05 0.669 0 -3.0 1e-06 
3.0 0.669 0 -3.0 1e-06 
0.05 0.67 0 -3.0 1e-06 
3.0 0.67 0 -3.0 1e-06 
0.05 0.671 0 -3.0 1e-06 
3.0 0.671 0 -3.0 1e-06 
0.05 0.672 0 -3.0 1e-06 
3.0 0.672 0 -3.0 1e-06 
0.05 0.673 0 -3.0 1e-06 
3.0 0.673 0 -3.0 1e-06 
0.05 0.674 0 -3.0 1e-06 
3.0 0.674 0 -3.0 1e-06 
0.05 0.675 0 -3.0 1e-06 
3.0 0.675 0 -3.0 1e-06 
0.05 0.676 0 -3.0 1e-06 
3.0 0.676 0 -3.0 1e-06 
0.05 0.677 0 -3.0 1e-06 
3.0 0.677 0 -3.0 1e-06 
0.05 0.678 0 -3.0 1e-06 
3.0 0.678 0 -3.0 1e-06 
0.05 0.679 0 -3.0 1e-06 
3.0 0.679 0 -3.0 1e-06 
0.05 0.68 0 -3.0 1e-06 
3.0 0.68 0 -3.0 1e-06 
0.05 0.681 0 -3.0 1e-06 
3.0 0.681 0 -3.0 1e-06 
0.05 0.682 0 -3.0 1e-06 
3.0 0.682 0 -3.0 1e-06 
0.05 0.683 0 -3.0 1e-06 
3.0 0.683 0 -3.0 1e-06 
0.05 0.684 0 -3.0 1e-06 
3.0 0.684 0 -3.0 1e-06 
0.05 0.685 0 -3.0 1e-06 
3.0 0.685 0 -3.0 1e-06 
0.05 0.686 0 -3.0 1e-06 
3.0 0.686 0 -3.0 1e-06 
0.05 0.687 0 -3.0 1e-06 
3.0 0.687 0 -3.0 1e-06 
0.05 0.688 0 -3.0 1e-06 
3.0 0.688 0 -3.0 1e-06 
0.05 0.689 0 -3.0 1e-06 
3.0 0.689 0 -3.0 1e-06 
0.05 0.69 0 -3.0 1e-06 
3.0 0.69 0 -3.0 1e-06 
0.05 0.691 0 -3.0 1e-06 
3.0 0.691 0 -3.0 1e-06 
0.05 0.692 0 -3.0 1e-06 
3.0 0.692 0 -3.0 1e-06 
0.05 0.693 0 -3.0 1e-06 
3.0 0.693 0 -3.0 1e-06 
0.05 0.694 0 -3.0 1e-06 
3.0 0.694 0 -3.0 1e-06 
0.05 0.695 0 -3.0 1e-06 
3.0 0.695 0 -3.0 1e-06 
0.05 0.696 0 -3.0 1e-06 
3.0 0.696 0 -3.0 1e-06 
0.05 0.697 0 -3.0 1e-06 
3.0 0.697 0 -3.0 1e-06 
0.05 0.698 0 -3.0 1e-06 
3.0 0.698 0 -3.0 1e-06 
0.05 0.699 0 -3.0 1e-06 
3.0 0.699 0 -3.0 1e-06 
0.05 0.7 0 -3.0 1e-06 
3.0 0.7 0 -3.0 1e-06 
0.05 0.701 0 -3.0 1e-06 
3.0 0.701 0 -3.0 1e-06 
0.05 0.702 0 -3.0 1e-06 
3.0 0.702 0 -3.0 1e-06 
0.05 0.703 0 -3.0 1e-06 
3.0 0.703 0 -3.0 1e-06 
0.05 0.704 0 -3.0 1e-06 
3.0 0.704 0 -3.0 1e-06 
0.05 0.705 0 -3.0 1e-06 
3.0 0.705 0 -3.0 1e-06 
0.05 0.706 0 -3.0 1e-06 
3.0 0.706 0 -3.0 1e-06 
0.05 0.707 0 -3.0 1e-06 
3.0 0.707 0 -3.0 1e-06 
0.05 0.708 0 -3.0 1e-06 
3.0 0.708 0 -3.0 1e-06 
0.05 0.709 0 -3.0 1e-06 
3.0 0.709 0 -3.0 1e-06 
0.05 0.71 0 -3.0 1e-06 
3.0 0.71 0 -3.0 1e-06 
0.05 0.711 0 -3.0 1e-06 
3.0 0.711 0 -3.0 1e-06 
0.05 0.712 0 -3.0 1e-06 
3.0 0.712 0 -3.0 1e-06 
0.05 0.713 0 -3.0 1e-06 
3.0 0.713 0 -3.0 1e-06 
0.05 0.714 0 -3.0 1e-06 
3.0 0.714 0 -3.0 1e-06 
0.05 0.715 0 -3.0 1e-06 
3.0 0.715 0 -3.0 1e-06 
0.05 0.716 0 -3.0 1e-06 
3.0 0.716 0 -3.0 1e-06 
0.05 0.717 0 -3.0 1e-06 
3.0 0.717 0 -3.0 1e-06 
0.05 0.718 0 -3.0 1e-06 
3.0 0.718 0 -3.0 1e-06 
0.05 0.719 0 -3.0 1e-06 
3.0 0.719 0 -3.0 1e-06 
0.05 0.72 0 -3.0 1e-06 
3.0 0.72 0 -3.0 1e-06 
0.05 0.721 0 -3.0 1e-06 
3.0 0.721 0 -3.0 1e-06 
0.05 0.722 0 -3.0 1e-06 
3.0 0.722 0 -3.0 1e-06 
0.05 0.723 0 -3.0 1e-06 
3.0 0.723 0 -3.0 1e-06 
0.05 0.724 0 -3.0 1e-06 
3.0 0.724 0 -3.0 1e-06 
0.05 0.725 0 -3.0 1e-06 
3.0 0.725 0 -3.0 1e-06 
0.05 0.726 0 -3.0 1e-06 
3.0 0.726 0 -3.0 1e-06 
0.05 0.727 0 -3.0 1e-06 
3.0 0.727 0 -3.0 1e-06 
0.05 0.728 0 -3.0 1e-06 
3.0 0.728 0 -3.0 1e-06 
0.05 0.729 0 -3.0 1e-06 
3.0 0.729 0 -3.0 1e-06 
0.05 0.73 0 -3.0 1e-06 
3.0 0.73 0 -3.0 1e-06 
0.05 0.731 0 -3.0 1e-06 
3.0 0.731 0 -3.0 1e-06 
0.05 0.732 0 -3.0 1e-06 
3.0 0.732 0 -3.0 1e-06 
0.05 0.733 0 -3.0 1e-06 
3.0 0.733 0 -3.0 1e-06 
0.05 0.734 0 -3.0 1e-06 
3.0 0.734 0 -3.0 1e-06 
0.05 0.735 0 -3.0 1e-06 
3.0 0.735 0 -3.0 1e-06 
0.05 0.736 0 -3.0 1e-06 
3.0 0.736 0 -3.0 1e-06 
0.05 0.737 0 -3.0 1e-06 
3.0 0.737 0 -3.0 1e-06 
0.05 0.738 0 -3.0 1e-06 
3.0 0.738 0 -3.0 1e-06 
0.05 0.739 0 -3.0 1e-06 
3.0 0.739 0 -3.0 1e-06 
0.05 0.74 0 -3.0 1e-06 
3.0 0.74 0 -3.0 1e-06 
0.05 0.741 0 -3.0 1e-06 
3.0 0.741 0 -3.0 1e-06 
0.05 0.742 0 -3.0 1e-06 
3.0 0.742 0 -3.0 1e-06 
0.05 0.743 0 -3.0 1e-06 
3.0 0.743 0 -3.0 1e-06 
0.05 0.744 0 -3.0 1e-06 
3.0 0.744 0 -3.0 1e-06 
0.05 0.745 0 -3.0 1e-06 
3.0 0.745 0 -3.0 1e-06 
0.05 0.746 0 -3.0 1e-06 
3.0 0.746 0 -3.0 1e-06 
0.05 0.747 0 -3.0 1e-06 
3.0 0.747 0 -3.0 1e-06 
0.05 0.748 0 -3.0 1e-06 
3.0 0.748 0 -3.0 1e-06 
0.05 0.749 0 -3.0 1e-06 
3.0 0.749 0 -3.0 1e-06 
0.05 0.75 0 -3.0 1e-06 
3.0 0.75 0 -3.0 1e-06 
0.05 0.751 0 -3.0 1e-06 
3.0 0.751 0 -3.0 1e-06 
0.05 0.752 0 -3.0 1e-06 
3.0 0.752 0 -3.0 1e-06 
0.05 0.753 0 -3.0 1e-06 
3.0 0.753 0 -3.0 1e-06 
0.05 0.754 0 -3.0 1e-06 
3.0 0.754 0 -3.0 1e-06 
0.05 0.755 0 -3.0 1e-06 
3.0 0.755 0 -3.0 1e-06 
0.05 0.756 0 -3.0 1e-06 
3.0 0.756 0 -3.0 1e-06 
0.05 0.757 0 -3.0 1e-06 
3.0 0.757 0 -3.0 1e-06 
0.05 0.758 0 -3.0 1e-06 
3.0 0.758 0 -3.0 1e-06 
0.05 0.759 0 -3.0 1e-06 
3.0 0.759 0 -3.0 1e-06 
0.05 0.76 0 -3.0 1e-06 
3.0 0.76 0 -3.0 1e-06 
0.05 0.761 0 -3.0 1e-06 
3.0 0.761 0 -3.0 1e-06 
0.05 0.762 0 -3.0 1e-06 
3.0 0.762 0 -3.0 1e-06 
0.05 0.763 0 -3.0 1e-06 
3.0 0.763 0 -3.0 1e-06 
0.05 0.764 0 -3.0 1e-06 
3.0 0.764 0 -3.0 1e-06 
0.05 0.765 0 -3.0 1e-06 
3.0 0.765 0 -3.0 1e-06 
0.05 0.766 0 -3.0 1e-06 
3.0 0.766 0 -3.0 1e-06 
0.05 0.767 0 -3.0 1e-06 
3.0 0.767 0 -3.0 1e-06 
0.05 0.768 0 -3.0 1e-06 
3.0 0.768 0 -3.0 1e-06 
0.05 0.769 0 -3.0 1e-06 
3.0 0.769 0 -3.0 1e-06 
0.05 0.77 0 -3.0 1e-06 
3.0 0.77 0 -3.0 1e-06 
0.05 0.771 0 -3.0 1e-06 
3.0 0.771 0 -3.0 1e-06 
0.05 0.772 0 -3.0 1e-06 
3.0 0.772 0 -3.0 1e-06 
0.05 0.773 0 -3.0 1e-06 
3.0 0.773 0 -3.0 1e-06 
0.05 0.774 0 -3.0 1e-06 
3.0 0.774 0 -3.0 1e-06 
0.05 0.775 0 -3.0 1e-06 
3.0 0.775 0 -3.0 1e-06 
0.05 0.776 0 -3.0 1e-06 
3.0 0.776 0 -3.0 1e-06 
0.05 0.777 0 -3.0 1e-06 
3.0 0.777 0 -3.0 1e-06 
0.05 0.778 0 -3.0 1e-06 
3.0 0.778 0 -3.0 1e-06 
0.05 0.779 0 -3.0 1e-06 
3.0 0.779 0 -3.0 1e-06 
0.05 0.78 0 -3.0 1e-06 
3.0 0.78 0 -3.0 1e-06 
0.05 0.781 0 -3.0 1e-06 
3.0 0.781 0 -3.0 1e-06 
0.05 0.782 0 -3.0 1e-06 
3.0 0.782 0 -3.0 1e-06 
0.05 0.783 0 -3.0 1e-06 
3.0 0.783 0 -3.0 1e-06 
0.05 0.784 0 -3.0 1e-06 
3.0 0.784 0 -3.0 1e-06 
0.05 0.785 0 -3.0 1e-06 
3.0 0.785 0 -3.0 1e-06 
0.05 0.786 0 -3.0 1e-06 
3.0 0.786 0 -3.0 1e-06 
0.05 0.787 0 -3.0 1e-06 
3.0 0.787 0 -3.0 1e-06 
0.05 0.788 0 -3.0 1e-06 
3.0 0.788 0 -3.0 1e-06 
0.05 0.789 0 -3.0 1e-06 
3.0 0.789 0 -3.0 1e-06 
0.05 0.79 0 -3.0 1e-06 
3.0 0.79 0 -3.0 1e-06 
0.05 0.791 0 -3.0 1e-06 
3.0 0.791 0 -3.0 1e-06 
0.05 0.792 0 -3.0 1e-06 
3.0 0.792 0 -3.0 1e-06 
0.05 0.793 0 -3.0 1e-06 
3.0 0.793 0 -3.0 1e-06 
0.05 0.794 0 -3.0 1e-06 
3.0 0.794 0 -3.0 1e-06 
0.05 0.795 0 -3.0 1e-06 
3.0 0.795 0 -3.0 1e-06 
0.05 0.796 0 -3.0 1e-06 
3.0 0.796 0 -3.0 1e-06 
0.05 0.797 0 -3.0 1e-06 
3.0 0.797 0 -3.0 1e-06 
0.05 0.798 0 -3.0 1e-06 
3.0 0.798 0 -3.0 1e-06 
0.05 0.799 0 -3.0 1e-06 
3.0 0.799 0 -3.0 1e-06 
0.05 0.8 0 -3.0 1e-06 
3.0 0.8 0 -3.0 1e-06 
0.05 0.801 0 -3.0 1e-06 
3.0 0.801 0 -3.0 1e-06 
0.05 0.802 0 -3.0 1e-06 
3.0 0.802 0 -3.0 1e-06 
0.05 0.803 0 -3.0 1e-06 
3.0 0.803 0 -3.0 1e-06 
0.05 0.804 0 -3.0 1e-06 
3.0 0.804 0 -3.0 1e-06 
0.05 0.805 0 -3.0 1e-06 
3.0 0.805 0 -3.0 1e-06 
0.05 0.806 0 -3.0 1e-06 
3.0 0.806 0 -3.0 1e-06 
0.05 0.807 0 -3.0 1e-06 
3.0 0.807 0 -3.0 1e-06 
0.05 0.808 0 -3.0 1e-06 
3.0 0.808 0 -3.0 1e-06 
0.05 0.809 0 -3.0 1e-06 
3.0 0.809 0 -3.0 1e-06 
0.05 0.81 0 -3.0 1e-06 
3.0 0.81 0 -3.0 1e-06 
0.05 0.811 0 -3.0 1e-06 
3.0 0.811 0 -3.0 1e-06 
0.05 0.812 0 -3.0 1e-06 
3.0 0.812 0 -3.0 1e-06 
0.05 0.813 0 -3.0 1e-06 
3.0 0.813 0 -3.0 1e-06 
0.05 0.814 0 -3.0 1e-06 
3.0 0.814 0 -3.0 1e-06 
0.05 0.815 0 -3.0 1e-06 
3.0 0.815 0 -3.0 1e-06 
0.05 0.816 0 -3.0 1e-06 
3.0 0.816 0 -3.0 1e-06 
0.05 0.817 0 -3.0 1e-06 
3.0 0.817 0 -3.0 1e-06 
0.05 0.818 0 -3.0 1e-06 
3.0 0.818 0 -3.0 1e-06 
0.05 0.819 0 -3.0 1e-06 
3.0 0.819 0 -3.0 1e-06 
0.05 0.82 0 -3.0 1e-06 
3.0 0.82 0 -3.0 1e-06 
0.05 0.821 0 -3.0 1e-06 
3.0 0.821 0 -3.0 1e-06 
0.05 0.822 0 -3.0 1e-06 
3.0 0.822 0 -3.0 1e-06 
0.05 0.823 0 -3.0 1e-06 
3.0 0.823 0 -3.0 1e-06 
0.05 0.824 0 -3.0 1e-06 
3.0 0.824 0 -3.0 1e-06 
0.05 0.825 0 -3.0 1e-06 
3.0 0.825 0 -3.0 1e-06 
0.05 0.826 0 -3.0 1e-06 
3.0 0.826 0 -3.0 1e-06 
0.05 0.827 0 -3.0 1e-06 
3.0 0.827 0 -3.0 1e-06 
0.05 0.828 0 -3.0 1e-06 
3.0 0.828 0 -3.0 1e-06 
0.05 0.829 0 -3.0 1e-06 
3.0 0.829 0 -3.0 1e-06 
0.05 0.83 0 -3.0 1e-06 
3.0 0.83 0 -3.0 1e-06 
0.05 0.831 0 -3.0 1e-06 
3.0 0.831 0 -3.0 1e-06 
0.05 0.832 0 -3.0 1e-06 
3.0 0.832 0 -3.0 1e-06 
0.05 0.833 0 -3.0 1e-06 
3.0 0.833 0 -3.0 1e-06 
0.05 0.834 0 -3.0 1e-06 
3.0 0.834 0 -3.0 1e-06 
0.05 0.835 0 -3.0 1e-06 
3.0 0.835 0 -3.0 1e-06 
0.05 0.836 0 -3.0 1e-06 
3.0 0.836 0 -3.0 1e-06 
0.05 0.837 0 -3.0 1e-06 
3.0 0.837 0 -3.0 1e-06 
0.05 0.838 0 -3.0 1e-06 
3.0 0.838 0 -3.0 1e-06 
0.05 0.839 0 -3.0 1e-06 
3.0 0.839 0 -3.0 1e-06 
0.05 0.84 0 -3.0 1e-06 
3.0 0.84 0 -3.0 1e-06 
0.05 0.841 0 -3.0 1e-06 
3.0 0.841 0 -3.0 1e-06 
0.05 0.842 0 -3.0 1e-06 
3.0 0.842 0 -3.0 1e-06 
0.05 0.843 0 -3.0 1e-06 
3.0 0.843 0 -3.0 1e-06 
0.05 0.844 0 -3.0 1e-06 
3.0 0.844 0 -3.0 1e-06 
0.05 0.845 0 -3.0 1e-06 
3.0 0.845 0 -3.0 1e-06 
0.05 0.846 0 -3.0 1e-06 
3.0 0.846 0 -3.0 1e-06 
0.05 0.847 0 -3.0 1e-06 
3.0 0.847 0 -3.0 1e-06 
0.05 0.848 0 -3.0 1e-06 
3.0 0.848 0 -3.0 1e-06 
0.05 0.849 0 -3.0 1e-06 
3.0 0.849 0 -3.0 1e-06 
0.05 0.85 0 -3.0 1e-06 
3.0 0.85 0 -3.0 1e-06 
0.05 0.851 0 -3.0 1e-06 
3.0 0.851 0 -3.0 1e-06 
0.05 0.852 0 -3.0 1e-06 
3.0 0.852 0 -3.0 1e-06 
0.05 0.853 0 -3.0 1e-06 
3.0 0.853 0 -3.0 1e-06 
0.05 0.854 0 -3.0 1e-06 
3.0 0.854 0 -3.0 1e-06 
0.05 0.855 0 -3.0 1e-06 
3.0 0.855 0 -3.0 1e-06 
0.05 0.856 0 -3.0 1e-06 
3.0 0.856 0 -3.0 1e-06 
0.05 0.857 0 -3.0 1e-06 
3.0 0.857 0 -3.0 1e-06 
0.05 0.858 0 -3.0 1e-06 
3.0 0.858 0 -3.0 1e-06 
0.05 0.859 0 -3.0 1e-06 
3.0 0.859 0 -3.0 1e-06 
0.05 0.86 0 -3.0 1e-06 
3.0 0.86 0 -3.0 1e-06 
0.05 0.861 0 -3.0 1e-06 
3.0 0.861 0 -3.0 1e-06 
0.05 0.862 0 -3.0 1e-06 
3.0 0.862 0 -3.0 1e-06 
0.05 0.863 0 -3.0 1e-06 
3.0 0.863 0 -3.0 1e-06 
0.05 0.864 0 -3.0 1e-06 
3.0 0.864 0 -3.0 1e-06 
0.05 0.865 0 -3.0 1e-06 
3.0 0.865 0 -3.0 1e-06 
0.05 0.866 0 -3.0 1e-06 
3.0 0.866 0 -3.0 1e-06 
0.05 0.867 0 -3.0 1e-06 
3.0 0.867 0 -3.0 1e-06 
0.05 0.868 0 -3.0 1e-06 
3.0 0.868 0 -3.0 1e-06 
0.05 0.869 0 -3.0 1e-06 
3.0 0.869 0 -3.0 1e-06 
0.05 0.87 0 -3.0 1e-06 
3.0 0.87 0 -3.0 1e-06 
0.05 0.871 0 -3.0 1e-06 
3.0 0.871 0 -3.0 1e-06 
0.05 0.872 0 -3.0 1e-06 
3.0 0.872 0 -3.0 1e-06 
0.05 0.873 0 -3.0 1e-06 
3.0 0.873 0 -3.0 1e-06 
0.05 0.874 0 -3.0 1e-06 
3.0 0.874 0 -3.0 1e-06 
0.05 0.875 0 -3.0 1e-06 
3.0 0.875 0 -3.0 1e-06 
0.05 0.876 0 -3.0 1e-06 
3.0 0.876 0 -3.0 1e-06 
0.05 0.877 0 -3.0 1e-06 
3.0 0.877 0 -3.0 1e-06 
0.05 0.878 0 -3.0 1e-06 
3.0 0.878 0 -3.0 1e-06 
0.05 0.879 0 -3.0 1e-06 
3.0 0.879 0 -3.0 1e-06 
0.05 0.88 0 -3.0 1e-06 
3.0 0.88 0 -3.0 1e-06 
0.05 0.881 0 -3.0 1e-06 
3.0 0.881 0 -3.0 1e-06 
0.05 0.882 0 -3.0 1e-06 
3.0 0.882 0 -3.0 1e-06 
0.05 0.883 0 -3.0 1e-06 
3.0 0.883 0 -3.0 1e-06 
0.05 0.884 0 -3.0 1e-06 
3.0 0.884 0 -3.0 1e-06 
0.05 0.885 0 -3.0 1e-06 
3.0 0.885 0 -3.0 1e-06 
0.05 0.886 0 -3.0 1e-06 
3.0 0.886 0 -3.0 1e-06 
0.05 0.887 0 -3.0 1e-06 
3.0 0.887 0 -3.0 1e-06 
0.05 0.888 0 -3.0 1e-06 
3.0 0.888 0 -3.0 1e-06 
0.05 0.889 0 -3.0 1e-06 
3.0 0.889 0 -3.0 1e-06 
0.05 0.89 0 -3.0 1e-06 
3.0 0.89 0 -3.0 1e-06 
0.05 0.891 0 -3.0 1e-06 
3.0 0.891 0 -3.0 1e-06 
0.05 0.892 0 -3.0 1e-06 
3.0 0.892 0 -3.0 1e-06 
0.05 0.893 0 -3.0 1e-06 
3.0 0.893 0 -3.0 1e-06 
0.05 0.894 0 -3.0 1e-06 
3.0 0.894 0 -3.0 1e-06 
0.05 0.895 0 -3.0 1e-06 
3.0 0.895 0 -3.0 1e-06 
0.05 0.896 0 -3.0 1e-06 
3.0 0.896 0 -3.0 1e-06 
0.05 0.897 0 -3.0 1e-06 
3.0 0.897 0 -3.0 1e-06 
0.05 0.898 0 -3.0 1e-06 
3.0 0.898 0 -3.0 1e-06 
0.05 0.899 0 -3.0 1e-06 
3.0 0.899 0 -3.0 1e-06 
0.05 0.9 0 -3.0 1e-06 
3.0 0.9 0 -3.0 1e-06 
0.05 0.901 0 -3.0 1e-06 
3.0 0.901 0 -3.0 1e-06 
0.05 0.902 0 -3.0 1e-06 
3.0 0.902 0 -3.0 1e-06 
0.05 0.903 0 -3.0 1e-06 
3.0 0.903 0 -3.0 1e-06 
0.05 0.904 0 -3.0 1e-06 
3.0 0.904 0 -3.0 1e-06 
0.05 0.905 0 -3.0 1e-06 
3.0 0.905 0 -3.0 1e-06 
0.05 0.906 0 -3.0 1e-06 
3.0 0.906 0 -3.0 1e-06 
0.05 0.907 0 -3.0 1e-06 
3.0 0.907 0 -3.0 1e-06 
0.05 0.908 0 -3.0 1e-06 
3.0 0.908 0 -3.0 1e-06 
0.05 0.909 0 -3.0 1e-06 
3.0 0.909 0 -3.0 1e-06 
0.05 0.91 0 -3.0 1e-06 
3.0 0.91 0 -3.0 1e-06 
0.05 0.911 0 -3.0 1e-06 
3.0 0.911 0 -3.0 1e-06 
0.05 0.912 0 -3.0 1e-06 
3.0 0.912 0 -3.0 1e-06 
0.05 0.913 0 -3.0 1e-06 
3.0 0.913 0 -3.0 1e-06 
0.05 0.914 0 -3.0 1e-06 
3.0 0.914 0 -3.0 1e-06 
0.05 0.915 0 -3.0 1e-06 
3.0 0.915 0 -3.0 1e-06 
0.05 0.916 0 -3.0 1e-06 
3.0 0.916 0 -3.0 1e-06 
0.05 0.917 0 -3.0 1e-06 
3.0 0.917 0 -3.0 1e-06 
0.05 0.918 0 -3.0 1e-06 
3.0 0.918 0 -3.0 1e-06 
0.05 0.919 0 -3.0 1e-06 
3.0 0.919 0 -3.0 1e-06 
0.05 0.92 0 -3.0 1e-06 
3.0 0.92 0 -3.0 1e-06 
0.05 0.921 0 -3.0 1e-06 
3.0 0.921 0 -3.0 1e-06 
0.05 0.922 0 -3.0 1e-06 
3.0 0.922 0 -3.0 1e-06 
0.05 0.923 0 -3.0 1e-06 
3.0 0.923 0 -3.0 1e-06 
0.05 0.924 0 -3.0 1e-06 
3.0 0.924 0 -3.0 1e-06 
0.05 0.925 0 -3.0 1e-06 
3.0 0.925 0 -3.0 1e-06 
0.05 0.926 0 -3.0 1e-06 
3.0 0.926 0 -3.0 1e-06 
0.05 0.927 0 -3.0 1e-06 
3.0 0.927 0 -3.0 1e-06 
0.05 0.928 0 -3.0 1e-06 
3.0 0.928 0 -3.0 1e-06 
0.05 0.929 0 -3.0 1e-06 
3.0 0.929 0 -3.0 1e-06 
0.05 0.93 0 -3.0 1e-06 
3.0 0.93 0 -3.0 1e-06 
0.05 0.931 0 -3.0 1e-06 
3.0 0.931 0 -3.0 1e-06 
0.05 0.932 0 -3.0 1e-06 
3.0 0.932 0 -3.0 1e-06 
0.05 0.933 0 -3.0 1e-06 
3.0 0.933 0 -3.0 1e-06 
0.05 0.934 0 -3.0 1e-06 
3.0 0.934 0 -3.0 1e-06 
0.05 0.935 0 -3.0 1e-06 
3.0 0.935 0 -3.0 1e-06 
0.05 0.936 0 -3.0 1e-06 
3.0 0.936 0 -3.0 1e-06 
0.05 0.937 0 -3.0 1e-06 
3.0 0.937 0 -3.0 1e-06 
0.05 0.938 0 -3.0 1e-06 
3.0 0.938 0 -3.0 1e-06 
0.05 0.939 0 -3.0 1e-06 
3.0 0.939 0 -3.0 1e-06 
0.05 0.94 0 -3.0 1e-06 
3.0 0.94 0 -3.0 1e-06 
0.05 0.941 0 -3.0 1e-06 
3.0 0.941 0 -3.0 1e-06 
0.05 0.942 0 -3.0 1e-06 
3.0 0.942 0 -3.0 1e-06 
0.05 0.943 0 -3.0 1e-06 
3.0 0.943 0 -3.0 1e-06 
0.05 0.944 0 -3.0 1e-06 
3.0 0.944 0 -3.0 1e-06 
0.05 0.945 0 -3.0 1e-06 
3.0 0.945 0 -3.0 1e-06 
0.05 0.946 0 -3.0 1e-06 
3.0 0.946 0 -3.0 1e-06 
0.05 0.947 0 -3.0 1e-06 
3.0 0.947 0 -3.0 1e-06 
0.05 0.948 0 -3.0 1e-06 
3.0 0.948 0 -3.0 1e-06 
0.05 0.949 0 -3.0 1e-06 
3.0 0.949 0 -3.0 1e-06 
0.05 0.95 0 -3.0 1e-06 
3.0 0.95 0 -3.0 1e-06 
0.05 0.951 0 -3.0 1e-06 
3.0 0.951 0 -3.0 1e-06 
0.05 0.952 0 -3.0 1e-06 
3.0 0.952 0 -3.0 1e-06 
0.05 0.953 0 -3.0 1e-06 
3.0 0.953 0 -3.0 1e-06 
0.05 0.954 0 -3.0 1e-06 
3.0 0.954 0 -3.0 1e-06 
0.05 0.955 0 -3.0 1e-06 
3.0 0.955 0 -3.0 1e-06 
0.05 0.956 0 -3.0 1e-06 
3.0 0.956 0 -3.0 1e-06 
0.05 0.957 0 -3.0 1e-06 
3.0 0.957 0 -3.0 1e-06 
0.05 0.958 0 -3.0 1e-06 
3.0 0.958 0 -3.0 1e-06 
0.05 0.959 0 -3.0 1e-06 
3.0 0.959 0 -3.0 1e-06 
0.05 0.96 0 -3.0 1e-06 
3.0 0.96 0 -3.0 1e-06 
0.05 0.961 0 -3.0 1e-06 
3.0 0.961 0 -3.0 1e-06 
0.05 0.962 0 -3.0 1e-06 
3.0 0.962 0 -3.0 1e-06 
0.05 0.963 0 -3.0 1e-06 
3.0 0.963 0 -3.0 1e-06 
0.05 0.964 0 -3.0 1e-06 
3.0 0.964 0 -3.0 1e-06 
0.05 0.965 0 -3.0 1e-06 
3.0 0.965 0 -3.0 1e-06 
0.05 0.966 0 -3.0 1e-06 
3.0 0.966 0 -3.0 1e-06 
0.05 0.967 0 -3.0 1e-06 
3.0 0.967 0 -3.0 1e-06 
0.05 0.968 0 -3.0 1e-06 
3.0 0.968 0 -3.0 1e-06 
0.05 0.969 0 -3.0 1e-06 
3.0 0.969 0 -3.0 1e-06 
0.05 0.97 0 -3.0 1e-06 
3.0 0.97 0 -3.0 1e-06 
0.05 0.971 0 -3.0 1e-06 
3.0 0.971 0 -3.0 1e-06 
0.05 0.972 0 -3.0 1e-06 
3.0 0.972 0 -3.0 1e-06 
0.05 0.973 0 -3.0 1e-06 
3.0 0.973 0 -3.0 1e-06 
0.05 0.974 0 -3.0 1e-06 
3.0 0.974 0 -3.0 1e-06 
0.05 0.975 0 -3.0 1e-06 
3.0 0.975 0 -3.0 1e-06 
0.05 0.976 0 -3.0 1e-06 
3.0 0.976 0 -3.0 1e-06 
0.05 0.977 0 -3.0 1e-06 
3.0 0.977 0 -3.0 1e-06 
0.05 0.978 0 -3.0 1e-06 
3.0 0.978 0 -3.0 1e-06 
0.05 0.979 0 -3.0 1e-06 
3.0 0.979 0 -3.0 1e-06 
0.05 0.98 0 -3.0 1e-06 
3.0 0.98 0 -3.0 1e-06 
0.05 0.981 0 -3.0 1e-06 
3.0 0.981 0 -3.0 1e-06 
0.05 0.982 0 -3.0 1e-06 
3.0 0.982 0 -3.0 1e-06 
0.05 0.983 0 -3.0 1e-06 
3.0 0.983 0 -3.0 1e-06 
0.05 0.984 0 -3.0 1e-06 
3.0 0.984 0 -3.0 1e-06 
0.05 0.985 0 -3.0 1e-06 
3.0 0.985 0 -3.0 1e-06 
0.05 0.986 0 -3.0 1e-06 
3.0 0.986 0 -3.0 1e-06 
0.05 0.987 0 -3.0 1e-06 
3.0 0.987 0 -3.0 1e-06 
0.05 0.988 0 -3.0 1e-06 
3.0 0.988 0 -3.0 1e-06 
0.05 0.989 0 -3.0 1e-06 
3.0 0.989 0 -3.0 1e-06 
0.05 0.99 0 -3.0 1e-06 
3.0 0.99 0 -3.0 1e-06 
0.05 0.991 0 -3.0 1e-06 
3.0 0.991 0 -3.0 1e-06 
0.05 0.992 0 -3.0 1e-06 
3.0 0.992 0 -3.0 1e-06 
0.05 0.993 0 -3.0 1e-06 
3.0 0.993 0 -3.0 1e-06 
0.05 0.994 0 -3.0 1e-06 
3.0 0.994 0 -3.0 1e-06 
0.05 0.995 0 -3.0 1e-06 
3.0 0.995 0 -3.0 1e-06 
0.05 0.996 0 -3.0 1e-06 
3.0 0.996 0 -3.0 1e-06 
0.05 0.997 0 -3.0 1e-06 
3.0 0.997 0 -3.0 1e-06 
0.05 0.998 0 -3.0 1e-06 
3.0 0.998 0 -3.0 1e-06 
0.05 0.999 0 -3.0 1e-06 
3.0 0.999 0 -3.0 1e-06 
0.05 1.0 0 -3.0 1e-06 
3.0 1.0 0 -3.0 1e-06 
0.05 1.001 0 -3.0 1e-06 
3.0 1.001 0 -3.0 1e-06 
0.05 1.002 0 -3.0 1e-06 
3.0 1.002 0 -3.0 1e-06 
0.05 1.003 0 -3.0 1e-06 
3.0 1.003 0 -3.0 1e-06 
0.05 1.004 0 -3.0 1e-06 
3.0 1.004 0 -3.0 1e-06 
0.05 1.005 0 -3.0 1e-06 
3.0 1.005 0 -3.0 1e-06 
0.05 1.006 0 -3.0 1e-06 
3.0 1.006 0 -3.0 1e-06 
0.05 1.007 0 -3.0 1e-06 
3.0 1.007 0 -3.0 1e-06 
0.05 1.008 0 -3.0 1e-06 
3.0 1.008 0 -3.0 1e-06 
0.05 1.009 0 -3.0 1e-06 
3.0 1.009 0 -3.0 1e-06 
0.05 1.01 0 -3.0 1e-06 
3.0 1.01 0 -3.0 1e-06 
0.05 1.011 0 -3.0 1e-06 
3.0 1.011 0 -3.0 1e-06 
0.05 1.012 0 -3.0 1e-06 
3.0 1.012 0 -3.0 1e-06 
0.05 1.013 0 -3.0 1e-06 
3.0 1.013 0 -3.0 1e-06 
0.05 1.014 0 -3.0 1e-06 
3.0 1.014 0 -3.0 1e-06 
0.05 1.015 0 -3.0 1e-06 
3.0 1.015 0 -3.0 1e-06 
0.05 1.016 0 -3.0 1e-06 
3.0 1.016 0 -3.0 1e-06 
0.05 1.017 0 -3.0 1e-06 
3.0 1.017 0 -3.0 1e-06 
0.05 1.018 0 -3.0 1e-06 
3.0 1.018 0 -3.0 1e-06 
0.05 1.019 0 -3.0 1e-06 
3.0 1.019 0 -3.0 1e-06 
0.05 1.02 0 -3.0 1e-06 
3.0 1.02 0 -3.0 1e-06 
0.05 1.021 0 -3.0 1e-06 
3.0 1.021 0 -3.0 1e-06 
0.05 1.022 0 -3.0 1e-06 
3.0 1.022 0 -3.0 1e-06 
0.05 1.023 0 -3.0 1e-06 
3.0 1.023 0 -3.0 1e-06 
0.05 1.024 0 -3.0 1e-06 
3.0 1.024 0 -3.0 1e-06 
0.05 1.025 0 -3.0 1e-06 
3.0 1.025 0 -3.0 1e-06 
0.05 1.026 0 -3.0 1e-06 
3.0 1.026 0 -3.0 1e-06 
0.05 1.027 0 -3.0 1e-06 
3.0 1.027 0 -3.0 1e-06 
0.05 1.028 0 -3.0 1e-06 
3.0 1.028 0 -3.0 1e-06 
0.05 1.029 0 -3.0 1e-06 
3.0 1.029 0 -3.0 1e-06 
0.05 1.03 0 -3.0 1e-06 
3.0 1.03 0 -3.0 1e-06 
0.05 1.031 0 -3.0 1e-06 
3.0 1.031 0 -3.0 1e-06 
0.05 1.032 0 -3.0 1e-06 
3.0 1.032 0 -3.0 1e-06 
0.05 1.033 0 -3.0 1e-06 
3.0 1.033 0 -3.0 1e-06 
0.05 1.034 0 -3.0 1e-06 
3.0 1.034 0 -3.0 1e-06 
0.05 1.035 0 -3.0 1e-06 
3.0 1.035 0 -3.0 1e-06 
0.05 1.036 0 -3.0 1e-06 
3.0 1.036 0 -3.0 1e-06 
0.05 1.037 0 -3.0 1e-06 
3.0 1.037 0 -3.0 1e-06 
0.05 1.038 0 -3.0 1e-06 
3.0 1.038 0 -3.0 1e-06 
0.05 1.039 0 -3.0 1e-06 
3.0 1.039 0 -3.0 1e-06 
0.05 1.04 0 -3.0 1e-06 
3.0 1.04 0 -3.0 1e-06 
0.05 1.041 0 -3.0 1e-06 
3.0 1.041 0 -3.0 1e-06 
0.05 1.042 0 -3.0 1e-06 
3.0 1.042 0 -3.0 1e-06 
0.05 1.043 0 -3.0 1e-06 
3.0 1.043 0 -3.0 1e-06 
0.05 1.044 0 -3.0 1e-06 
3.0 1.044 0 -3.0 1e-06 
0.05 1.045 0 -3.0 1e-06 
3.0 1.045 0 -3.0 1e-06 
0.05 1.046 0 -3.0 1e-06 
3.0 1.046 0 -3.0 1e-06 
0.05 1.047 0 -3.0 1e-06 
3.0 1.047 0 -3.0 1e-06 
0.05 1.048 0 -3.0 1e-06 
3.0 1.048 0 -3.0 1e-06 
0.05 1.049 0 -3.0 1e-06 
3.0 1.049 0 -3.0 1e-06 
0.05 1.05 0 -3.0 1e-06 
3.0 1.05 0 -3.0 1e-06 
0.05 1.051 0 -3.0 1e-06 
3.0 1.051 0 -3.0 1e-06 
0.05 1.052 0 -3.0 1e-06 
3.0 1.052 0 -3.0 1e-06 
0.05 1.053 0 -3.0 1e-06 
3.0 1.053 0 -3.0 1e-06 
0.05 1.054 0 -3.0 1e-06 
3.0 1.054 0 -3.0 1e-06 
0.05 1.055 0 -3.0 1e-06 
3.0 1.055 0 -3.0 1e-06 
0.05 1.056 0 -3.0 1e-06 
3.0 1.056 0 -3.0 1e-06 
0.05 1.057 0 -3.0 1e-06 
3.0 1.057 0 -3.0 1e-06 
0.05 1.058 0 -3.0 1e-06 
3.0 1.058 0 -3.0 1e-06 
0.05 1.059 0 -3.0 1e-06 
3.0 1.059 0 -3.0 1e-06 
0.05 1.06 0 -3.0 1e-06 
3.0 1.06 0 -3.0 1e-06 
0.05 1.061 0 -3.0 1e-06 
3.0 1.061 0 -3.0 1e-06 
0.05 1.062 0 -3.0 1e-06 
3.0 1.062 0 -3.0 1e-06 
0.05 1.063 0 -3.0 1e-06 
3.0 1.063 0 -3.0 1e-06 
0.05 1.064 0 -3.0 1e-06 
3.0 1.064 0 -3.0 1e-06 
0.05 1.065 0 -3.0 1e-06 
3.0 1.065 0 -3.0 1e-06 
0.05 1.066 0 -3.0 1e-06 
3.0 1.066 0 -3.0 1e-06 
0.05 1.067 0 -3.0 1e-06 
3.0 1.067 0 -3.0 1e-06 
0.05 1.068 0 -3.0 1e-06 
3.0 1.068 0 -3.0 1e-06 
0.05 1.069 0 -3.0 1e-06 
3.0 1.069 0 -3.0 1e-06 
0.05 1.07 0 -3.0 1e-06 
3.0 1.07 0 -3.0 1e-06 
0.05 1.071 0 -3.0 1e-06 
3.0 1.071 0 -3.0 1e-06 
0.05 1.072 0 -3.0 1e-06 
3.0 1.072 0 -3.0 1e-06 
0.05 1.073 0 -3.0 1e-06 
3.0 1.073 0 -3.0 1e-06 
0.05 1.074 0 -3.0 1e-06 
3.0 1.074 0 -3.0 1e-06 
0.05 1.075 0 -3.0 1e-06 
3.0 1.075 0 -3.0 1e-06 
0.05 1.076 0 -3.0 1e-06 
3.0 1.076 0 -3.0 1e-06 
0.05 1.077 0 -3.0 1e-06 
3.0 1.077 0 -3.0 1e-06 
0.05 1.078 0 -3.0 1e-06 
3.0 1.078 0 -3.0 1e-06 
0.05 1.079 0 -3.0 1e-06 
3.0 1.079 0 -3.0 1e-06 
0.05 1.08 0 -3.0 1e-06 
3.0 1.08 0 -3.0 1e-06 
0.05 1.081 0 -3.0 1e-06 
3.0 1.081 0 -3.0 1e-06 
0.05 1.082 0 -3.0 1e-06 
3.0 1.082 0 -3.0 1e-06 
0.05 1.083 0 -3.0 1e-06 
3.0 1.083 0 -3.0 1e-06 
0.05 1.084 0 -3.0 1e-06 
3.0 1.084 0 -3.0 1e-06 
0.05 1.085 0 -3.0 1e-06 
3.0 1.085 0 -3.0 1e-06 
0.05 1.086 0 -3.0 1e-06 
3.0 1.086 0 -3.0 1e-06 
0.05 1.087 0 -3.0 1e-06 
3.0 1.087 0 -3.0 1e-06 
0.05 1.088 0 -3.0 1e-06 
3.0 1.088 0 -3.0 1e-06 
0.05 1.089 0 -3.0 1e-06 
3.0 1.089 0 -3.0 1e-06 
0.05 1.09 0 -3.0 1e-06 
3.0 1.09 0 -3.0 1e-06 
0.05 1.091 0 -3.0 1e-06 
3.0 1.091 0 -3.0 1e-06 
0.05 1.092 0 -3.0 1e-06 
3.0 1.092 0 -3.0 1e-06 
0.05 1.093 0 -3.0 1e-06 
3.0 1.093 0 -3.0 1e-06 
0.05 1.094 0 -3.0 1e-06 
3.0 1.094 0 -3.0 1e-06 
0.05 1.095 0 -3.0 1e-06 
3.0 1.095 0 -3.0 1e-06 
0.05 1.096 0 -3.0 1e-06 
3.0 1.096 0 -3.0 1e-06 
0.05 1.097 0 -3.0 1e-06 
3.0 1.097 0 -3.0 1e-06 
0.05 1.098 0 -3.0 1e-06 
3.0 1.098 0 -3.0 1e-06 
0.05 1.099 0 -3.0 1e-06 
3.0 1.099 0 -3.0 1e-06 
0.05 1.1 0 -3.0 1e-06 
3.0 1.1 0 -3.0 1e-06 
0.05 1.101 0 -3.0 1e-06 
3.0 1.101 0 -3.0 1e-06 
0.05 1.102 0 -3.0 1e-06 
3.0 1.102 0 -3.0 1e-06 
0.05 1.103 0 -3.0 1e-06 
3.0 1.103 0 -3.0 1e-06 
0.05 1.104 0 -3.0 1e-06 
3.0 1.104 0 -3.0 1e-06 
0.05 1.105 0 -3.0 1e-06 
3.0 1.105 0 -3.0 1e-06 
0.05 1.106 0 -3.0 1e-06 
3.0 1.106 0 -3.0 1e-06 
0.05 1.107 0 -3.0 1e-06 
3.0 1.107 0 -3.0 1e-06 
0.05 1.108 0 -3.0 1e-06 
3.0 1.108 0 -3.0 1e-06 
0.05 1.109 0 -3.0 1e-06 
3.0 1.109 0 -3.0 1e-06 
0.05 1.11 0 -3.0 1e-06 
3.0 1.11 0 -3.0 1e-06 
0.05 1.111 0 -3.0 1e-06 
3.0 1.111 0 -3.0 1e-06 
0.05 1.112 0 -3.0 1e-06 
3.0 1.112 0 -3.0 1e-06 
0.05 1.113 0 -3.0 1e-06 
3.0 1.113 0 -3.0 1e-06 
0.05 1.114 0 -3.0 1e-06 
3.0 1.114 0 -3.0 1e-06 
0.05 1.115 0 -3.0 1e-06 
3.0 1.115 0 -3.0 1e-06 
0.05 1.116 0 -3.0 1e-06 
3.0 1.116 0 -3.0 1e-06 
0.05 1.117 0 -3.0 1e-06 
3.0 1.117 0 -3.0 1e-06 
0.05 1.118 0 -3.0 1e-06 
3.0 1.118 0 -3.0 1e-06 
0.05 1.119 0 -3.0 1e-06 
3.0 1.119 0 -3.0 1e-06 
0.05 1.12 0 -3.0 1e-06 
3.0 1.12 0 -3.0 1e-06 
0.05 1.121 0 -3.0 1e-06 
3.0 1.121 0 -3.0 1e-06 
0.05 1.122 0 -3.0 1e-06 
3.0 1.122 0 -3.0 1e-06 
0.05 1.123 0 -3.0 1e-06 
3.0 1.123 0 -3.0 1e-06 
0.05 1.124 0 -3.0 1e-06 
3.0 1.124 0 -3.0 1e-06 
0.05 1.125 0 -3.0 1e-06 
3.0 1.125 0 -3.0 1e-06 
0.05 1.126 0 -3.0 1e-06 
3.0 1.126 0 -3.0 1e-06 
0.05 1.127 0 -3.0 1e-06 
3.0 1.127 0 -3.0 1e-06 
0.05 1.128 0 -3.0 1e-06 
3.0 1.128 0 -3.0 1e-06 
0.05 1.129 0 -3.0 1e-06 
3.0 1.129 0 -3.0 1e-06 
0.05 1.13 0 -3.0 1e-06 
3.0 1.13 0 -3.0 1e-06 
0.05 1.131 0 -3.0 1e-06 
3.0 1.131 0 -3.0 1e-06 
0.05 1.132 0 -3.0 1e-06 
3.0 1.132 0 -3.0 1e-06 
0.05 1.133 0 -3.0 1e-06 
3.0 1.133 0 -3.0 1e-06 
0.05 1.134 0 -3.0 1e-06 
3.0 1.134 0 -3.0 1e-06 
0.05 1.135 0 -3.0 1e-06 
3.0 1.135 0 -3.0 1e-06 
0.05 1.136 0 -3.0 1e-06 
3.0 1.136 0 -3.0 1e-06 
0.05 1.137 0 -3.0 1e-06 
3.0 1.137 0 -3.0 1e-06 
0.05 1.138 0 -3.0 1e-06 
3.0 1.138 0 -3.0 1e-06 
0.05 1.139 0 -3.0 1e-06 
3.0 1.139 0 -3.0 1e-06 
0.05 1.14 0 -3.0 1e-06 
3.0 1.14 0 -3.0 1e-06 
0.05 1.141 0 -3.0 1e-06 
3.0 1.141 0 -3.0 1e-06 
0.05 1.142 0 -3.0 1e-06 
3.0 1.142 0 -3.0 1e-06 
0.05 1.143 0 -3.0 1e-06 
3.0 1.143 0 -3.0 1e-06 
0.05 1.144 0 -3.0 1e-06 
3.0 1.144 0 -3.0 1e-06 
0.05 1.145 0 -3.0 1e-06 
3.0 1.145 0 -3.0 1e-06 
0.05 1.146 0 -3.0 1e-06 
3.0 1.146 0 -3.0 1e-06 
0.05 1.147 0 -3.0 1e-06 
3.0 1.147 0 -3.0 1e-06 
0.05 1.148 0 -3.0 1e-06 
3.0 1.148 0 -3.0 1e-06 
0.05 1.149 0 -3.0 1e-06 
3.0 1.149 0 -3.0 1e-06 
0.05 1.15 0 -3.0 1e-06 
3.0 1.15 0 -3.0 1e-06 
0.05 1.151 0 -3.0 1e-06 
3.0 1.151 0 -3.0 1e-06 
0.05 1.152 0 -3.0 1e-06 
3.0 1.152 0 -3.0 1e-06 
0.05 1.153 0 -3.0 1e-06 
3.0 1.153 0 -3.0 1e-06 
0.05 1.154 0 -3.0 1e-06 
3.0 1.154 0 -3.0 1e-06 
0.05 1.155 0 -3.0 1e-06 
3.0 1.155 0 -3.0 1e-06 
0.05 1.156 0 -3.0 1e-06 
3.0 1.156 0 -3.0 1e-06 
0.05 1.157 0 -3.0 1e-06 
3.0 1.157 0 -3.0 1e-06 
0.05 1.158 0 -3.0 1e-06 
3.0 1.158 0 -3.0 1e-06 
0.05 1.159 0 -3.0 1e-06 
3.0 1.159 0 -3.0 1e-06 
0.05 1.16 0 -3.0 1e-06 
3.0 1.16 0 -3.0 1e-06 
0.05 1.161 0 -3.0 1e-06 
3.0 1.161 0 -3.0 1e-06 
0.05 1.162 0 -3.0 1e-06 
3.0 1.162 0 -3.0 1e-06 
0.05 1.163 0 -3.0 1e-06 
3.0 1.163 0 -3.0 1e-06 
0.05 1.164 0 -3.0 1e-06 
3.0 1.164 0 -3.0 1e-06 
0.05 1.165 0 -3.0 1e-06 
3.0 1.165 0 -3.0 1e-06 
0.05 1.166 0 -3.0 1e-06 
3.0 1.166 0 -3.0 1e-06 
0.05 1.167 0 -3.0 1e-06 
3.0 1.167 0 -3.0 1e-06 
0.05 1.168 0 -3.0 1e-06 
3.0 1.168 0 -3.0 1e-06 
0.05 1.169 0 -3.0 1e-06 
3.0 1.169 0 -3.0 1e-06 
0.05 1.17 0 -3.0 1e-06 
3.0 1.17 0 -3.0 1e-06 
0.05 1.171 0 -3.0 1e-06 
3.0 1.171 0 -3.0 1e-06 
0.05 1.172 0 -3.0 1e-06 
3.0 1.172 0 -3.0 1e-06 
0.05 1.173 0 -3.0 1e-06 
3.0 1.173 0 -3.0 1e-06 
0.05 1.174 0 -3.0 1e-06 
3.0 1.174 0 -3.0 1e-06 
0.05 1.175 0 -3.0 1e-06 
3.0 1.175 0 -3.0 1e-06 
0.05 1.176 0 -3.0 1e-06 
3.0 1.176 0 -3.0 1e-06 
0.05 1.177 0 -3.0 1e-06 
3.0 1.177 0 -3.0 1e-06 
0.05 1.178 0 -3.0 1e-06 
3.0 1.178 0 -3.0 1e-06 
0.05 1.179 0 -3.0 1e-06 
3.0 1.179 0 -3.0 1e-06 
0.05 1.18 0 -3.0 1e-06 
3.0 1.18 0 -3.0 1e-06 
0.05 1.181 0 -3.0 1e-06 
3.0 1.181 0 -3.0 1e-06 
0.05 1.182 0 -3.0 1e-06 
3.0 1.182 0 -3.0 1e-06 
0.05 1.183 0 -3.0 1e-06 
3.0 1.183 0 -3.0 1e-06 
0.05 1.184 0 -3.0 1e-06 
3.0 1.184 0 -3.0 1e-06 
0.05 1.185 0 -3.0 1e-06 
3.0 1.185 0 -3.0 1e-06 
0.05 1.186 0 -3.0 1e-06 
3.0 1.186 0 -3.0 1e-06 
0.05 1.187 0 -3.0 1e-06 
3.0 1.187 0 -3.0 1e-06 
0.05 1.188 0 -3.0 1e-06 
3.0 1.188 0 -3.0 1e-06 
0.05 1.189 0 -3.0 1e-06 
3.0 1.189 0 -3.0 1e-06 
0.05 1.19 0 -3.0 1e-06 
3.0 1.19 0 -3.0 1e-06 
0.05 1.191 0 -3.0 1e-06 
3.0 1.191 0 -3.0 1e-06 
0.05 1.192 0 -3.0 1e-06 
3.0 1.192 0 -3.0 1e-06 
0.05 1.193 0 -3.0 1e-06 
3.0 1.193 0 -3.0 1e-06 
0.05 1.194 0 -3.0 1e-06 
3.0 1.194 0 -3.0 1e-06 
0.05 1.195 0 -3.0 1e-06 
3.0 1.195 0 -3.0 1e-06 
0.05 1.196 0 -3.0 1e-06 
3.0 1.196 0 -3.0 1e-06 
0.05 1.197 0 -3.0 1e-06 
3.0 1.197 0 -3.0 1e-06 
0.05 1.198 0 -3.0 1e-06 
3.0 1.198 0 -3.0 1e-06 
0.05 1.199 0 -3.0 1e-06 
3.0 1.199 0 -3.0 1e-06 
0.05 1.2 0 -3.0 1e-06 
3.0 1.2 0 -3.0 1e-06 
0.05 1.201 0 -3.0 1e-06 
3.0 1.201 0 -3.0 1e-06 
0.05 1.202 0 -3.0 1e-06 
3.0 1.202 0 -3.0 1e-06 
0.05 1.203 0 -3.0 1e-06 
3.0 1.203 0 -3.0 1e-06 
0.05 1.204 0 -3.0 1e-06 
3.0 1.204 0 -3.0 1e-06 
0.05 1.205 0 -3.0 1e-06 
3.0 1.205 0 -3.0 1e-06 
0.05 1.206 0 -3.0 1e-06 
3.0 1.206 0 -3.0 1e-06 
0.05 1.207 0 -3.0 1e-06 
3.0 1.207 0 -3.0 1e-06 
0.05 1.208 0 -3.0 1e-06 
3.0 1.208 0 -3.0 1e-06 
0.05 1.209 0 -3.0 1e-06 
3.0 1.209 0 -3.0 1e-06 
0.05 1.21 0 -3.0 1e-06 
3.0 1.21 0 -3.0 1e-06 
0.05 1.211 0 -3.0 1e-06 
3.0 1.211 0 -3.0 1e-06 
0.05 1.212 0 -3.0 1e-06 
3.0 1.212 0 -3.0 1e-06 
0.05 1.213 0 -3.0 1e-06 
3.0 1.213 0 -3.0 1e-06 
0.05 1.214 0 -3.0 1e-06 
3.0 1.214 0 -3.0 1e-06 
0.05 1.215 0 -3.0 1e-06 
3.0 1.215 0 -3.0 1e-06 
0.05 1.216 0 -3.0 1e-06 
3.0 1.216 0 -3.0 1e-06 
0.05 1.217 0 -3.0 1e-06 
3.0 1.217 0 -3.0 1e-06 
0.05 1.218 0 -3.0 1e-06 
3.0 1.218 0 -3.0 1e-06 
0.05 1.219 0 -3.0 1e-06 
3.0 1.219 0 -3.0 1e-06 
0.05 1.22 0 -3.0 1e-06 
3.0 1.22 0 -3.0 1e-06 
0.05 1.221 0 -3.0 1e-06 
3.0 1.221 0 -3.0 1e-06 
0.05 1.222 0 -3.0 1e-06 
3.0 1.222 0 -3.0 1e-06 
0.05 1.223 0 -3.0 1e-06 
3.0 1.223 0 -3.0 1e-06 
0.05 1.224 0 -3.0 1e-06 
3.0 1.224 0 -3.0 1e-06 
0.05 1.225 0 -3.0 1e-06 
3.0 1.225 0 -3.0 1e-06 
0.05 1.226 0 -3.0 1e-06 
3.0 1.226 0 -3.0 1e-06 
0.05 1.227 0 -3.0 1e-06 
3.0 1.227 0 -3.0 1e-06 
0.05 1.228 0 -3.0 1e-06 
3.0 1.228 0 -3.0 1e-06 
0.05 1.229 0 -3.0 1e-06 
3.0 1.229 0 -3.0 1e-06 
0.05 1.23 0 -3.0 1e-06 
3.0 1.23 0 -3.0 1e-06 
0.05 1.231 0 -3.0 1e-06 
3.0 1.231 0 -3.0 1e-06 
0.05 1.232 0 -3.0 1e-06 
3.0 1.232 0 -3.0 1e-06 
0.05 1.233 0 -3.0 1e-06 
3.0 1.233 0 -3.0 1e-06 
0.05 1.234 0 -3.0 1e-06 
3.0 1.234 0 -3.0 1e-06 
0.05 1.235 0 -3.0 1e-06 
3.0 1.235 0 -3.0 1e-06 
0.05 1.236 0 -3.0 1e-06 
3.0 1.236 0 -3.0 1e-06 
0.05 1.237 0 -3.0 1e-06 
3.0 1.237 0 -3.0 1e-06 
0.05 1.238 0 -3.0 1e-06 
3.0 1.238 0 -3.0 1e-06 
0.05 1.239 0 -3.0 1e-06 
3.0 1.239 0 -3.0 1e-06 
0.05 1.24 0 -3.0 1e-06 
3.0 1.24 0 -3.0 1e-06 
0.05 1.241 0 -3.0 1e-06 
3.0 1.241 0 -3.0 1e-06 
0.05 1.242 0 -3.0 1e-06 
3.0 1.242 0 -3.0 1e-06 
0.05 1.243 0 -3.0 1e-06 
3.0 1.243 0 -3.0 1e-06 
0.05 1.244 0 -3.0 1e-06 
3.0 1.244 0 -3.0 1e-06 
0.05 1.245 0 -3.0 1e-06 
3.0 1.245 0 -3.0 1e-06 
0.05 1.246 0 -3.0 1e-06 
3.0 1.246 0 -3.0 1e-06 
0.05 1.247 0 -3.0 1e-06 
3.0 1.247 0 -3.0 1e-06 
0.05 1.248 0 -3.0 1e-06 
3.0 1.248 0 -3.0 1e-06 
0.05 1.249 0 -3.0 1e-06 
3.0 1.249 0 -3.0 1e-06 
0.05 1.25 0 -3.0 1e-06 
3.0 1.25 0 -3.0 1e-06 
0.05 1.251 0 -3.0 1e-06 
3.0 1.251 0 -3.0 1e-06 
0.05 1.252 0 -3.0 1e-06 
3.0 1.252 0 -3.0 1e-06 
0.05 1.253 0 -3.0 1e-06 
3.0 1.253 0 -3.0 1e-06 
0.05 1.254 0 -3.0 1e-06 
3.0 1.254 0 -3.0 1e-06 
0.05 1.255 0 -3.0 1e-06 
3.0 1.255 0 -3.0 1e-06 
0.05 1.256 0 -3.0 1e-06 
3.0 1.256 0 -3.0 1e-06 
0.05 1.257 0 -3.0 1e-06 
3.0 1.257 0 -3.0 1e-06 
0.05 1.258 0 -3.0 1e-06 
3.0 1.258 0 -3.0 1e-06 
0.05 1.259 0 -3.0 1e-06 
3.0 1.259 0 -3.0 1e-06 
0.05 1.26 0 -3.0 1e-06 
3.0 1.26 0 -3.0 1e-06 
0.05 1.261 0 -3.0 1e-06 
3.0 1.261 0 -3.0 1e-06 
0.05 1.262 0 -3.0 1e-06 
3.0 1.262 0 -3.0 1e-06 
0.05 1.263 0 -3.0 1e-06 
3.0 1.263 0 -3.0 1e-06 
0.05 1.264 0 -3.0 1e-06 
3.0 1.264 0 -3.0 1e-06 
0.05 1.265 0 -3.0 1e-06 
3.0 1.265 0 -3.0 1e-06 
0.05 1.266 0 -3.0 1e-06 
3.0 1.266 0 -3.0 1e-06 
0.05 1.267 0 -3.0 1e-06 
3.0 1.267 0 -3.0 1e-06 
0.05 1.268 0 -3.0 1e-06 
3.0 1.268 0 -3.0 1e-06 
0.05 1.269 0 -3.0 1e-06 
3.0 1.269 0 -3.0 1e-06 
0.05 1.27 0 -3.0 1e-06 
3.0 1.27 0 -3.0 1e-06 
0.05 1.271 0 -3.0 1e-06 
3.0 1.271 0 -3.0 1e-06 
0.05 1.272 0 -3.0 1e-06 
3.0 1.272 0 -3.0 1e-06 
0.05 1.273 0 -3.0 1e-06 
3.0 1.273 0 -3.0 1e-06 
0.05 1.274 0 -3.0 1e-06 
3.0 1.274 0 -3.0 1e-06 
0.05 1.275 0 -3.0 1e-06 
3.0 1.275 0 -3.0 1e-06 
0.05 1.276 0 -3.0 1e-06 
3.0 1.276 0 -3.0 1e-06 
0.05 1.277 0 -3.0 1e-06 
3.0 1.277 0 -3.0 1e-06 
0.05 1.278 0 -3.0 1e-06 
3.0 1.278 0 -3.0 1e-06 
0.05 1.279 0 -3.0 1e-06 
3.0 1.279 0 -3.0 1e-06 
0.05 1.28 0 -3.0 1e-06 
3.0 1.28 0 -3.0 1e-06 
0.05 1.281 0 -3.0 1e-06 
3.0 1.281 0 -3.0 1e-06 
0.05 1.282 0 -3.0 1e-06 
3.0 1.282 0 -3.0 1e-06 
0.05 1.283 0 -3.0 1e-06 
3.0 1.283 0 -3.0 1e-06 
0.05 1.284 0 -3.0 1e-06 
3.0 1.284 0 -3.0 1e-06 
0.05 1.285 0 -3.0 1e-06 
3.0 1.285 0 -3.0 1e-06 
0.05 1.286 0 -3.0 1e-06 
3.0 1.286 0 -3.0 1e-06 
0.05 1.287 0 -3.0 1e-06 
3.0 1.287 0 -3.0 1e-06 
0.05 1.288 0 -3.0 1e-06 
3.0 1.288 0 -3.0 1e-06 
0.05 1.289 0 -3.0 1e-06 
3.0 1.289 0 -3.0 1e-06 
0.05 1.29 0 -3.0 1e-06 
3.0 1.29 0 -3.0 1e-06 
0.05 1.291 0 -3.0 1e-06 
3.0 1.291 0 -3.0 1e-06 
0.05 1.292 0 -3.0 1e-06 
3.0 1.292 0 -3.0 1e-06 
0.05 1.293 0 -3.0 1e-06 
3.0 1.293 0 -3.0 1e-06 
0.05 1.294 0 -3.0 1e-06 
3.0 1.294 0 -3.0 1e-06 
0.05 1.295 0 -3.0 1e-06 
3.0 1.295 0 -3.0 1e-06 
0.05 1.296 0 -3.0 1e-06 
3.0 1.296 0 -3.0 1e-06 
0.05 1.297 0 -3.0 1e-06 
3.0 1.297 0 -3.0 1e-06 
0.05 1.298 0 -3.0 1e-06 
3.0 1.298 0 -3.0 1e-06 
0.05 1.299 0 -3.0 1e-06 
3.0 1.299 0 -3.0 1e-06 
0.05 1.3 0 -3.0 1e-06 
3.0 1.3 0 -3.0 1e-06 
0.05 1.301 0 -3.0 1e-06 
3.0 1.301 0 -3.0 1e-06 
0.05 1.302 0 -3.0 1e-06 
3.0 1.302 0 -3.0 1e-06 
0.05 1.303 0 -3.0 1e-06 
3.0 1.303 0 -3.0 1e-06 
0.05 1.304 0 -3.0 1e-06 
3.0 1.304 0 -3.0 1e-06 
0.05 1.305 0 -3.0 1e-06 
3.0 1.305 0 -3.0 1e-06 
0.05 1.306 0 -3.0 1e-06 
3.0 1.306 0 -3.0 1e-06 
0.05 1.307 0 -3.0 1e-06 
3.0 1.307 0 -3.0 1e-06 
0.05 1.308 0 -3.0 1e-06 
3.0 1.308 0 -3.0 1e-06 
0.05 1.309 0 -3.0 1e-06 
3.0 1.309 0 -3.0 1e-06 
0.05 1.31 0 -3.0 1e-06 
3.0 1.31 0 -3.0 1e-06 
0.05 1.311 0 -3.0 1e-06 
3.0 1.311 0 -3.0 1e-06 
0.05 1.312 0 -3.0 1e-06 
3.0 1.312 0 -3.0 1e-06 
0.05 1.313 0 -3.0 1e-06 
3.0 1.313 0 -3.0 1e-06 
0.05 1.314 0 -3.0 1e-06 
3.0 1.314 0 -3.0 1e-06 
0.05 1.315 0 -3.0 1e-06 
3.0 1.315 0 -3.0 1e-06 
0.05 1.316 0 -3.0 1e-06 
3.0 1.316 0 -3.0 1e-06 
0.05 1.317 0 -3.0 1e-06 
3.0 1.317 0 -3.0 1e-06 
0.05 1.318 0 -3.0 1e-06 
3.0 1.318 0 -3.0 1e-06 
0.05 1.319 0 -3.0 1e-06 
3.0 1.319 0 -3.0 1e-06 
0.05 1.32 0 -3.0 1e-06 
3.0 1.32 0 -3.0 1e-06 
0.05 1.321 0 -3.0 1e-06 
3.0 1.321 0 -3.0 1e-06 
0.05 1.322 0 -3.0 1e-06 
3.0 1.322 0 -3.0 1e-06 
0.05 1.323 0 -3.0 1e-06 
3.0 1.323 0 -3.0 1e-06 
0.05 1.324 0 -3.0 1e-06 
3.0 1.324 0 -3.0 1e-06 
0.05 1.325 0 -3.0 1e-06 
3.0 1.325 0 -3.0 1e-06 
0.05 1.326 0 -3.0 1e-06 
3.0 1.326 0 -3.0 1e-06 
0.05 1.327 0 -3.0 1e-06 
3.0 1.327 0 -3.0 1e-06 
0.05 1.328 0 -3.0 1e-06 
3.0 1.328 0 -3.0 1e-06 
0.05 1.329 0 -3.0 1e-06 
3.0 1.329 0 -3.0 1e-06 
0.05 1.33 0 -3.0 1e-06 
3.0 1.33 0 -3.0 1e-06 
0.05 1.331 0 -3.0 1e-06 
3.0 1.331 0 -3.0 1e-06 
0.05 1.332 0 -3.0 1e-06 
3.0 1.332 0 -3.0 1e-06 
0.05 1.333 0 -3.0 1e-06 
3.0 1.333 0 -3.0 1e-06 
0.05 1.334 0 -3.0 1e-06 
3.0 1.334 0 -3.0 1e-06 
0.05 1.335 0 -3.0 1e-06 
3.0 1.335 0 -3.0 1e-06 
0.05 1.336 0 -3.0 1e-06 
3.0 1.336 0 -3.0 1e-06 
0.05 1.337 0 -3.0 1e-06 
3.0 1.337 0 -3.0 1e-06 
0.05 1.338 0 -3.0 1e-06 
3.0 1.338 0 -3.0 1e-06 
0.05 1.339 0 -3.0 1e-06 
3.0 1.339 0 -3.0 1e-06 
0.05 1.34 0 -3.0 1e-06 
3.0 1.34 0 -3.0 1e-06 
0.05 1.341 0 -3.0 1e-06 
3.0 1.341 0 -3.0 1e-06 
0.05 1.342 0 -3.0 1e-06 
3.0 1.342 0 -3.0 1e-06 
0.05 1.343 0 -3.0 1e-06 
3.0 1.343 0 -3.0 1e-06 
0.05 1.344 0 -3.0 1e-06 
3.0 1.344 0 -3.0 1e-06 
0.05 1.345 0 -3.0 1e-06 
3.0 1.345 0 -3.0 1e-06 
0.05 1.346 0 -3.0 1e-06 
3.0 1.346 0 -3.0 1e-06 
0.05 1.347 0 -3.0 1e-06 
3.0 1.347 0 -3.0 1e-06 
0.05 1.348 0 -3.0 1e-06 
3.0 1.348 0 -3.0 1e-06 
0.05 1.349 0 -3.0 1e-06 
3.0 1.349 0 -3.0 1e-06 
0.05 1.35 0 -3.0 1e-06 
3.0 1.35 0 -3.0 1e-06 
0.05 1.351 0 -3.0 1e-06 
3.0 1.351 0 -3.0 1e-06 
0.05 1.352 0 -3.0 1e-06 
3.0 1.352 0 -3.0 1e-06 
0.05 1.353 0 -3.0 1e-06 
3.0 1.353 0 -3.0 1e-06 
0.05 1.354 0 -3.0 1e-06 
3.0 1.354 0 -3.0 1e-06 
0.05 1.355 0 -3.0 1e-06 
3.0 1.355 0 -3.0 1e-06 
0.05 1.356 0 -3.0 1e-06 
3.0 1.356 0 -3.0 1e-06 
0.05 1.357 0 -3.0 1e-06 
3.0 1.357 0 -3.0 1e-06 
0.05 1.358 0 -3.0 1e-06 
3.0 1.358 0 -3.0 1e-06 
0.05 1.359 0 -3.0 1e-06 
3.0 1.359 0 -3.0 1e-06 
0.05 1.36 0 -3.0 1e-06 
3.0 1.36 0 -3.0 1e-06 
0.05 1.361 0 -3.0 1e-06 
3.0 1.361 0 -3.0 1e-06 
0.05 1.362 0 -3.0 1e-06 
3.0 1.362 0 -3.0 1e-06 
0.05 1.363 0 -3.0 1e-06 
3.0 1.363 0 -3.0 1e-06 
0.05 1.364 0 -3.0 1e-06 
3.0 1.364 0 -3.0 1e-06 
0.05 1.365 0 -3.0 1e-06 
3.0 1.365 0 -3.0 1e-06 
0.05 1.366 0 -3.0 1e-06 
3.0 1.366 0 -3.0 1e-06 
0.05 1.367 0 -3.0 1e-06 
3.0 1.367 0 -3.0 1e-06 
0.05 1.368 0 -3.0 1e-06 
3.0 1.368 0 -3.0 1e-06 
0.05 1.369 0 -3.0 1e-06 
3.0 1.369 0 -3.0 1e-06 
0.05 1.37 0 -3.0 1e-06 
3.0 1.37 0 -3.0 1e-06 
0.05 1.371 0 -3.0 1e-06 
3.0 1.371 0 -3.0 1e-06 
0.05 1.372 0 -3.0 1e-06 
3.0 1.372 0 -3.0 1e-06 
0.05 1.373 0 -3.0 1e-06 
3.0 1.373 0 -3.0 1e-06 
0.05 1.374 0 -3.0 1e-06 
3.0 1.374 0 -3.0 1e-06 
0.05 1.375 0 -3.0 1e-06 
3.0 1.375 0 -3.0 1e-06 
0.05 1.376 0 -3.0 1e-06 
3.0 1.376 0 -3.0 1e-06 
0.05 1.377 0 -3.0 1e-06 
3.0 1.377 0 -3.0 1e-06 
0.05 1.378 0 -3.0 1e-06 
3.0 1.378 0 -3.0 1e-06 
0.05 1.379 0 -3.0 1e-06 
3.0 1.379 0 -3.0 1e-06 
0.05 1.38 0 -3.0 1e-06 
3.0 1.38 0 -3.0 1e-06 
0.05 1.381 0 -3.0 1e-06 
3.0 1.381 0 -3.0 1e-06 
0.05 1.382 0 -3.0 1e-06 
3.0 1.382 0 -3.0 1e-06 
0.05 1.383 0 -3.0 1e-06 
3.0 1.383 0 -3.0 1e-06 
0.05 1.384 0 -3.0 1e-06 
3.0 1.384 0 -3.0 1e-06 
0.05 1.385 0 -3.0 1e-06 
3.0 1.385 0 -3.0 1e-06 
0.05 1.386 0 -3.0 1e-06 
3.0 1.386 0 -3.0 1e-06 
0.05 1.387 0 -3.0 1e-06 
3.0 1.387 0 -3.0 1e-06 
0.05 1.388 0 -3.0 1e-06 
3.0 1.388 0 -3.0 1e-06 
0.05 1.389 0 -3.0 1e-06 
3.0 1.389 0 -3.0 1e-06 
0.05 1.39 0 -3.0 1e-06 
3.0 1.39 0 -3.0 1e-06 
0.05 1.391 0 -3.0 1e-06 
3.0 1.391 0 -3.0 1e-06 
0.05 1.392 0 -3.0 1e-06 
3.0 1.392 0 -3.0 1e-06 
0.05 1.393 0 -3.0 1e-06 
3.0 1.393 0 -3.0 1e-06 
0.05 1.394 0 -3.0 1e-06 
3.0 1.394 0 -3.0 1e-06 
0.05 1.395 0 -3.0 1e-06 
3.0 1.395 0 -3.0 1e-06 
0.05 1.396 0 -3.0 1e-06 
3.0 1.396 0 -3.0 1e-06 
0.05 1.397 0 -3.0 1e-06 
3.0 1.397 0 -3.0 1e-06 
0.05 1.398 0 -3.0 1e-06 
3.0 1.398 0 -3.0 1e-06 
0.05 1.399 0 -3.0 1e-06 
3.0 1.399 0 -3.0 1e-06 
0.05 1.4 0 -3.0 1e-06 
3.0 1.4 0 -3.0 1e-06 
0.05 1.401 0 -3.0 1e-06 
3.0 1.401 0 -3.0 1e-06 
0.05 1.402 0 -3.0 1e-06 
3.0 1.402 0 -3.0 1e-06 
0.05 1.403 0 -3.0 1e-06 
3.0 1.403 0 -3.0 1e-06 
0.05 1.404 0 -3.0 1e-06 
3.0 1.404 0 -3.0 1e-06 
0.05 1.405 0 -3.0 1e-06 
3.0 1.405 0 -3.0 1e-06 
0.05 1.406 0 -3.0 1e-06 
3.0 1.406 0 -3.0 1e-06 
0.05 1.407 0 -3.0 1e-06 
3.0 1.407 0 -3.0 1e-06 
0.05 1.408 0 -3.0 1e-06 
3.0 1.408 0 -3.0 1e-06 
0.05 1.409 0 -3.0 1e-06 
3.0 1.409 0 -3.0 1e-06 
0.05 1.41 0 -3.0 1e-06 
3.0 1.41 0 -3.0 1e-06 
0.05 1.411 0 -3.0 1e-06 
3.0 1.411 0 -3.0 1e-06 
0.05 1.412 0 -3.0 1e-06 
3.0 1.412 0 -3.0 1e-06 
0.05 1.413 0 -3.0 1e-06 
3.0 1.413 0 -3.0 1e-06 
0.05 1.414 0 -3.0 1e-06 
3.0 1.414 0 -3.0 1e-06 
0.05 1.415 0 -3.0 1e-06 
3.0 1.415 0 -3.0 1e-06 
0.05 1.416 0 -3.0 1e-06 
3.0 1.416 0 -3.0 1e-06 
0.05 1.417 0 -3.0 1e-06 
3.0 1.417 0 -3.0 1e-06 
0.05 1.418 0 -3.0 1e-06 
3.0 1.418 0 -3.0 1e-06 
0.05 1.419 0 -3.0 1e-06 
3.0 1.419 0 -3.0 1e-06 
0.05 1.42 0 -3.0 1e-06 
3.0 1.42 0 -3.0 1e-06 
0.05 1.421 0 -3.0 1e-06 
3.0 1.421 0 -3.0 1e-06 
0.05 1.422 0 -3.0 1e-06 
3.0 1.422 0 -3.0 1e-06 
0.05 1.423 0 -3.0 1e-06 
3.0 1.423 0 -3.0 1e-06 
0.05 1.424 0 -3.0 1e-06 
3.0 1.424 0 -3.0 1e-06 
0.05 1.425 0 -3.0 1e-06 
3.0 1.425 0 -3.0 1e-06 
0.05 1.426 0 -3.0 1e-06 
3.0 1.426 0 -3.0 1e-06 
0.05 1.427 0 -3.0 1e-06 
3.0 1.427 0 -3.0 1e-06 
0.05 1.428 0 -3.0 1e-06 
3.0 1.428 0 -3.0 1e-06 
0.05 1.429 0 -3.0 1e-06 
3.0 1.429 0 -3.0 1e-06 
0.05 1.43 0 -3.0 1e-06 
3.0 1.43 0 -3.0 1e-06 
0.05 1.431 0 -3.0 1e-06 
3.0 1.431 0 -3.0 1e-06 
0.05 1.432 0 -3.0 1e-06 
3.0 1.432 0 -3.0 1e-06 
0.05 1.433 0 -3.0 1e-06 
3.0 1.433 0 -3.0 1e-06 
0.05 1.434 0 -3.0 1e-06 
3.0 1.434 0 -3.0 1e-06 
0.05 1.435 0 -3.0 1e-06 
3.0 1.435 0 -3.0 1e-06 
0.05 1.436 0 -3.0 1e-06 
3.0 1.436 0 -3.0 1e-06 
0.05 1.437 0 -3.0 1e-06 
3.0 1.437 0 -3.0 1e-06 
0.05 1.438 0 -3.0 1e-06 
3.0 1.438 0 -3.0 1e-06 
0.05 1.439 0 -3.0 1e-06 
3.0 1.439 0 -3.0 1e-06 
0.05 1.44 0 -3.0 1e-06 
3.0 1.44 0 -3.0 1e-06 
0.05 1.441 0 -3.0 1e-06 
3.0 1.441 0 -3.0 1e-06 
0.05 1.442 0 -3.0 1e-06 
3.0 1.442 0 -3.0 1e-06 
0.05 1.443 0 -3.0 1e-06 
3.0 1.443 0 -3.0 1e-06 
0.05 1.444 0 -3.0 1e-06 
3.0 1.444 0 -3.0 1e-06 
0.05 1.445 0 -3.0 1e-06 
3.0 1.445 0 -3.0 1e-06 
0.05 1.446 0 -3.0 1e-06 
3.0 1.446 0 -3.0 1e-06 
0.05 1.447 0 -3.0 1e-06 
3.0 1.447 0 -3.0 1e-06 
0.05 1.448 0 -3.0 1e-06 
3.0 1.448 0 -3.0 1e-06 
0.05 1.449 0 -3.0 1e-06 
3.0 1.449 0 -3.0 1e-06 
0.05 1.45 0 -3.0 1e-06 
3.0 1.45 0 -3.0 1e-06 
0.05 1.451 0 -3.0 1e-06 
3.0 1.451 0 -3.0 1e-06 
0.05 1.452 0 -3.0 1e-06 
3.0 1.452 0 -3.0 1e-06 
0.05 1.453 0 -3.0 1e-06 
3.0 1.453 0 -3.0 1e-06 
0.05 1.454 0 -3.0 1e-06 
3.0 1.454 0 -3.0 1e-06 
0.05 1.455 0 -3.0 1e-06 
3.0 1.455 0 -3.0 1e-06 
0.05 1.456 0 -3.0 1e-06 
3.0 1.456 0 -3.0 1e-06 
0.05 1.457 0 -3.0 1e-06 
3.0 1.457 0 -3.0 1e-06 
0.05 1.458 0 -3.0 1e-06 
3.0 1.458 0 -3.0 1e-06 
0.05 1.459 0 -3.0 1e-06 
3.0 1.459 0 -3.0 1e-06 
0.05 1.46 0 -3.0 1e-06 
3.0 1.46 0 -3.0 1e-06 
0.05 1.461 0 -3.0 1e-06 
3.0 1.461 0 -3.0 1e-06 
0.05 1.462 0 -3.0 1e-06 
3.0 1.462 0 -3.0 1e-06 
0.05 1.463 0 -3.0 1e-06 
3.0 1.463 0 -3.0 1e-06 
0.05 1.464 0 -3.0 1e-06 
3.0 1.464 0 -3.0 1e-06 
0.05 1.465 0 -3.0 1e-06 
3.0 1.465 0 -3.0 1e-06 
0.05 1.466 0 -3.0 1e-06 
3.0 1.466 0 -3.0 1e-06 
0.05 1.467 0 -3.0 1e-06 
3.0 1.467 0 -3.0 1e-06 
0.05 1.468 0 -3.0 1e-06 
3.0 1.468 0 -3.0 1e-06 
0.05 1.469 0 -3.0 1e-06 
3.0 1.469 0 -3.0 1e-06 
0.05 1.47 0 -3.0 1e-06 
3.0 1.47 0 -3.0 1e-06 
0.05 1.471 0 -3.0 1e-06 
3.0 1.471 0 -3.0 1e-06 
0.05 1.472 0 -3.0 1e-06 
3.0 1.472 0 -3.0 1e-06 
0.05 1.473 0 -3.0 1e-06 
3.0 1.473 0 -3.0 1e-06 
0.05 1.474 0 -3.0 1e-06 
3.0 1.474 0 -3.0 1e-06 
0.05 1.475 0 -3.0 1e-06 
3.0 1.475 0 -3.0 1e-06 
0.05 1.476 0 -3.0 1e-06 
3.0 1.476 0 -3.0 1e-06 
0.05 1.477 0 -3.0 1e-06 
3.0 1.477 0 -3.0 1e-06 
0.05 1.478 0 -3.0 1e-06 
3.0 1.478 0 -3.0 1e-06 
0.05 1.479 0 -3.0 1e-06 
3.0 1.479 0 -3.0 1e-06 
0.05 1.48 0 -3.0 1e-06 
3.0 1.48 0 -3.0 1e-06 
0.05 1.481 0 -3.0 1e-06 
3.0 1.481 0 -3.0 1e-06 
0.05 1.482 0 -3.0 1e-06 
3.0 1.482 0 -3.0 1e-06 
0.05 1.483 0 -3.0 1e-06 
3.0 1.483 0 -3.0 1e-06 
0.05 1.484 0 -3.0 1e-06 
3.0 1.484 0 -3.0 1e-06 
0.05 1.485 0 -3.0 1e-06 
3.0 1.485 0 -3.0 1e-06 
0.05 1.486 0 -3.0 1e-06 
3.0 1.486 0 -3.0 1e-06 
0.05 1.487 0 -3.0 1e-06 
3.0 1.487 0 -3.0 1e-06 
0.05 1.488 0 -3.0 1e-06 
3.0 1.488 0 -3.0 1e-06 
0.05 1.489 0 -3.0 1e-06 
3.0 1.489 0 -3.0 1e-06 
0.05 1.49 0 -3.0 1e-06 
3.0 1.49 0 -3.0 1e-06 
0.05 1.491 0 -3.0 1e-06 
3.0 1.491 0 -3.0 1e-06 
0.05 1.492 0 -3.0 1e-06 
3.0 1.492 0 -3.0 1e-06 
0.05 1.493 0 -3.0 1e-06 
3.0 1.493 0 -3.0 1e-06 
0.05 1.494 0 -3.0 1e-06 
3.0 1.494 0 -3.0 1e-06 
0.05 1.495 0 -3.0 1e-06 
3.0 1.495 0 -3.0 1e-06 
0.05 1.496 0 -3.0 1e-06 
3.0 1.496 0 -3.0 1e-06 
0.05 1.497 0 -3.0 1e-06 
3.0 1.497 0 -3.0 1e-06 
0.05 1.498 0 -3.0 1e-06 
3.0 1.498 0 -3.0 1e-06 
0.05 1.499 0 -3.0 1e-06 
3.0 1.499 0 -3.0 1e-06 
0.05 1.5 0 -3.0 1e-06 
3.0 1.5 0 -3.0 1e-06 
0.05 1.501 0 -3.0 1e-06 
3.0 1.501 0 -3.0 1e-06 
0.05 1.502 0 -3.0 1e-06 
3.0 1.502 0 -3.0 1e-06 
0.05 1.503 0 -3.0 1e-06 
3.0 1.503 0 -3.0 1e-06 
0.05 1.504 0 -3.0 1e-06 
3.0 1.504 0 -3.0 1e-06 
0.05 1.505 0 -3.0 1e-06 
3.0 1.505 0 -3.0 1e-06 
0.05 1.506 0 -3.0 1e-06 
3.0 1.506 0 -3.0 1e-06 
0.05 1.507 0 -3.0 1e-06 
3.0 1.507 0 -3.0 1e-06 
0.05 1.508 0 -3.0 1e-06 
3.0 1.508 0 -3.0 1e-06 
0.05 1.509 0 -3.0 1e-06 
3.0 1.509 0 -3.0 1e-06 
0.05 1.51 0 -3.0 1e-06 
3.0 1.51 0 -3.0 1e-06 
0.05 1.511 0 -3.0 1e-06 
3.0 1.511 0 -3.0 1e-06 
0.05 1.512 0 -3.0 1e-06 
3.0 1.512 0 -3.0 1e-06 
0.05 1.513 0 -3.0 1e-06 
3.0 1.513 0 -3.0 1e-06 
0.05 1.514 0 -3.0 1e-06 
3.0 1.514 0 -3.0 1e-06 
0.05 1.515 0 -3.0 1e-06 
3.0 1.515 0 -3.0 1e-06 
0.05 1.516 0 -3.0 1e-06 
3.0 1.516 0 -3.0 1e-06 
0.05 1.517 0 -3.0 1e-06 
3.0 1.517 0 -3.0 1e-06 
0.05 1.518 0 -3.0 1e-06 
3.0 1.518 0 -3.0 1e-06 
0.05 1.519 0 -3.0 1e-06 
3.0 1.519 0 -3.0 1e-06 
0.05 1.52 0 -3.0 1e-06 
3.0 1.52 0 -3.0 1e-06 
0.05 1.521 0 -3.0 1e-06 
3.0 1.521 0 -3.0 1e-06 
0.05 1.522 0 -3.0 1e-06 
3.0 1.522 0 -3.0 1e-06 
0.05 1.523 0 -3.0 1e-06 
3.0 1.523 0 -3.0 1e-06 
0.05 1.524 0 -3.0 1e-06 
3.0 1.524 0 -3.0 1e-06 
0.05 1.525 0 -3.0 1e-06 
3.0 1.525 0 -3.0 1e-06 
0.05 1.526 0 -3.0 1e-06 
3.0 1.526 0 -3.0 1e-06 
0.05 1.527 0 -3.0 1e-06 
3.0 1.527 0 -3.0 1e-06 
0.05 1.528 0 -3.0 1e-06 
3.0 1.528 0 -3.0 1e-06 
0.05 1.529 0 -3.0 1e-06 
3.0 1.529 0 -3.0 1e-06 
0.05 1.53 0 -3.0 1e-06 
3.0 1.53 0 -3.0 1e-06 
0.05 1.531 0 -3.0 1e-06 
3.0 1.531 0 -3.0 1e-06 
0.05 1.532 0 -3.0 1e-06 
3.0 1.532 0 -3.0 1e-06 
0.05 1.533 0 -3.0 1e-06 
3.0 1.533 0 -3.0 1e-06 
0.05 1.534 0 -3.0 1e-06 
3.0 1.534 0 -3.0 1e-06 
0.05 1.535 0 -3.0 1e-06 
3.0 1.535 0 -3.0 1e-06 
0.05 1.536 0 -3.0 1e-06 
3.0 1.536 0 -3.0 1e-06 
0.05 1.537 0 -3.0 1e-06 
3.0 1.537 0 -3.0 1e-06 
0.05 1.538 0 -3.0 1e-06 
3.0 1.538 0 -3.0 1e-06 
0.05 1.539 0 -3.0 1e-06 
3.0 1.539 0 -3.0 1e-06 
0.05 1.54 0 -3.0 1e-06 
3.0 1.54 0 -3.0 1e-06 
0.05 1.541 0 -3.0 1e-06 
3.0 1.541 0 -3.0 1e-06 
0.05 1.542 0 -3.0 1e-06 
3.0 1.542 0 -3.0 1e-06 
0.05 1.543 0 -3.0 1e-06 
3.0 1.543 0 -3.0 1e-06 
0.05 1.544 0 -3.0 1e-06 
3.0 1.544 0 -3.0 1e-06 
0.05 1.545 0 -3.0 1e-06 
3.0 1.545 0 -3.0 1e-06 
0.05 1.546 0 -3.0 1e-06 
3.0 1.546 0 -3.0 1e-06 
0.05 1.547 0 -3.0 1e-06 
3.0 1.547 0 -3.0 1e-06 
0.05 1.548 0 -3.0 1e-06 
3.0 1.548 0 -3.0 1e-06 
0.05 1.549 0 -3.0 1e-06 
3.0 1.549 0 -3.0 1e-06 
0.05 1.55 0 -3.0 1e-06 
3.0 1.55 0 -3.0 1e-06 
0.05 1.551 0 -3.0 1e-06 
3.0 1.551 0 -3.0 1e-06 
0.05 1.552 0 -3.0 1e-06 
3.0 1.552 0 -3.0 1e-06 
0.05 1.553 0 -3.0 1e-06 
3.0 1.553 0 -3.0 1e-06 
0.05 1.554 0 -3.0 1e-06 
3.0 1.554 0 -3.0 1e-06 
0.05 1.555 0 -3.0 1e-06 
3.0 1.555 0 -3.0 1e-06 
0.05 1.556 0 -3.0 1e-06 
3.0 1.556 0 -3.0 1e-06 
0.05 1.557 0 -3.0 1e-06 
3.0 1.557 0 -3.0 1e-06 
0.05 1.558 0 -3.0 1e-06 
3.0 1.558 0 -3.0 1e-06 
0.05 1.559 0 -3.0 1e-06 
3.0 1.559 0 -3.0 1e-06 
0.05 1.56 0 -3.0 1e-06 
3.0 1.56 0 -3.0 1e-06 
0.05 1.561 0 -3.0 1e-06 
3.0 1.561 0 -3.0 1e-06 
0.05 1.562 0 -3.0 1e-06 
3.0 1.562 0 -3.0 1e-06 
0.05 1.563 0 -3.0 1e-06 
3.0 1.563 0 -3.0 1e-06 
0.05 1.564 0 -3.0 1e-06 
3.0 1.564 0 -3.0 1e-06 
0.05 1.565 0 -3.0 1e-06 
3.0 1.565 0 -3.0 1e-06 
0.05 1.566 0 -3.0 1e-06 
3.0 1.566 0 -3.0 1e-06 
0.05 1.567 0 -3.0 1e-06 
3.0 1.567 0 -3.0 1e-06 
0.05 1.568 0 -3.0 1e-06 
3.0 1.568 0 -3.0 1e-06 
0.05 1.569 0 -3.0 1e-06 
3.0 1.569 0 -3.0 1e-06 
0.05 1.57 0 -3.0 1e-06 
3.0 1.57 0 -3.0 1e-06 
0.05 1.571 0 -3.0 1e-06 
3.0 1.571 0 -3.0 1e-06 
0.05 1.572 0 -3.0 1e-06 
3.0 1.572 0 -3.0 1e-06 
0.05 1.573 0 -3.0 1e-06 
3.0 1.573 0 -3.0 1e-06 
0.05 1.574 0 -3.0 1e-06 
3.0 1.574 0 -3.0 1e-06 
0.05 1.575 0 -3.0 1e-06 
3.0 1.575 0 -3.0 1e-06 
0.05 1.576 0 -3.0 1e-06 
3.0 1.576 0 -3.0 1e-06 
0.05 1.577 0 -3.0 1e-06 
3.0 1.577 0 -3.0 1e-06 
0.05 1.578 0 -3.0 1e-06 
3.0 1.578 0 -3.0 1e-06 
0.05 1.579 0 -3.0 1e-06 
3.0 1.579 0 -3.0 1e-06 
0.05 1.58 0 -3.0 1e-06 
3.0 1.58 0 -3.0 1e-06 
0.05 1.581 0 -3.0 1e-06 
3.0 1.581 0 -3.0 1e-06 
0.05 1.582 0 -3.0 1e-06 
3.0 1.582 0 -3.0 1e-06 
0.05 1.583 0 -3.0 1e-06 
3.0 1.583 0 -3.0 1e-06 
0.05 1.584 0 -3.0 1e-06 
3.0 1.584 0 -3.0 1e-06 
0.05 1.585 0 -3.0 1e-06 
3.0 1.585 0 -3.0 1e-06 
0.05 1.586 0 -3.0 1e-06 
3.0 1.586 0 -3.0 1e-06 
0.05 1.587 0 -3.0 1e-06 
3.0 1.587 0 -3.0 1e-06 
0.05 1.588 0 -3.0 1e-06 
3.0 1.588 0 -3.0 1e-06 
0.05 1.589 0 -3.0 1e-06 
3.0 1.589 0 -3.0 1e-06 
0.05 1.59 0 -3.0 1e-06 
3.0 1.59 0 -3.0 1e-06 
0.05 1.591 0 -3.0 1e-06 
3.0 1.591 0 -3.0 1e-06 
0.05 1.592 0 -3.0 1e-06 
3.0 1.592 0 -3.0 1e-06 
0.05 1.593 0 -3.0 1e-06 
3.0 1.593 0 -3.0 1e-06 
0.05 1.594 0 -3.0 1e-06 
3.0 1.594 0 -3.0 1e-06 
0.05 1.595 0 -3.0 1e-06 
3.0 1.595 0 -3.0 1e-06 
0.05 1.596 0 -3.0 1e-06 
3.0 1.596 0 -3.0 1e-06 
0.05 1.597 0 -3.0 1e-06 
3.0 1.597 0 -3.0 1e-06 
0.05 1.598 0 -3.0 1e-06 
3.0 1.598 0 -3.0 1e-06 
0.05 1.599 0 -3.0 1e-06 
3.0 1.599 0 -3.0 1e-06 
0.05 1.6 0 -3.0 1e-06 
3.0 1.6 0 -3.0 1e-06 
0.05 1.601 0 -3.0 1e-06 
3.0 1.601 0 -3.0 1e-06 
0.05 1.602 0 -3.0 1e-06 
3.0 1.602 0 -3.0 1e-06 
0.05 1.603 0 -3.0 1e-06 
3.0 1.603 0 -3.0 1e-06 
0.05 1.604 0 -3.0 1e-06 
3.0 1.604 0 -3.0 1e-06 
0.05 1.605 0 -3.0 1e-06 
3.0 1.605 0 -3.0 1e-06 
0.05 1.606 0 -3.0 1e-06 
3.0 1.606 0 -3.0 1e-06 
0.05 1.607 0 -3.0 1e-06 
3.0 1.607 0 -3.0 1e-06 
0.05 1.608 0 -3.0 1e-06 
3.0 1.608 0 -3.0 1e-06 
0.05 1.609 0 -3.0 1e-06 
3.0 1.609 0 -3.0 1e-06 
0.05 1.61 0 -3.0 1e-06 
3.0 1.61 0 -3.0 1e-06 
0.05 1.611 0 -3.0 1e-06 
3.0 1.611 0 -3.0 1e-06 
0.05 1.612 0 -3.0 1e-06 
3.0 1.612 0 -3.0 1e-06 
0.05 1.613 0 -3.0 1e-06 
3.0 1.613 0 -3.0 1e-06 
0.05 1.614 0 -3.0 1e-06 
3.0 1.614 0 -3.0 1e-06 
0.05 1.615 0 -3.0 1e-06 
3.0 1.615 0 -3.0 1e-06 
0.05 1.616 0 -3.0 1e-06 
3.0 1.616 0 -3.0 1e-06 
0.05 1.617 0 -3.0 1e-06 
3.0 1.617 0 -3.0 1e-06 
0.05 1.618 0 -3.0 1e-06 
3.0 1.618 0 -3.0 1e-06 
0.05 1.619 0 -3.0 1e-06 
3.0 1.619 0 -3.0 1e-06 
0.05 1.62 0 -3.0 1e-06 
3.0 1.62 0 -3.0 1e-06 
0.05 1.621 0 -3.0 1e-06 
3.0 1.621 0 -3.0 1e-06 
0.05 1.622 0 -3.0 1e-06 
3.0 1.622 0 -3.0 1e-06 
0.05 1.623 0 -3.0 1e-06 
3.0 1.623 0 -3.0 1e-06 
0.05 1.624 0 -3.0 1e-06 
3.0 1.624 0 -3.0 1e-06 
0.05 1.625 0 -3.0 1e-06 
3.0 1.625 0 -3.0 1e-06 
0.05 1.626 0 -3.0 1e-06 
3.0 1.626 0 -3.0 1e-06 
0.05 1.627 0 -3.0 1e-06 
3.0 1.627 0 -3.0 1e-06 
0.05 1.628 0 -3.0 1e-06 
3.0 1.628 0 -3.0 1e-06 
0.05 1.629 0 -3.0 1e-06 
3.0 1.629 0 -3.0 1e-06 
0.05 1.63 0 -3.0 1e-06 
3.0 1.63 0 -3.0 1e-06 
0.05 1.631 0 -3.0 1e-06 
3.0 1.631 0 -3.0 1e-06 
0.05 1.632 0 -3.0 1e-06 
3.0 1.632 0 -3.0 1e-06 
0.05 1.633 0 -3.0 1e-06 
3.0 1.633 0 -3.0 1e-06 
0.05 1.634 0 -3.0 1e-06 
3.0 1.634 0 -3.0 1e-06 
0.05 1.635 0 -3.0 1e-06 
3.0 1.635 0 -3.0 1e-06 
0.05 1.636 0 -3.0 1e-06 
3.0 1.636 0 -3.0 1e-06 
0.05 1.637 0 -3.0 1e-06 
3.0 1.637 0 -3.0 1e-06 
0.05 1.638 0 -3.0 1e-06 
3.0 1.638 0 -3.0 1e-06 
0.05 1.639 0 -3.0 1e-06 
3.0 1.639 0 -3.0 1e-06 
0.05 1.64 0 -3.0 1e-06 
3.0 1.64 0 -3.0 1e-06 
0.05 1.641 0 -3.0 1e-06 
3.0 1.641 0 -3.0 1e-06 
0.05 1.642 0 -3.0 1e-06 
3.0 1.642 0 -3.0 1e-06 
0.05 1.643 0 -3.0 1e-06 
3.0 1.643 0 -3.0 1e-06 
0.05 1.644 0 -3.0 1e-06 
3.0 1.644 0 -3.0 1e-06 
0.05 1.645 0 -3.0 1e-06 
3.0 1.645 0 -3.0 1e-06 
0.05 1.646 0 -3.0 1e-06 
3.0 1.646 0 -3.0 1e-06 
0.05 1.647 0 -3.0 1e-06 
3.0 1.647 0 -3.0 1e-06 
0.05 1.648 0 -3.0 1e-06 
3.0 1.648 0 -3.0 1e-06 
0.05 1.649 0 -3.0 1e-06 
3.0 1.649 0 -3.0 1e-06 
0.05 1.65 0 -3.0 1e-06 
3.0 1.65 0 -3.0 1e-06 
0.05 1.651 0 -3.0 1e-06 
3.0 1.651 0 -3.0 1e-06 
0.05 1.652 0 -3.0 1e-06 
3.0 1.652 0 -3.0 1e-06 
0.05 1.653 0 -3.0 1e-06 
3.0 1.653 0 -3.0 1e-06 
0.05 1.654 0 -3.0 1e-06 
3.0 1.654 0 -3.0 1e-06 
0.05 1.655 0 -3.0 1e-06 
3.0 1.655 0 -3.0 1e-06 
0.05 1.656 0 -3.0 1e-06 
3.0 1.656 0 -3.0 1e-06 
0.05 1.657 0 -3.0 1e-06 
3.0 1.657 0 -3.0 1e-06 
0.05 1.658 0 -3.0 1e-06 
3.0 1.658 0 -3.0 1e-06 
0.05 1.659 0 -3.0 1e-06 
3.0 1.659 0 -3.0 1e-06 
0.05 1.66 0 -3.0 1e-06 
3.0 1.66 0 -3.0 1e-06 
0.05 1.661 0 -3.0 1e-06 
3.0 1.661 0 -3.0 1e-06 
0.05 1.662 0 -3.0 1e-06 
3.0 1.662 0 -3.0 1e-06 
0.05 1.663 0 -3.0 1e-06 
3.0 1.663 0 -3.0 1e-06 
0.05 1.664 0 -3.0 1e-06 
3.0 1.664 0 -3.0 1e-06 
0.05 1.665 0 -3.0 1e-06 
3.0 1.665 0 -3.0 1e-06 
0.05 1.666 0 -3.0 1e-06 
3.0 1.666 0 -3.0 1e-06 
0.05 1.667 0 -3.0 1e-06 
3.0 1.667 0 -3.0 1e-06 
0.05 1.668 0 -3.0 1e-06 
3.0 1.668 0 -3.0 1e-06 
0.05 1.669 0 -3.0 1e-06 
3.0 1.669 0 -3.0 1e-06 
0.05 1.67 0 -3.0 1e-06 
3.0 1.67 0 -3.0 1e-06 
0.05 1.671 0 -3.0 1e-06 
3.0 1.671 0 -3.0 1e-06 
0.05 1.672 0 -3.0 1e-06 
3.0 1.672 0 -3.0 1e-06 
0.05 1.673 0 -3.0 1e-06 
3.0 1.673 0 -3.0 1e-06 
0.05 1.674 0 -3.0 1e-06 
3.0 1.674 0 -3.0 1e-06 
0.05 1.675 0 -3.0 1e-06 
3.0 1.675 0 -3.0 1e-06 
0.05 1.676 0 -3.0 1e-06 
3.0 1.676 0 -3.0 1e-06 
0.05 1.677 0 -3.0 1e-06 
3.0 1.677 0 -3.0 1e-06 
0.05 1.678 0 -3.0 1e-06 
3.0 1.678 0 -3.0 1e-06 
0.05 1.679 0 -3.0 1e-06 
3.0 1.679 0 -3.0 1e-06 
0.05 1.68 0 -3.0 1e-06 
3.0 1.68 0 -3.0 1e-06 
0.05 1.681 0 -3.0 1e-06 
3.0 1.681 0 -3.0 1e-06 
0.05 1.682 0 -3.0 1e-06 
3.0 1.682 0 -3.0 1e-06 
0.05 1.683 0 -3.0 1e-06 
3.0 1.683 0 -3.0 1e-06 
0.05 1.684 0 -3.0 1e-06 
3.0 1.684 0 -3.0 1e-06 
0.05 1.685 0 -3.0 1e-06 
3.0 1.685 0 -3.0 1e-06 
0.05 1.686 0 -3.0 1e-06 
3.0 1.686 0 -3.0 1e-06 
0.05 1.687 0 -3.0 1e-06 
3.0 1.687 0 -3.0 1e-06 
0.05 1.688 0 -3.0 1e-06 
3.0 1.688 0 -3.0 1e-06 
0.05 1.689 0 -3.0 1e-06 
3.0 1.689 0 -3.0 1e-06 
0.05 1.69 0 -3.0 1e-06 
3.0 1.69 0 -3.0 1e-06 
0.05 1.691 0 -3.0 1e-06 
3.0 1.691 0 -3.0 1e-06 
0.05 1.692 0 -3.0 1e-06 
3.0 1.692 0 -3.0 1e-06 
0.05 1.693 0 -3.0 1e-06 
3.0 1.693 0 -3.0 1e-06 
0.05 1.694 0 -3.0 1e-06 
3.0 1.694 0 -3.0 1e-06 
0.05 1.695 0 -3.0 1e-06 
3.0 1.695 0 -3.0 1e-06 
0.05 1.696 0 -3.0 1e-06 
3.0 1.696 0 -3.0 1e-06 
0.05 1.697 0 -3.0 1e-06 
3.0 1.697 0 -3.0 1e-06 
0.05 1.698 0 -3.0 1e-06 
3.0 1.698 0 -3.0 1e-06 
0.05 1.699 0 -3.0 1e-06 
3.0 1.699 0 -3.0 1e-06 
0.05 1.7 0 -3.0 1e-06 
3.0 1.7 0 -3.0 1e-06 
0.05 1.701 0 -3.0 1e-06 
3.0 1.701 0 -3.0 1e-06 
0.05 1.702 0 -3.0 1e-06 
3.0 1.702 0 -3.0 1e-06 
0.05 1.703 0 -3.0 1e-06 
3.0 1.703 0 -3.0 1e-06 
0.05 1.704 0 -3.0 1e-06 
3.0 1.704 0 -3.0 1e-06 
0.05 1.705 0 -3.0 1e-06 
3.0 1.705 0 -3.0 1e-06 
0.05 1.706 0 -3.0 1e-06 
3.0 1.706 0 -3.0 1e-06 
0.05 1.707 0 -3.0 1e-06 
3.0 1.707 0 -3.0 1e-06 
0.05 1.708 0 -3.0 1e-06 
3.0 1.708 0 -3.0 1e-06 
0.05 1.709 0 -3.0 1e-06 
3.0 1.709 0 -3.0 1e-06 
0.05 1.71 0 -3.0 1e-06 
3.0 1.71 0 -3.0 1e-06 
0.05 1.711 0 -3.0 1e-06 
3.0 1.711 0 -3.0 1e-06 
0.05 1.712 0 -3.0 1e-06 
3.0 1.712 0 -3.0 1e-06 
0.05 1.713 0 -3.0 1e-06 
3.0 1.713 0 -3.0 1e-06 
0.05 1.714 0 -3.0 1e-06 
3.0 1.714 0 -3.0 1e-06 
0.05 1.715 0 -3.0 1e-06 
3.0 1.715 0 -3.0 1e-06 
0.05 1.716 0 -3.0 1e-06 
3.0 1.716 0 -3.0 1e-06 
0.05 1.717 0 -3.0 1e-06 
3.0 1.717 0 -3.0 1e-06 
0.05 1.718 0 -3.0 1e-06 
3.0 1.718 0 -3.0 1e-06 
0.05 1.719 0 -3.0 1e-06 
3.0 1.719 0 -3.0 1e-06 
0.05 1.72 0 -3.0 1e-06 
3.0 1.72 0 -3.0 1e-06 
0.05 1.721 0 -3.0 1e-06 
3.0 1.721 0 -3.0 1e-06 
0.05 1.722 0 -3.0 1e-06 
3.0 1.722 0 -3.0 1e-06 
0.05 1.723 0 -3.0 1e-06 
3.0 1.723 0 -3.0 1e-06 
0.05 1.724 0 -3.0 1e-06 
3.0 1.724 0 -3.0 1e-06 
0.05 1.725 0 -3.0 1e-06 
3.0 1.725 0 -3.0 1e-06 
0.05 1.726 0 -3.0 1e-06 
3.0 1.726 0 -3.0 1e-06 
0.05 1.727 0 -3.0 1e-06 
3.0 1.727 0 -3.0 1e-06 
0.05 1.728 0 -3.0 1e-06 
3.0 1.728 0 -3.0 1e-06 
0.05 1.729 0 -3.0 1e-06 
3.0 1.729 0 -3.0 1e-06 
0.05 1.73 0 -3.0 1e-06 
3.0 1.73 0 -3.0 1e-06 
0.05 1.731 0 -3.0 1e-06 
3.0 1.731 0 -3.0 1e-06 
0.05 1.732 0 -3.0 1e-06 
3.0 1.732 0 -3.0 1e-06 
0.05 1.733 0 -3.0 1e-06 
3.0 1.733 0 -3.0 1e-06 
0.05 1.734 0 -3.0 1e-06 
3.0 1.734 0 -3.0 1e-06 
0.05 1.735 0 -3.0 1e-06 
3.0 1.735 0 -3.0 1e-06 
0.05 1.736 0 -3.0 1e-06 
3.0 1.736 0 -3.0 1e-06 
0.05 1.737 0 -3.0 1e-06 
3.0 1.737 0 -3.0 1e-06 
0.05 1.738 0 -3.0 1e-06 
3.0 1.738 0 -3.0 1e-06 
0.05 1.739 0 -3.0 1e-06 
3.0 1.739 0 -3.0 1e-06 
0.05 1.74 0 -3.0 1e-06 
3.0 1.74 0 -3.0 1e-06 
0.05 1.741 0 -3.0 1e-06 
3.0 1.741 0 -3.0 1e-06 
0.05 1.742 0 -3.0 1e-06 
3.0 1.742 0 -3.0 1e-06 
0.05 1.743 0 -3.0 1e-06 
3.0 1.743 0 -3.0 1e-06 
0.05 1.744 0 -3.0 1e-06 
3.0 1.744 0 -3.0 1e-06 
0.05 1.745 0 -3.0 1e-06 
3.0 1.745 0 -3.0 1e-06 
0.05 1.746 0 -3.0 1e-06 
3.0 1.746 0 -3.0 1e-06 
0.05 1.747 0 -3.0 1e-06 
3.0 1.747 0 -3.0 1e-06 
0.05 1.748 0 -3.0 1e-06 
3.0 1.748 0 -3.0 1e-06 
0.05 1.749 0 -3.0 1e-06 
3.0 1.749 0 -3.0 1e-06 
0.05 1.75 0 -3.0 1e-06 
3.0 1.75 0 -3.0 1e-06 
0.05 1.751 0 -3.0 1e-06 
3.0 1.751 0 -3.0 1e-06 
0.05 1.752 0 -3.0 1e-06 
3.0 1.752 0 -3.0 1e-06 
0.05 1.753 0 -3.0 1e-06 
3.0 1.753 0 -3.0 1e-06 
0.05 1.754 0 -3.0 1e-06 
3.0 1.754 0 -3.0 1e-06 
0.05 1.755 0 -3.0 1e-06 
3.0 1.755 0 -3.0 1e-06 
0.05 1.756 0 -3.0 1e-06 
3.0 1.756 0 -3.0 1e-06 
0.05 1.757 0 -3.0 1e-06 
3.0 1.757 0 -3.0 1e-06 
0.05 1.758 0 -3.0 1e-06 
3.0 1.758 0 -3.0 1e-06 
0.05 1.759 0 -3.0 1e-06 
3.0 1.759 0 -3.0 1e-06 
0.05 1.76 0 -3.0 1e-06 
3.0 1.76 0 -3.0 1e-06 
0.05 1.761 0 -3.0 1e-06 
3.0 1.761 0 -3.0 1e-06 
0.05 1.762 0 -3.0 1e-06 
3.0 1.762 0 -3.0 1e-06 
0.05 1.763 0 -3.0 1e-06 
3.0 1.763 0 -3.0 1e-06 
0.05 1.764 0 -3.0 1e-06 
3.0 1.764 0 -3.0 1e-06 
0.05 1.765 0 -3.0 1e-06 
3.0 1.765 0 -3.0 1e-06 
0.05 1.766 0 -3.0 1e-06 
3.0 1.766 0 -3.0 1e-06 
0.05 1.767 0 -3.0 1e-06 
3.0 1.767 0 -3.0 1e-06 
0.05 1.768 0 -3.0 1e-06 
3.0 1.768 0 -3.0 1e-06 
0.05 1.769 0 -3.0 1e-06 
3.0 1.769 0 -3.0 1e-06 
0.05 1.77 0 -3.0 1e-06 
3.0 1.77 0 -3.0 1e-06 
0.05 1.771 0 -3.0 1e-06 
3.0 1.771 0 -3.0 1e-06 
0.05 1.772 0 -3.0 1e-06 
3.0 1.772 0 -3.0 1e-06 
0.05 1.773 0 -3.0 1e-06 
3.0 1.773 0 -3.0 1e-06 
0.05 1.774 0 -3.0 1e-06 
3.0 1.774 0 -3.0 1e-06 
0.05 1.775 0 -3.0 1e-06 
3.0 1.775 0 -3.0 1e-06 
0.05 1.776 0 -3.0 1e-06 
3.0 1.776 0 -3.0 1e-06 
0.05 1.777 0 -3.0 1e-06 
3.0 1.777 0 -3.0 1e-06 
0.05 1.778 0 -3.0 1e-06 
3.0 1.778 0 -3.0 1e-06 
0.05 1.779 0 -3.0 1e-06 
3.0 1.779 0 -3.0 1e-06 
0.05 1.78 0 -3.0 1e-06 
3.0 1.78 0 -3.0 1e-06 
0.05 1.781 0 -3.0 1e-06 
3.0 1.781 0 -3.0 1e-06 
0.05 1.782 0 -3.0 1e-06 
3.0 1.782 0 -3.0 1e-06 
0.05 1.783 0 -3.0 1e-06 
3.0 1.783 0 -3.0 1e-06 
0.05 1.784 0 -3.0 1e-06 
3.0 1.784 0 -3.0 1e-06 
0.05 1.785 0 -3.0 1e-06 
3.0 1.785 0 -3.0 1e-06 
0.05 1.786 0 -3.0 1e-06 
3.0 1.786 0 -3.0 1e-06 
0.05 1.787 0 -3.0 1e-06 
3.0 1.787 0 -3.0 1e-06 
0.05 1.788 0 -3.0 1e-06 
3.0 1.788 0 -3.0 1e-06 
0.05 1.789 0 -3.0 1e-06 
3.0 1.789 0 -3.0 1e-06 
0.05 1.79 0 -3.0 1e-06 
3.0 1.79 0 -3.0 1e-06 
0.05 1.791 0 -3.0 1e-06 
3.0 1.791 0 -3.0 1e-06 
0.05 1.792 0 -3.0 1e-06 
3.0 1.792 0 -3.0 1e-06 
0.05 1.793 0 -3.0 1e-06 
3.0 1.793 0 -3.0 1e-06 
0.05 1.794 0 -3.0 1e-06 
3.0 1.794 0 -3.0 1e-06 
0.05 1.795 0 -3.0 1e-06 
3.0 1.795 0 -3.0 1e-06 
0.05 1.796 0 -3.0 1e-06 
3.0 1.796 0 -3.0 1e-06 
0.05 1.797 0 -3.0 1e-06 
3.0 1.797 0 -3.0 1e-06 
0.05 1.798 0 -3.0 1e-06 
3.0 1.798 0 -3.0 1e-06 
0.05 1.799 0 -3.0 1e-06 
3.0 1.799 0 -3.0 1e-06 
0.05 1.8 0 -3.0 1e-06 
3.0 1.8 0 -3.0 1e-06 
0.05 1.801 0 -3.0 1e-06 
3.0 1.801 0 -3.0 1e-06 
0.05 1.802 0 -3.0 1e-06 
3.0 1.802 0 -3.0 1e-06 
0.05 1.803 0 -3.0 1e-06 
3.0 1.803 0 -3.0 1e-06 
0.05 1.804 0 -3.0 1e-06 
3.0 1.804 0 -3.0 1e-06 
0.05 1.805 0 -3.0 1e-06 
3.0 1.805 0 -3.0 1e-06 
0.05 1.806 0 -3.0 1e-06 
3.0 1.806 0 -3.0 1e-06 
0.05 1.807 0 -3.0 1e-06 
3.0 1.807 0 -3.0 1e-06 
0.05 1.808 0 -3.0 1e-06 
3.0 1.808 0 -3.0 1e-06 
0.05 1.809 0 -3.0 1e-06 
3.0 1.809 0 -3.0 1e-06 
0.05 1.81 0 -3.0 1e-06 
3.0 1.81 0 -3.0 1e-06 
0.05 1.811 0 -3.0 1e-06 
3.0 1.811 0 -3.0 1e-06 
0.05 1.812 0 -3.0 1e-06 
3.0 1.812 0 -3.0 1e-06 
0.05 1.813 0 -3.0 1e-06 
3.0 1.813 0 -3.0 1e-06 
0.05 1.814 0 -3.0 1e-06 
3.0 1.814 0 -3.0 1e-06 
0.05 1.815 0 -3.0 1e-06 
3.0 1.815 0 -3.0 1e-06 
0.05 1.816 0 -3.0 1e-06 
3.0 1.816 0 -3.0 1e-06 
0.05 1.817 0 -3.0 1e-06 
3.0 1.817 0 -3.0 1e-06 
0.05 1.818 0 -3.0 1e-06 
3.0 1.818 0 -3.0 1e-06 
0.05 1.819 0 -3.0 1e-06 
3.0 1.819 0 -3.0 1e-06 
0.05 1.82 0 -3.0 1e-06 
3.0 1.82 0 -3.0 1e-06 
0.05 1.821 0 -3.0 1e-06 
3.0 1.821 0 -3.0 1e-06 
0.05 1.822 0 -3.0 1e-06 
3.0 1.822 0 -3.0 1e-06 
0.05 1.823 0 -3.0 1e-06 
3.0 1.823 0 -3.0 1e-06 
0.05 1.824 0 -3.0 1e-06 
3.0 1.824 0 -3.0 1e-06 
0.05 1.825 0 -3.0 1e-06 
3.0 1.825 0 -3.0 1e-06 
0.05 1.826 0 -3.0 1e-06 
3.0 1.826 0 -3.0 1e-06 
0.05 1.827 0 -3.0 1e-06 
3.0 1.827 0 -3.0 1e-06 
0.05 1.828 0 -3.0 1e-06 
3.0 1.828 0 -3.0 1e-06 
0.05 1.829 0 -3.0 1e-06 
3.0 1.829 0 -3.0 1e-06 
0.05 1.83 0 -3.0 1e-06 
3.0 1.83 0 -3.0 1e-06 
0.05 1.831 0 -3.0 1e-06 
3.0 1.831 0 -3.0 1e-06 
0.05 1.832 0 -3.0 1e-06 
3.0 1.832 0 -3.0 1e-06 
0.05 1.833 0 -3.0 1e-06 
3.0 1.833 0 -3.0 1e-06 
0.05 1.834 0 -3.0 1e-06 
3.0 1.834 0 -3.0 1e-06 
0.05 1.835 0 -3.0 1e-06 
3.0 1.835 0 -3.0 1e-06 
0.05 1.836 0 -3.0 1e-06 
3.0 1.836 0 -3.0 1e-06 
0.05 1.837 0 -3.0 1e-06 
3.0 1.837 0 -3.0 1e-06 
0.05 1.838 0 -3.0 1e-06 
3.0 1.838 0 -3.0 1e-06 
0.05 1.839 0 -3.0 1e-06 
3.0 1.839 0 -3.0 1e-06 
0.05 1.84 0 -3.0 1e-06 
3.0 1.84 0 -3.0 1e-06 
0.05 1.841 0 -3.0 1e-06 
3.0 1.841 0 -3.0 1e-06 
0.05 1.842 0 -3.0 1e-06 
3.0 1.842 0 -3.0 1e-06 
0.05 1.843 0 -3.0 1e-06 
3.0 1.843 0 -3.0 1e-06 
0.05 1.844 0 -3.0 1e-06 
3.0 1.844 0 -3.0 1e-06 
0.05 1.845 0 -3.0 1e-06 
3.0 1.845 0 -3.0 1e-06 
0.05 1.846 0 -3.0 1e-06 
3.0 1.846 0 -3.0 1e-06 
0.05 1.847 0 -3.0 1e-06 
3.0 1.847 0 -3.0 1e-06 
0.05 1.848 0 -3.0 1e-06 
3.0 1.848 0 -3.0 1e-06 
0.05 1.849 0 -3.0 1e-06 
3.0 1.849 0 -3.0 1e-06 
0.05 1.85 0 -3.0 1e-06 
3.0 1.85 0 -3.0 1e-06 
0.05 1.851 0 -3.0 1e-06 
3.0 1.851 0 -3.0 1e-06 
0.05 1.852 0 -3.0 1e-06 
3.0 1.852 0 -3.0 1e-06 
0.05 1.853 0 -3.0 1e-06 
3.0 1.853 0 -3.0 1e-06 
0.05 1.854 0 -3.0 1e-06 
3.0 1.854 0 -3.0 1e-06 
0.05 1.855 0 -3.0 1e-06 
3.0 1.855 0 -3.0 1e-06 
0.05 1.856 0 -3.0 1e-06 
3.0 1.856 0 -3.0 1e-06 
0.05 1.857 0 -3.0 1e-06 
3.0 1.857 0 -3.0 1e-06 
0.05 1.858 0 -3.0 1e-06 
3.0 1.858 0 -3.0 1e-06 
0.05 1.859 0 -3.0 1e-06 
3.0 1.859 0 -3.0 1e-06 
0.05 1.86 0 -3.0 1e-06 
3.0 1.86 0 -3.0 1e-06 
0.05 1.861 0 -3.0 1e-06 
3.0 1.861 0 -3.0 1e-06 
0.05 1.862 0 -3.0 1e-06 
3.0 1.862 0 -3.0 1e-06 
0.05 1.863 0 -3.0 1e-06 
3.0 1.863 0 -3.0 1e-06 
0.05 1.864 0 -3.0 1e-06 
3.0 1.864 0 -3.0 1e-06 
0.05 1.865 0 -3.0 1e-06 
3.0 1.865 0 -3.0 1e-06 
0.05 1.866 0 -3.0 1e-06 
3.0 1.866 0 -3.0 1e-06 
0.05 1.867 0 -3.0 1e-06 
3.0 1.867 0 -3.0 1e-06 
0.05 1.868 0 -3.0 1e-06 
3.0 1.868 0 -3.0 1e-06 
0.05 1.869 0 -3.0 1e-06 
3.0 1.869 0 -3.0 1e-06 
0.05 1.87 0 -3.0 1e-06 
3.0 1.87 0 -3.0 1e-06 
0.05 1.871 0 -3.0 1e-06 
3.0 1.871 0 -3.0 1e-06 
0.05 1.872 0 -3.0 1e-06 
3.0 1.872 0 -3.0 1e-06 
0.05 1.873 0 -3.0 1e-06 
3.0 1.873 0 -3.0 1e-06 
0.05 1.874 0 -3.0 1e-06 
3.0 1.874 0 -3.0 1e-06 
0.05 1.875 0 -3.0 1e-06 
3.0 1.875 0 -3.0 1e-06 
0.05 1.876 0 -3.0 1e-06 
3.0 1.876 0 -3.0 1e-06 
0.05 1.877 0 -3.0 1e-06 
3.0 1.877 0 -3.0 1e-06 
0.05 1.878 0 -3.0 1e-06 
3.0 1.878 0 -3.0 1e-06 
0.05 1.879 0 -3.0 1e-06 
3.0 1.879 0 -3.0 1e-06 
0.05 1.88 0 -3.0 1e-06 
3.0 1.88 0 -3.0 1e-06 
0.05 1.881 0 -3.0 1e-06 
3.0 1.881 0 -3.0 1e-06 
0.05 1.882 0 -3.0 1e-06 
3.0 1.882 0 -3.0 1e-06 
0.05 1.883 0 -3.0 1e-06 
3.0 1.883 0 -3.0 1e-06 
0.05 1.884 0 -3.0 1e-06 
3.0 1.884 0 -3.0 1e-06 
0.05 1.885 0 -3.0 1e-06 
3.0 1.885 0 -3.0 1e-06 
0.05 1.886 0 -3.0 1e-06 
3.0 1.886 0 -3.0 1e-06 
0.05 1.887 0 -3.0 1e-06 
3.0 1.887 0 -3.0 1e-06 
0.05 1.888 0 -3.0 1e-06 
3.0 1.888 0 -3.0 1e-06 
0.05 1.889 0 -3.0 1e-06 
3.0 1.889 0 -3.0 1e-06 
0.05 1.89 0 -3.0 1e-06 
3.0 1.89 0 -3.0 1e-06 
0.05 1.891 0 -3.0 1e-06 
3.0 1.891 0 -3.0 1e-06 
0.05 1.892 0 -3.0 1e-06 
3.0 1.892 0 -3.0 1e-06 
0.05 1.893 0 -3.0 1e-06 
3.0 1.893 0 -3.0 1e-06 
0.05 1.894 0 -3.0 1e-06 
3.0 1.894 0 -3.0 1e-06 
0.05 1.895 0 -3.0 1e-06 
3.0 1.895 0 -3.0 1e-06 
0.05 1.896 0 -3.0 1e-06 
3.0 1.896 0 -3.0 1e-06 
0.05 1.897 0 -3.0 1e-06 
3.0 1.897 0 -3.0 1e-06 
0.05 1.898 0 -3.0 1e-06 
3.0 1.898 0 -3.0 1e-06 
0.05 1.899 0 -3.0 1e-06 
3.0 1.899 0 -3.0 1e-06 
0.05 1.9 0 -3.0 1e-06 
3.0 1.9 0 -3.0 1e-06 
0.05 1.901 0 -3.0 1e-06 
3.0 1.901 0 -3.0 1e-06 
0.05 1.902 0 -3.0 1e-06 
3.0 1.902 0 -3.0 1e-06 
0.05 1.903 0 -3.0 1e-06 
3.0 1.903 0 -3.0 1e-06 
0.05 1.904 0 -3.0 1e-06 
3.0 1.904 0 -3.0 1e-06 
0.05 1.905 0 -3.0 1e-06 
3.0 1.905 0 -3.0 1e-06 
0.05 1.906 0 -3.0 1e-06 
3.0 1.906 0 -3.0 1e-06 
0.05 1.907 0 -3.0 1e-06 
3.0 1.907 0 -3.0 1e-06 
0.05 1.908 0 -3.0 1e-06 
3.0 1.908 0 -3.0 1e-06 
0.05 1.909 0 -3.0 1e-06 
3.0 1.909 0 -3.0 1e-06 
0.05 1.91 0 -3.0 1e-06 
3.0 1.91 0 -3.0 1e-06 
0.05 1.911 0 -3.0 1e-06 
3.0 1.911 0 -3.0 1e-06 
0.05 1.912 0 -3.0 1e-06 
3.0 1.912 0 -3.0 1e-06 
0.05 1.913 0 -3.0 1e-06 
3.0 1.913 0 -3.0 1e-06 
0.05 1.914 0 -3.0 1e-06 
3.0 1.914 0 -3.0 1e-06 
0.05 1.915 0 -3.0 1e-06 
3.0 1.915 0 -3.0 1e-06 
0.05 1.916 0 -3.0 1e-06 
3.0 1.916 0 -3.0 1e-06 
0.05 1.917 0 -3.0 1e-06 
3.0 1.917 0 -3.0 1e-06 
0.05 1.918 0 -3.0 1e-06 
3.0 1.918 0 -3.0 1e-06 
0.05 1.919 0 -3.0 1e-06 
3.0 1.919 0 -3.0 1e-06 
0.05 1.92 0 -3.0 1e-06 
3.0 1.92 0 -3.0 1e-06 
0.05 1.921 0 -3.0 1e-06 
3.0 1.921 0 -3.0 1e-06 
0.05 1.922 0 -3.0 1e-06 
3.0 1.922 0 -3.0 1e-06 
0.05 1.923 0 -3.0 1e-06 
3.0 1.923 0 -3.0 1e-06 
0.05 1.924 0 -3.0 1e-06 
3.0 1.924 0 -3.0 1e-06 
0.05 1.925 0 -3.0 1e-06 
3.0 1.925 0 -3.0 1e-06 
0.05 1.926 0 -3.0 1e-06 
3.0 1.926 0 -3.0 1e-06 
0.05 1.927 0 -3.0 1e-06 
3.0 1.927 0 -3.0 1e-06 
0.05 1.928 0 -3.0 1e-06 
3.0 1.928 0 -3.0 1e-06 
0.05 1.929 0 -3.0 1e-06 
3.0 1.929 0 -3.0 1e-06 
0.05 1.93 0 -3.0 1e-06 
3.0 1.93 0 -3.0 1e-06 
0.05 1.931 0 -3.0 1e-06 
3.0 1.931 0 -3.0 1e-06 
0.05 1.932 0 -3.0 1e-06 
3.0 1.932 0 -3.0 1e-06 
0.05 1.933 0 -3.0 1e-06 
3.0 1.933 0 -3.0 1e-06 
0.05 1.934 0 -3.0 1e-06 
3.0 1.934 0 -3.0 1e-06 
0.05 1.935 0 -3.0 1e-06 
3.0 1.935 0 -3.0 1e-06 
0.05 1.936 0 -3.0 1e-06 
3.0 1.936 0 -3.0 1e-06 
0.05 1.937 0 -3.0 1e-06 
3.0 1.937 0 -3.0 1e-06 
0.05 1.938 0 -3.0 1e-06 
3.0 1.938 0 -3.0 1e-06 
0.05 1.939 0 -3.0 1e-06 
3.0 1.939 0 -3.0 1e-06 
0.05 1.94 0 -3.0 1e-06 
3.0 1.94 0 -3.0 1e-06 
0.05 1.941 0 -3.0 1e-06 
3.0 1.941 0 -3.0 1e-06 
0.05 1.942 0 -3.0 1e-06 
3.0 1.942 0 -3.0 1e-06 
0.05 1.943 0 -3.0 1e-06 
3.0 1.943 0 -3.0 1e-06 
0.05 1.944 0 -3.0 1e-06 
3.0 1.944 0 -3.0 1e-06 
0.05 1.945 0 -3.0 1e-06 
3.0 1.945 0 -3.0 1e-06 
0.05 1.946 0 -3.0 1e-06 
3.0 1.946 0 -3.0 1e-06 
0.05 1.947 0 -3.0 1e-06 
3.0 1.947 0 -3.0 1e-06 
0.05 1.948 0 -3.0 1e-06 
3.0 1.948 0 -3.0 1e-06 
0.05 1.949 0 -3.0 1e-06 
3.0 1.949 0 -3.0 1e-06 
0.05 1.95 0 -3.0 1e-06 
3.0 1.95 0 -3.0 1e-06 
0.05 1.951 0 -3.0 1e-06 
3.0 1.951 0 -3.0 1e-06 
0.05 1.952 0 -3.0 1e-06 
3.0 1.952 0 -3.0 1e-06 
0.05 1.953 0 -3.0 1e-06 
3.0 1.953 0 -3.0 1e-06 
0.05 1.954 0 -3.0 1e-06 
3.0 1.954 0 -3.0 1e-06 
0.05 1.955 0 -3.0 1e-06 
3.0 1.955 0 -3.0 1e-06 
0.05 1.956 0 -3.0 1e-06 
3.0 1.956 0 -3.0 1e-06 
0.05 1.957 0 -3.0 1e-06 
3.0 1.957 0 -3.0 1e-06 
0.05 1.958 0 -3.0 1e-06 
3.0 1.958 0 -3.0 1e-06 
0.05 1.959 0 -3.0 1e-06 
3.0 1.959 0 -3.0 1e-06 
0.05 1.96 0 -3.0 1e-06 
3.0 1.96 0 -3.0 1e-06 
0.05 1.961 0 -3.0 1e-06 
3.0 1.961 0 -3.0 1e-06 
0.05 1.962 0 -3.0 1e-06 
3.0 1.962 0 -3.0 1e-06 
0.05 1.963 0 -3.0 1e-06 
3.0 1.963 0 -3.0 1e-06 
0.05 1.964 0 -3.0 1e-06 
3.0 1.964 0 -3.0 1e-06 
0.05 1.965 0 -3.0 1e-06 
3.0 1.965 0 -3.0 1e-06 
0.05 1.966 0 -3.0 1e-06 
3.0 1.966 0 -3.0 1e-06 
0.05 1.967 0 -3.0 1e-06 
3.0 1.967 0 -3.0 1e-06 
0.05 1.968 0 -3.0 1e-06 
3.0 1.968 0 -3.0 1e-06 
0.05 1.969 0 -3.0 1e-06 
3.0 1.969 0 -3.0 1e-06 
0.05 1.97 0 -3.0 1e-06 
3.0 1.97 0 -3.0 1e-06 
0.05 1.971 0 -3.0 1e-06 
3.0 1.971 0 -3.0 1e-06 
0.05 1.972 0 -3.0 1e-06 
3.0 1.972 0 -3.0 1e-06 
0.05 1.973 0 -3.0 1e-06 
3.0 1.973 0 -3.0 1e-06 
0.05 1.974 0 -3.0 1e-06 
3.0 1.974 0 -3.0 1e-06 
0.05 1.975 0 -3.0 1e-06 
3.0 1.975 0 -3.0 1e-06 
0.05 1.976 0 -3.0 1e-06 
3.0 1.976 0 -3.0 1e-06 
0.05 1.977 0 -3.0 1e-06 
3.0 1.977 0 -3.0 1e-06 
0.05 1.978 0 -3.0 1e-06 
3.0 1.978 0 -3.0 1e-06 
0.05 1.979 0 -3.0 1e-06 
3.0 1.979 0 -3.0 1e-06 
0.05 1.98 0 -3.0 1e-06 
3.0 1.98 0 -3.0 1e-06 
0.05 1.981 0 -3.0 1e-06 
3.0 1.981 0 -3.0 1e-06 
0.05 1.982 0 -3.0 1e-06 
3.0 1.982 0 -3.0 1e-06 
0.05 1.983 0 -3.0 1e-06 
3.0 1.983 0 -3.0 1e-06 
0.05 1.984 0 -3.0 1e-06 
3.0 1.984 0 -3.0 1e-06 
0.05 1.985 0 -3.0 1e-06 
3.0 1.985 0 -3.0 1e-06 
0.05 1.986 0 -3.0 1e-06 
3.0 1.986 0 -3.0 1e-06 
0.05 1.987 0 -3.0 1e-06 
3.0 1.987 0 -3.0 1e-06 
0.05 1.988 0 -3.0 1e-06 
3.0 1.988 0 -3.0 1e-06 
0.05 1.989 0 -3.0 1e-06 
3.0 1.989 0 -3.0 1e-06 
0.05 1.99 0 -3.0 1e-06 
3.0 1.99 0 -3.0 1e-06 
0.05 1.991 0 -3.0 1e-06 
3.0 1.991 0 -3.0 1e-06 
0.05 1.992 0 -3.0 1e-06 
3.0 1.992 0 -3.0 1e-06 
0.05 1.993 0 -3.0 1e-06 
3.0 1.993 0 -3.0 1e-06 
0.05 1.994 0 -3.0 1e-06 
3.0 1.994 0 -3.0 1e-06 
0.05 1.995 0 -3.0 1e-06 
3.0 1.995 0 -3.0 1e-06 
0.05 1.996 0 -3.0 1e-06 
3.0 1.996 0 -3.0 1e-06 
0.05 1.997 0 -3.0 1e-06 
3.0 1.997 0 -3.0 1e-06 
0.05 1.998 0 -3.0 1e-06 
3.0 1.998 0 -3.0 1e-06 
0.05 1.999 0 -3.0 1e-06 
3.0 1.999 0 -3.0 1e-06 
0.05 2.0 0 -3.0 1e-06 
3.0 2.0 0 -3.0 1e-06 
0.05 2.001 0 -3.0 1e-06 
3.0 2.001 0 -3.0 1e-06 
0.05 2.002 0 -3.0 1e-06 
3.0 2.002 0 -3.0 1e-06 
0.05 2.003 0 -3.0 1e-06 
3.0 2.003 0 -3.0 1e-06 
0.05 2.004 0 -3.0 1e-06 
3.0 2.004 0 -3.0 1e-06 
0.05 2.005 0 -3.0 1e-06 
3.0 2.005 0 -3.0 1e-06 
0.05 2.006 0 -3.0 1e-06 
3.0 2.006 0 -3.0 1e-06 
0.05 2.007 0 -3.0 1e-06 
3.0 2.007 0 -3.0 1e-06 
0.05 2.008 0 -3.0 1e-06 
3.0 2.008 0 -3.0 1e-06 
0.05 2.009 0 -3.0 1e-06 
3.0 2.009 0 -3.0 1e-06 
0.05 2.01 0 -3.0 1e-06 
3.0 2.01 0 -3.0 1e-06 
0.05 2.011 0 -3.0 1e-06 
3.0 2.011 0 -3.0 1e-06 
0.05 2.012 0 -3.0 1e-06 
3.0 2.012 0 -3.0 1e-06 
0.05 2.013 0 -3.0 1e-06 
3.0 2.013 0 -3.0 1e-06 
0.05 2.014 0 -3.0 1e-06 
3.0 2.014 0 -3.0 1e-06 
0.05 2.015 0 -3.0 1e-06 
3.0 2.015 0 -3.0 1e-06 
0.05 2.016 0 -3.0 1e-06 
3.0 2.016 0 -3.0 1e-06 
0.05 2.017 0 -3.0 1e-06 
3.0 2.017 0 -3.0 1e-06 
0.05 2.018 0 -3.0 1e-06 
3.0 2.018 0 -3.0 1e-06 
0.05 2.019 0 -3.0 1e-06 
3.0 2.019 0 -3.0 1e-06 
0.05 2.02 0 -3.0 1e-06 
3.0 2.02 0 -3.0 1e-06 
0.05 2.021 0 -3.0 1e-06 
3.0 2.021 0 -3.0 1e-06 
0.05 2.022 0 -3.0 1e-06 
3.0 2.022 0 -3.0 1e-06 
0.05 2.023 0 -3.0 1e-06 
3.0 2.023 0 -3.0 1e-06 
0.05 2.024 0 -3.0 1e-06 
3.0 2.024 0 -3.0 1e-06 
0.05 2.025 0 -3.0 1e-06 
3.0 2.025 0 -3.0 1e-06 
0.05 2.026 0 -3.0 1e-06 
3.0 2.026 0 -3.0 1e-06 
0.05 2.027 0 -3.0 1e-06 
3.0 2.027 0 -3.0 1e-06 
0.05 2.028 0 -3.0 1e-06 
3.0 2.028 0 -3.0 1e-06 
0.05 2.029 0 -3.0 1e-06 
3.0 2.029 0 -3.0 1e-06 
0.05 2.03 0 -3.0 1e-06 
3.0 2.03 0 -3.0 1e-06 
0.05 2.031 0 -3.0 1e-06 
3.0 2.031 0 -3.0 1e-06 
0.05 2.032 0 -3.0 1e-06 
3.0 2.032 0 -3.0 1e-06 
0.05 2.033 0 -3.0 1e-06 
3.0 2.033 0 -3.0 1e-06 
0.05 2.034 0 -3.0 1e-06 
3.0 2.034 0 -3.0 1e-06 
0.05 2.035 0 -3.0 1e-06 
3.0 2.035 0 -3.0 1e-06 
0.05 2.036 0 -3.0 1e-06 
3.0 2.036 0 -3.0 1e-06 
0.05 2.037 0 -3.0 1e-06 
3.0 2.037 0 -3.0 1e-06 
0.05 2.038 0 -3.0 1e-06 
3.0 2.038 0 -3.0 1e-06 
0.05 2.039 0 -3.0 1e-06 
3.0 2.039 0 -3.0 1e-06 
0.05 2.04 0 -3.0 1e-06 
3.0 2.04 0 -3.0 1e-06 
0.05 2.041 0 -3.0 1e-06 
3.0 2.041 0 -3.0 1e-06 
0.05 2.042 0 -3.0 1e-06 
3.0 2.042 0 -3.0 1e-06 
0.05 2.043 0 -3.0 1e-06 
3.0 2.043 0 -3.0 1e-06 
0.05 2.044 0 -3.0 1e-06 
3.0 2.044 0 -3.0 1e-06 
0.05 2.045 0 -3.0 1e-06 
3.0 2.045 0 -3.0 1e-06 
0.05 2.046 0 -3.0 1e-06 
3.0 2.046 0 -3.0 1e-06 
0.05 2.047 0 -3.0 1e-06 
3.0 2.047 0 -3.0 1e-06 
0.05 2.048 0 -3.0 1e-06 
3.0 2.048 0 -3.0 1e-06 
0.05 2.049 0 -3.0 1e-06 
3.0 2.049 0 -3.0 1e-06 
0.05 2.05 0 -3.0 1e-06 
3.0 2.05 0 -3.0 1e-06 
0.05 2.051 0 -3.0 1e-06 
3.0 2.051 0 -3.0 1e-06 
0.05 2.052 0 -3.0 1e-06 
3.0 2.052 0 -3.0 1e-06 
0.05 2.053 0 -3.0 1e-06 
3.0 2.053 0 -3.0 1e-06 
0.05 2.054 0 -3.0 1e-06 
3.0 2.054 0 -3.0 1e-06 
0.05 2.055 0 -3.0 1e-06 
3.0 2.055 0 -3.0 1e-06 
0.05 2.056 0 -3.0 1e-06 
3.0 2.056 0 -3.0 1e-06 
0.05 2.057 0 -3.0 1e-06 
3.0 2.057 0 -3.0 1e-06 
0.05 2.058 0 -3.0 1e-06 
3.0 2.058 0 -3.0 1e-06 
0.05 2.059 0 -3.0 1e-06 
3.0 2.059 0 -3.0 1e-06 
0.05 2.06 0 -3.0 1e-06 
3.0 2.06 0 -3.0 1e-06 
0.05 2.061 0 -3.0 1e-06 
3.0 2.061 0 -3.0 1e-06 
0.05 2.062 0 -3.0 1e-06 
3.0 2.062 0 -3.0 1e-06 
0.05 2.063 0 -3.0 1e-06 
3.0 2.063 0 -3.0 1e-06 
0.05 2.064 0 -3.0 1e-06 
3.0 2.064 0 -3.0 1e-06 
0.05 2.065 0 -3.0 1e-06 
3.0 2.065 0 -3.0 1e-06 
0.05 2.066 0 -3.0 1e-06 
3.0 2.066 0 -3.0 1e-06 
0.05 2.067 0 -3.0 1e-06 
3.0 2.067 0 -3.0 1e-06 
0.05 2.068 0 -3.0 1e-06 
3.0 2.068 0 -3.0 1e-06 
0.05 2.069 0 -3.0 1e-06 
3.0 2.069 0 -3.0 1e-06 
0.05 2.07 0 -3.0 1e-06 
3.0 2.07 0 -3.0 1e-06 
0.05 2.071 0 -3.0 1e-06 
3.0 2.071 0 -3.0 1e-06 
0.05 2.072 0 -3.0 1e-06 
3.0 2.072 0 -3.0 1e-06 
0.05 2.073 0 -3.0 1e-06 
3.0 2.073 0 -3.0 1e-06 
0.05 2.074 0 -3.0 1e-06 
3.0 2.074 0 -3.0 1e-06 
0.05 2.075 0 -3.0 1e-06 
3.0 2.075 0 -3.0 1e-06 
0.05 2.076 0 -3.0 1e-06 
3.0 2.076 0 -3.0 1e-06 
0.05 2.077 0 -3.0 1e-06 
3.0 2.077 0 -3.0 1e-06 
0.05 2.078 0 -3.0 1e-06 
3.0 2.078 0 -3.0 1e-06 
0.05 2.079 0 -3.0 1e-06 
3.0 2.079 0 -3.0 1e-06 
0.05 2.08 0 -3.0 1e-06 
3.0 2.08 0 -3.0 1e-06 
0.05 2.081 0 -3.0 1e-06 
3.0 2.081 0 -3.0 1e-06 
0.05 2.082 0 -3.0 1e-06 
3.0 2.082 0 -3.0 1e-06 
0.05 2.083 0 -3.0 1e-06 
3.0 2.083 0 -3.0 1e-06 
0.05 2.084 0 -3.0 1e-06 
3.0 2.084 0 -3.0 1e-06 
0.05 2.085 0 -3.0 1e-06 
3.0 2.085 0 -3.0 1e-06 
0.05 2.086 0 -3.0 1e-06 
3.0 2.086 0 -3.0 1e-06 
0.05 2.087 0 -3.0 1e-06 
3.0 2.087 0 -3.0 1e-06 
0.05 2.088 0 -3.0 1e-06 
3.0 2.088 0 -3.0 1e-06 
0.05 2.089 0 -3.0 1e-06 
3.0 2.089 0 -3.0 1e-06 
0.05 2.09 0 -3.0 1e-06 
3.0 2.09 0 -3.0 1e-06 
0.05 2.091 0 -3.0 1e-06 
3.0 2.091 0 -3.0 1e-06 
0.05 2.092 0 -3.0 1e-06 
3.0 2.092 0 -3.0 1e-06 
0.05 2.093 0 -3.0 1e-06 
3.0 2.093 0 -3.0 1e-06 
0.05 2.094 0 -3.0 1e-06 
3.0 2.094 0 -3.0 1e-06 
0.05 2.095 0 -3.0 1e-06 
3.0 2.095 0 -3.0 1e-06 
0.05 2.096 0 -3.0 1e-06 
3.0 2.096 0 -3.0 1e-06 
0.05 2.097 0 -3.0 1e-06 
3.0 2.097 0 -3.0 1e-06 
0.05 2.098 0 -3.0 1e-06 
3.0 2.098 0 -3.0 1e-06 
0.05 2.099 0 -3.0 1e-06 
3.0 2.099 0 -3.0 1e-06 
0.05 2.1 0 -3.0 1e-06 
3.0 2.1 0 -3.0 1e-06 
0.05 2.101 0 -3.0 1e-06 
3.0 2.101 0 -3.0 1e-06 
0.05 2.102 0 -3.0 1e-06 
3.0 2.102 0 -3.0 1e-06 
0.05 2.103 0 -3.0 1e-06 
3.0 2.103 0 -3.0 1e-06 
0.05 2.104 0 -3.0 1e-06 
3.0 2.104 0 -3.0 1e-06 
0.05 2.105 0 -3.0 1e-06 
3.0 2.105 0 -3.0 1e-06 
0.05 2.106 0 -3.0 1e-06 
3.0 2.106 0 -3.0 1e-06 
0.05 2.107 0 -3.0 1e-06 
3.0 2.107 0 -3.0 1e-06 
0.05 2.108 0 -3.0 1e-06 
3.0 2.108 0 -3.0 1e-06 
0.05 2.109 0 -3.0 1e-06 
3.0 2.109 0 -3.0 1e-06 
0.05 2.11 0 -3.0 1e-06 
3.0 2.11 0 -3.0 1e-06 
0.05 2.111 0 -3.0 1e-06 
3.0 2.111 0 -3.0 1e-06 
0.05 2.112 0 -3.0 1e-06 
3.0 2.112 0 -3.0 1e-06 
0.05 2.113 0 -3.0 1e-06 
3.0 2.113 0 -3.0 1e-06 
0.05 2.114 0 -3.0 1e-06 
3.0 2.114 0 -3.0 1e-06 
0.05 2.115 0 -3.0 1e-06 
3.0 2.115 0 -3.0 1e-06 
0.05 2.116 0 -3.0 1e-06 
3.0 2.116 0 -3.0 1e-06 
0.05 2.117 0 -3.0 1e-06 
3.0 2.117 0 -3.0 1e-06 
0.05 2.118 0 -3.0 1e-06 
3.0 2.118 0 -3.0 1e-06 
0.05 2.119 0 -3.0 1e-06 
3.0 2.119 0 -3.0 1e-06 
0.05 2.12 0 -3.0 1e-06 
3.0 2.12 0 -3.0 1e-06 
0.05 2.121 0 -3.0 1e-06 
3.0 2.121 0 -3.0 1e-06 
0.05 2.122 0 -3.0 1e-06 
3.0 2.122 0 -3.0 1e-06 
0.05 2.123 0 -3.0 1e-06 
3.0 2.123 0 -3.0 1e-06 
0.05 2.124 0 -3.0 1e-06 
3.0 2.124 0 -3.0 1e-06 
0.05 2.125 0 -3.0 1e-06 
3.0 2.125 0 -3.0 1e-06 
0.05 2.126 0 -3.0 1e-06 
3.0 2.126 0 -3.0 1e-06 
0.05 2.127 0 -3.0 1e-06 
3.0 2.127 0 -3.0 1e-06 
0.05 2.128 0 -3.0 1e-06 
3.0 2.128 0 -3.0 1e-06 
0.05 2.129 0 -3.0 1e-06 
3.0 2.129 0 -3.0 1e-06 
0.05 2.13 0 -3.0 1e-06 
3.0 2.13 0 -3.0 1e-06 
0.05 2.131 0 -3.0 1e-06 
3.0 2.131 0 -3.0 1e-06 
0.05 2.132 0 -3.0 1e-06 
3.0 2.132 0 -3.0 1e-06 
0.05 2.133 0 -3.0 1e-06 
3.0 2.133 0 -3.0 1e-06 
0.05 2.134 0 -3.0 1e-06 
3.0 2.134 0 -3.0 1e-06 
0.05 2.135 0 -3.0 1e-06 
3.0 2.135 0 -3.0 1e-06 
0.05 2.136 0 -3.0 1e-06 
3.0 2.136 0 -3.0 1e-06 
0.05 2.137 0 -3.0 1e-06 
3.0 2.137 0 -3.0 1e-06 
0.05 2.138 0 -3.0 1e-06 
3.0 2.138 0 -3.0 1e-06 
0.05 2.139 0 -3.0 1e-06 
3.0 2.139 0 -3.0 1e-06 
0.05 2.14 0 -3.0 1e-06 
3.0 2.14 0 -3.0 1e-06 
0.05 2.141 0 -3.0 1e-06 
3.0 2.141 0 -3.0 1e-06 
0.05 2.142 0 -3.0 1e-06 
3.0 2.142 0 -3.0 1e-06 
0.05 2.143 0 -3.0 1e-06 
3.0 2.143 0 -3.0 1e-06 
0.05 2.144 0 -3.0 1e-06 
3.0 2.144 0 -3.0 1e-06 
0.05 2.145 0 -3.0 1e-06 
3.0 2.145 0 -3.0 1e-06 
0.05 2.146 0 -3.0 1e-06 
3.0 2.146 0 -3.0 1e-06 
0.05 2.147 0 -3.0 1e-06 
3.0 2.147 0 -3.0 1e-06 
0.05 2.148 0 -3.0 1e-06 
3.0 2.148 0 -3.0 1e-06 
0.05 2.149 0 -3.0 1e-06 
3.0 2.149 0 -3.0 1e-06 
0.05 2.15 0 -3.0 1e-06 
3.0 2.15 0 -3.0 1e-06 
0.05 2.151 0 -3.0 1e-06 
3.0 2.151 0 -3.0 1e-06 
0.05 2.152 0 -3.0 1e-06 
3.0 2.152 0 -3.0 1e-06 
0.05 2.153 0 -3.0 1e-06 
3.0 2.153 0 -3.0 1e-06 
0.05 2.154 0 -3.0 1e-06 
3.0 2.154 0 -3.0 1e-06 
0.05 2.155 0 -3.0 1e-06 
3.0 2.155 0 -3.0 1e-06 
0.05 2.156 0 -3.0 1e-06 
3.0 2.156 0 -3.0 1e-06 
0.05 2.157 0 -3.0 1e-06 
3.0 2.157 0 -3.0 1e-06 
0.05 2.158 0 -3.0 1e-06 
3.0 2.158 0 -3.0 1e-06 
0.05 2.159 0 -3.0 1e-06 
3.0 2.159 0 -3.0 1e-06 
0.05 2.16 0 -3.0 1e-06 
3.0 2.16 0 -3.0 1e-06 
0.05 2.161 0 -3.0 1e-06 
3.0 2.161 0 -3.0 1e-06 
0.05 2.162 0 -3.0 1e-06 
3.0 2.162 0 -3.0 1e-06 
0.05 2.163 0 -3.0 1e-06 
3.0 2.163 0 -3.0 1e-06 
0.05 2.164 0 -3.0 1e-06 
3.0 2.164 0 -3.0 1e-06 
0.05 2.165 0 -3.0 1e-06 
3.0 2.165 0 -3.0 1e-06 
0.05 2.166 0 -3.0 1e-06 
3.0 2.166 0 -3.0 1e-06 
0.05 2.167 0 -3.0 1e-06 
3.0 2.167 0 -3.0 1e-06 
0.05 2.168 0 -3.0 1e-06 
3.0 2.168 0 -3.0 1e-06 
0.05 2.169 0 -3.0 1e-06 
3.0 2.169 0 -3.0 1e-06 
0.05 2.17 0 -3.0 1e-06 
3.0 2.17 0 -3.0 1e-06 
0.05 2.171 0 -3.0 1e-06 
3.0 2.171 0 -3.0 1e-06 
0.05 2.172 0 -3.0 1e-06 
3.0 2.172 0 -3.0 1e-06 
0.05 2.173 0 -3.0 1e-06 
3.0 2.173 0 -3.0 1e-06 
0.05 2.174 0 -3.0 1e-06 
3.0 2.174 0 -3.0 1e-06 
0.05 2.175 0 -3.0 1e-06 
3.0 2.175 0 -3.0 1e-06 
0.05 2.176 0 -3.0 1e-06 
3.0 2.176 0 -3.0 1e-06 
0.05 2.177 0 -3.0 1e-06 
3.0 2.177 0 -3.0 1e-06 
0.05 2.178 0 -3.0 1e-06 
3.0 2.178 0 -3.0 1e-06 
0.05 2.179 0 -3.0 1e-06 
3.0 2.179 0 -3.0 1e-06 
0.05 2.18 0 -3.0 1e-06 
3.0 2.18 0 -3.0 1e-06 
0.05 2.181 0 -3.0 1e-06 
3.0 2.181 0 -3.0 1e-06 
0.05 2.182 0 -3.0 1e-06 
3.0 2.182 0 -3.0 1e-06 
0.05 2.183 0 -3.0 1e-06 
3.0 2.183 0 -3.0 1e-06 
0.05 2.184 0 -3.0 1e-06 
3.0 2.184 0 -3.0 1e-06 
0.05 2.185 0 -3.0 1e-06 
3.0 2.185 0 -3.0 1e-06 
0.05 2.186 0 -3.0 1e-06 
3.0 2.186 0 -3.0 1e-06 
0.05 2.187 0 -3.0 1e-06 
3.0 2.187 0 -3.0 1e-06 
0.05 2.188 0 -3.0 1e-06 
3.0 2.188 0 -3.0 1e-06 
0.05 2.189 0 -3.0 1e-06 
3.0 2.189 0 -3.0 1e-06 
0.05 2.19 0 -3.0 1e-06 
3.0 2.19 0 -3.0 1e-06 
0.05 2.191 0 -3.0 1e-06 
3.0 2.191 0 -3.0 1e-06 
0.05 2.192 0 -3.0 1e-06 
3.0 2.192 0 -3.0 1e-06 
0.05 2.193 0 -3.0 1e-06 
3.0 2.193 0 -3.0 1e-06 
0.05 2.194 0 -3.0 1e-06 
3.0 2.194 0 -3.0 1e-06 
0.05 2.195 0 -3.0 1e-06 
3.0 2.195 0 -3.0 1e-06 
0.05 2.196 0 -3.0 1e-06 
3.0 2.196 0 -3.0 1e-06 
0.05 2.197 0 -3.0 1e-06 
3.0 2.197 0 -3.0 1e-06 
0.05 2.198 0 -3.0 1e-06 
3.0 2.198 0 -3.0 1e-06 
0.05 2.199 0 -3.0 1e-06 
3.0 2.199 0 -3.0 1e-06 
0.05 2.2 0 -3.0 1e-06 
3.0 2.2 0 -3.0 1e-06 
0.05 2.201 0 -3.0 1e-06 
3.0 2.201 0 -3.0 1e-06 
0.05 2.202 0 -3.0 1e-06 
3.0 2.202 0 -3.0 1e-06 
0.05 2.203 0 -3.0 1e-06 
3.0 2.203 0 -3.0 1e-06 
0.05 2.204 0 -3.0 1e-06 
3.0 2.204 0 -3.0 1e-06 
0.05 2.205 0 -3.0 1e-06 
3.0 2.205 0 -3.0 1e-06 
0.05 2.206 0 -3.0 1e-06 
3.0 2.206 0 -3.0 1e-06 
0.05 2.207 0 -3.0 1e-06 
3.0 2.207 0 -3.0 1e-06 
0.05 2.208 0 -3.0 1e-06 
3.0 2.208 0 -3.0 1e-06 
0.05 2.209 0 -3.0 1e-06 
3.0 2.209 0 -3.0 1e-06 
0.05 2.21 0 -3.0 1e-06 
3.0 2.21 0 -3.0 1e-06 
0.05 2.211 0 -3.0 1e-06 
3.0 2.211 0 -3.0 1e-06 
0.05 2.212 0 -3.0 1e-06 
3.0 2.212 0 -3.0 1e-06 
0.05 2.213 0 -3.0 1e-06 
3.0 2.213 0 -3.0 1e-06 
0.05 2.214 0 -3.0 1e-06 
3.0 2.214 0 -3.0 1e-06 
0.05 2.215 0 -3.0 1e-06 
3.0 2.215 0 -3.0 1e-06 
0.05 2.216 0 -3.0 1e-06 
3.0 2.216 0 -3.0 1e-06 
0.05 2.217 0 -3.0 1e-06 
3.0 2.217 0 -3.0 1e-06 
0.05 2.218 0 -3.0 1e-06 
3.0 2.218 0 -3.0 1e-06 
0.05 2.219 0 -3.0 1e-06 
3.0 2.219 0 -3.0 1e-06 
0.05 2.22 0 -3.0 1e-06 
3.0 2.22 0 -3.0 1e-06 
0.05 2.221 0 -3.0 1e-06 
3.0 2.221 0 -3.0 1e-06 
0.05 2.222 0 -3.0 1e-06 
3.0 2.222 0 -3.0 1e-06 
0.05 2.223 0 -3.0 1e-06 
3.0 2.223 0 -3.0 1e-06 
0.05 2.224 0 -3.0 1e-06 
3.0 2.224 0 -3.0 1e-06 
0.05 2.225 0 -3.0 1e-06 
3.0 2.225 0 -3.0 1e-06 
0.05 2.226 0 -3.0 1e-06 
3.0 2.226 0 -3.0 1e-06 
0.05 2.227 0 -3.0 1e-06 
3.0 2.227 0 -3.0 1e-06 
0.05 2.228 0 -3.0 1e-06 
3.0 2.228 0 -3.0 1e-06 
0.05 2.229 0 -3.0 1e-06 
3.0 2.229 0 -3.0 1e-06 
0.05 2.23 0 -3.0 1e-06 
3.0 2.23 0 -3.0 1e-06 
0.05 2.231 0 -3.0 1e-06 
3.0 2.231 0 -3.0 1e-06 
0.05 2.232 0 -3.0 1e-06 
3.0 2.232 0 -3.0 1e-06 
0.05 2.233 0 -3.0 1e-06 
3.0 2.233 0 -3.0 1e-06 
0.05 2.234 0 -3.0 1e-06 
3.0 2.234 0 -3.0 1e-06 
0.05 2.235 0 -3.0 1e-06 
3.0 2.235 0 -3.0 1e-06 
0.05 2.236 0 -3.0 1e-06 
3.0 2.236 0 -3.0 1e-06 
0.05 2.237 0 -3.0 1e-06 
3.0 2.237 0 -3.0 1e-06 
0.05 2.238 0 -3.0 1e-06 
3.0 2.238 0 -3.0 1e-06 
0.05 2.239 0 -3.0 1e-06 
3.0 2.239 0 -3.0 1e-06 
0.05 2.24 0 -3.0 1e-06 
3.0 2.24 0 -3.0 1e-06 
0.05 2.241 0 -3.0 1e-06 
3.0 2.241 0 -3.0 1e-06 
0.05 2.242 0 -3.0 1e-06 
3.0 2.242 0 -3.0 1e-06 
0.05 2.243 0 -3.0 1e-06 
3.0 2.243 0 -3.0 1e-06 
0.05 2.244 0 -3.0 1e-06 
3.0 2.244 0 -3.0 1e-06 
0.05 2.245 0 -3.0 1e-06 
3.0 2.245 0 -3.0 1e-06 
0.05 2.246 0 -3.0 1e-06 
3.0 2.246 0 -3.0 1e-06 
0.05 2.247 0 -3.0 1e-06 
3.0 2.247 0 -3.0 1e-06 
0.05 2.248 0 -3.0 1e-06 
3.0 2.248 0 -3.0 1e-06 
0.05 2.249 0 -3.0 1e-06 
3.0 2.249 0 -3.0 1e-06 
0.05 2.25 0 -3.0 1e-06 
3.0 2.25 0 -3.0 1e-06 
0.05 2.251 0 -3.0 1e-06 
3.0 2.251 0 -3.0 1e-06 
0.05 2.252 0 -3.0 1e-06 
3.0 2.252 0 -3.0 1e-06 
0.05 2.253 0 -3.0 1e-06 
3.0 2.253 0 -3.0 1e-06 
0.05 2.254 0 -3.0 1e-06 
3.0 2.254 0 -3.0 1e-06 
0.05 2.255 0 -3.0 1e-06 
3.0 2.255 0 -3.0 1e-06 
0.05 2.256 0 -3.0 1e-06 
3.0 2.256 0 -3.0 1e-06 
0.05 2.257 0 -3.0 1e-06 
3.0 2.257 0 -3.0 1e-06 
0.05 2.258 0 -3.0 1e-06 
3.0 2.258 0 -3.0 1e-06 
0.05 2.259 0 -3.0 1e-06 
3.0 2.259 0 -3.0 1e-06 
0.05 2.26 0 -3.0 1e-06 
3.0 2.26 0 -3.0 1e-06 
0.05 2.261 0 -3.0 1e-06 
3.0 2.261 0 -3.0 1e-06 
0.05 2.262 0 -3.0 1e-06 
3.0 2.262 0 -3.0 1e-06 
0.05 2.263 0 -3.0 1e-06 
3.0 2.263 0 -3.0 1e-06 
0.05 2.264 0 -3.0 1e-06 
3.0 2.264 0 -3.0 1e-06 
0.05 2.265 0 -3.0 1e-06 
3.0 2.265 0 -3.0 1e-06 
0.05 2.266 0 -3.0 1e-06 
3.0 2.266 0 -3.0 1e-06 
0.05 2.267 0 -3.0 1e-06 
3.0 2.267 0 -3.0 1e-06 
0.05 2.268 0 -3.0 1e-06 
3.0 2.268 0 -3.0 1e-06 
0.05 2.269 0 -3.0 1e-06 
3.0 2.269 0 -3.0 1e-06 
0.05 2.27 0 -3.0 1e-06 
3.0 2.27 0 -3.0 1e-06 
0.05 2.271 0 -3.0 1e-06 
3.0 2.271 0 -3.0 1e-06 
0.05 2.272 0 -3.0 1e-06 
3.0 2.272 0 -3.0 1e-06 
0.05 2.273 0 -3.0 1e-06 
3.0 2.273 0 -3.0 1e-06 
0.05 2.274 0 -3.0 1e-06 
3.0 2.274 0 -3.0 1e-06 
0.05 2.275 0 -3.0 1e-06 
3.0 2.275 0 -3.0 1e-06 
0.05 2.276 0 -3.0 1e-06 
3.0 2.276 0 -3.0 1e-06 
0.05 2.277 0 -3.0 1e-06 
3.0 2.277 0 -3.0 1e-06 
0.05 2.278 0 -3.0 1e-06 
3.0 2.278 0 -3.0 1e-06 
0.05 2.279 0 -3.0 1e-06 
3.0 2.279 0 -3.0 1e-06 
0.05 2.28 0 -3.0 1e-06 
3.0 2.28 0 -3.0 1e-06 
0.05 2.281 0 -3.0 1e-06 
3.0 2.281 0 -3.0 1e-06 
0.05 2.282 0 -3.0 1e-06 
3.0 2.282 0 -3.0 1e-06 
0.05 2.283 0 -3.0 1e-06 
3.0 2.283 0 -3.0 1e-06 
0.05 2.284 0 -3.0 1e-06 
3.0 2.284 0 -3.0 1e-06 
0.05 2.285 0 -3.0 1e-06 
3.0 2.285 0 -3.0 1e-06 
0.05 2.286 0 -3.0 1e-06 
3.0 2.286 0 -3.0 1e-06 
0.05 2.287 0 -3.0 1e-06 
3.0 2.287 0 -3.0 1e-06 
0.05 2.288 0 -3.0 1e-06 
3.0 2.288 0 -3.0 1e-06 
0.05 2.289 0 -3.0 1e-06 
3.0 2.289 0 -3.0 1e-06 
0.05 2.29 0 -3.0 1e-06 
3.0 2.29 0 -3.0 1e-06 
0.05 2.291 0 -3.0 1e-06 
3.0 2.291 0 -3.0 1e-06 
0.05 2.292 0 -3.0 1e-06 
3.0 2.292 0 -3.0 1e-06 
0.05 2.293 0 -3.0 1e-06 
3.0 2.293 0 -3.0 1e-06 
0.05 2.294 0 -3.0 1e-06 
3.0 2.294 0 -3.0 1e-06 
0.05 2.295 0 -3.0 1e-06 
3.0 2.295 0 -3.0 1e-06 
0.05 2.296 0 -3.0 1e-06 
3.0 2.296 0 -3.0 1e-06 
0.05 2.297 0 -3.0 1e-06 
3.0 2.297 0 -3.0 1e-06 
0.05 2.298 0 -3.0 1e-06 
3.0 2.298 0 -3.0 1e-06 
0.05 2.299 0 -3.0 1e-06 
3.0 2.299 0 -3.0 1e-06 
0.05 2.3 0 -3.0 1e-06 
3.0 2.3 0 -3.0 1e-06 
0.05 2.301 0 -3.0 1e-06 
3.0 2.301 0 -3.0 1e-06 
0.05 2.302 0 -3.0 1e-06 
3.0 2.302 0 -3.0 1e-06 
0.05 2.303 0 -3.0 1e-06 
3.0 2.303 0 -3.0 1e-06 
0.05 2.304 0 -3.0 1e-06 
3.0 2.304 0 -3.0 1e-06 
0.05 2.305 0 -3.0 1e-06 
3.0 2.305 0 -3.0 1e-06 
0.05 2.306 0 -3.0 1e-06 
3.0 2.306 0 -3.0 1e-06 
0.05 2.307 0 -3.0 1e-06 
3.0 2.307 0 -3.0 1e-06 
0.05 2.308 0 -3.0 1e-06 
3.0 2.308 0 -3.0 1e-06 
0.05 2.309 0 -3.0 1e-06 
3.0 2.309 0 -3.0 1e-06 
0.05 2.31 0 -3.0 1e-06 
3.0 2.31 0 -3.0 1e-06 
0.05 2.311 0 -3.0 1e-06 
3.0 2.311 0 -3.0 1e-06 
0.05 2.312 0 -3.0 1e-06 
3.0 2.312 0 -3.0 1e-06 
0.05 2.313 0 -3.0 1e-06 
3.0 2.313 0 -3.0 1e-06 
0.05 2.314 0 -3.0 1e-06 
3.0 2.314 0 -3.0 1e-06 
0.05 2.315 0 -3.0 1e-06 
3.0 2.315 0 -3.0 1e-06 
0.05 2.316 0 -3.0 1e-06 
3.0 2.316 0 -3.0 1e-06 
0.05 2.317 0 -3.0 1e-06 
3.0 2.317 0 -3.0 1e-06 
0.05 2.318 0 -3.0 1e-06 
3.0 2.318 0 -3.0 1e-06 
0.05 2.319 0 -3.0 1e-06 
3.0 2.319 0 -3.0 1e-06 
0.05 2.32 0 -3.0 1e-06 
3.0 2.32 0 -3.0 1e-06 
0.05 2.321 0 -3.0 1e-06 
3.0 2.321 0 -3.0 1e-06 
0.05 2.322 0 -3.0 1e-06 
3.0 2.322 0 -3.0 1e-06 
0.05 2.323 0 -3.0 1e-06 
3.0 2.323 0 -3.0 1e-06 
0.05 2.324 0 -3.0 1e-06 
3.0 2.324 0 -3.0 1e-06 
0.05 2.325 0 -3.0 1e-06 
3.0 2.325 0 -3.0 1e-06 
0.05 2.326 0 -3.0 1e-06 
3.0 2.326 0 -3.0 1e-06 
0.05 2.327 0 -3.0 1e-06 
3.0 2.327 0 -3.0 1e-06 
0.05 2.328 0 -3.0 1e-06 
3.0 2.328 0 -3.0 1e-06 
0.05 2.329 0 -3.0 1e-06 
3.0 2.329 0 -3.0 1e-06 
0.05 2.33 0 -3.0 1e-06 
3.0 2.33 0 -3.0 1e-06 
0.05 2.331 0 -3.0 1e-06 
3.0 2.331 0 -3.0 1e-06 
0.05 2.332 0 -3.0 1e-06 
3.0 2.332 0 -3.0 1e-06 
0.05 2.333 0 -3.0 1e-06 
3.0 2.333 0 -3.0 1e-06 
0.05 2.334 0 -3.0 1e-06 
3.0 2.334 0 -3.0 1e-06 
0.05 2.335 0 -3.0 1e-06 
3.0 2.335 0 -3.0 1e-06 
0.05 2.336 0 -3.0 1e-06 
3.0 2.336 0 -3.0 1e-06 
0.05 2.337 0 -3.0 1e-06 
3.0 2.337 0 -3.0 1e-06 
0.05 2.338 0 -3.0 1e-06 
3.0 2.338 0 -3.0 1e-06 
0.05 2.339 0 -3.0 1e-06 
3.0 2.339 0 -3.0 1e-06 
0.05 2.34 0 -3.0 1e-06 
3.0 2.34 0 -3.0 1e-06 
0.05 2.341 0 -3.0 1e-06 
3.0 2.341 0 -3.0 1e-06 
0.05 2.342 0 -3.0 1e-06 
3.0 2.342 0 -3.0 1e-06 
0.05 2.343 0 -3.0 1e-06 
3.0 2.343 0 -3.0 1e-06 
0.05 2.344 0 -3.0 1e-06 
3.0 2.344 0 -3.0 1e-06 
0.05 2.345 0 -3.0 1e-06 
3.0 2.345 0 -3.0 1e-06 
0.05 2.346 0 -3.0 1e-06 
3.0 2.346 0 -3.0 1e-06 
0.05 2.347 0 -3.0 1e-06 
3.0 2.347 0 -3.0 1e-06 
0.05 2.348 0 -3.0 1e-06 
3.0 2.348 0 -3.0 1e-06 
0.05 2.349 0 -3.0 1e-06 
3.0 2.349 0 -3.0 1e-06 
0.05 2.35 0 -3.0 1e-06 
3.0 2.35 0 -3.0 1e-06 
0.05 2.351 0 -3.0 1e-06 
3.0 2.351 0 -3.0 1e-06 
0.05 2.352 0 -3.0 1e-06 
3.0 2.352 0 -3.0 1e-06 
0.05 2.353 0 -3.0 1e-06 
3.0 2.353 0 -3.0 1e-06 
0.05 2.354 0 -3.0 1e-06 
3.0 2.354 0 -3.0 1e-06 
0.05 2.355 0 -3.0 1e-06 
3.0 2.355 0 -3.0 1e-06 
0.05 2.356 0 -3.0 1e-06 
3.0 2.356 0 -3.0 1e-06 
0.05 2.357 0 -3.0 1e-06 
3.0 2.357 0 -3.0 1e-06 
0.05 2.358 0 -3.0 1e-06 
3.0 2.358 0 -3.0 1e-06 
0.05 2.359 0 -3.0 1e-06 
3.0 2.359 0 -3.0 1e-06 
0.05 2.36 0 -3.0 1e-06 
3.0 2.36 0 -3.0 1e-06 
0.05 2.361 0 -3.0 1e-06 
3.0 2.361 0 -3.0 1e-06 
0.05 2.362 0 -3.0 1e-06 
3.0 2.362 0 -3.0 1e-06 
0.05 2.363 0 -3.0 1e-06 
3.0 2.363 0 -3.0 1e-06 
0.05 2.364 0 -3.0 1e-06 
3.0 2.364 0 -3.0 1e-06 
0.05 2.365 0 -3.0 1e-06 
3.0 2.365 0 -3.0 1e-06 
0.05 2.366 0 -3.0 1e-06 
3.0 2.366 0 -3.0 1e-06 
0.05 2.367 0 -3.0 1e-06 
3.0 2.367 0 -3.0 1e-06 
0.05 2.368 0 -3.0 1e-06 
3.0 2.368 0 -3.0 1e-06 
0.05 2.369 0 -3.0 1e-06 
3.0 2.369 0 -3.0 1e-06 
0.05 2.37 0 -3.0 1e-06 
3.0 2.37 0 -3.0 1e-06 
0.05 2.371 0 -3.0 1e-06 
3.0 2.371 0 -3.0 1e-06 
0.05 2.372 0 -3.0 1e-06 
3.0 2.372 0 -3.0 1e-06 
0.05 2.373 0 -3.0 1e-06 
3.0 2.373 0 -3.0 1e-06 
0.05 2.374 0 -3.0 1e-06 
3.0 2.374 0 -3.0 1e-06 
0.05 2.375 0 -3.0 1e-06 
3.0 2.375 0 -3.0 1e-06 
0.05 2.376 0 -3.0 1e-06 
3.0 2.376 0 -3.0 1e-06 
0.05 2.377 0 -3.0 1e-06 
3.0 2.377 0 -3.0 1e-06 
0.05 2.378 0 -3.0 1e-06 
3.0 2.378 0 -3.0 1e-06 
0.05 2.379 0 -3.0 1e-06 
3.0 2.379 0 -3.0 1e-06 
0.05 2.38 0 -3.0 1e-06 
3.0 2.38 0 -3.0 1e-06 
0.05 2.381 0 -3.0 1e-06 
3.0 2.381 0 -3.0 1e-06 
0.05 2.382 0 -3.0 1e-06 
3.0 2.382 0 -3.0 1e-06 
0.05 2.383 0 -3.0 1e-06 
3.0 2.383 0 -3.0 1e-06 
0.05 2.384 0 -3.0 1e-06 
3.0 2.384 0 -3.0 1e-06 
0.05 2.385 0 -3.0 1e-06 
3.0 2.385 0 -3.0 1e-06 
0.05 2.386 0 -3.0 1e-06 
3.0 2.386 0 -3.0 1e-06 
0.05 2.387 0 -3.0 1e-06 
3.0 2.387 0 -3.0 1e-06 
0.05 2.388 0 -3.0 1e-06 
3.0 2.388 0 -3.0 1e-06 
0.05 2.389 0 -3.0 1e-06 
3.0 2.389 0 -3.0 1e-06 
0.05 2.39 0 -3.0 1e-06 
3.0 2.39 0 -3.0 1e-06 
0.05 2.391 0 -3.0 1e-06 
3.0 2.391 0 -3.0 1e-06 
0.05 2.392 0 -3.0 1e-06 
3.0 2.392 0 -3.0 1e-06 
0.05 2.393 0 -3.0 1e-06 
3.0 2.393 0 -3.0 1e-06 
0.05 2.394 0 -3.0 1e-06 
3.0 2.394 0 -3.0 1e-06 
0.05 2.395 0 -3.0 1e-06 
3.0 2.395 0 -3.0 1e-06 
0.05 2.396 0 -3.0 1e-06 
3.0 2.396 0 -3.0 1e-06 
0.05 2.397 0 -3.0 1e-06 
3.0 2.397 0 -3.0 1e-06 
0.05 2.398 0 -3.0 1e-06 
3.0 2.398 0 -3.0 1e-06 
0.05 2.399 0 -3.0 1e-06 
3.0 2.399 0 -3.0 1e-06 
0.05 2.4 0 -3.0 1e-06 
3.0 2.4 0 -3.0 1e-06 
0.05 2.401 0 -3.0 1e-06 
3.0 2.401 0 -3.0 1e-06 
0.05 2.402 0 -3.0 1e-06 
3.0 2.402 0 -3.0 1e-06 
0.05 2.403 0 -3.0 1e-06 
3.0 2.403 0 -3.0 1e-06 
0.05 2.404 0 -3.0 1e-06 
3.0 2.404 0 -3.0 1e-06 
0.05 2.405 0 -3.0 1e-06 
3.0 2.405 0 -3.0 1e-06 
0.05 2.406 0 -3.0 1e-06 
3.0 2.406 0 -3.0 1e-06 
0.05 2.407 0 -3.0 1e-06 
3.0 2.407 0 -3.0 1e-06 
0.05 2.408 0 -3.0 1e-06 
3.0 2.408 0 -3.0 1e-06 
0.05 2.409 0 -3.0 1e-06 
3.0 2.409 0 -3.0 1e-06 
0.05 2.41 0 -3.0 1e-06 
3.0 2.41 0 -3.0 1e-06 
0.05 2.411 0 -3.0 1e-06 
3.0 2.411 0 -3.0 1e-06 
0.05 2.412 0 -3.0 1e-06 
3.0 2.412 0 -3.0 1e-06 
0.05 2.413 0 -3.0 1e-06 
3.0 2.413 0 -3.0 1e-06 
0.05 2.414 0 -3.0 1e-06 
3.0 2.414 0 -3.0 1e-06 
0.05 2.415 0 -3.0 1e-06 
3.0 2.415 0 -3.0 1e-06 
0.05 2.416 0 -3.0 1e-06 
3.0 2.416 0 -3.0 1e-06 
0.05 2.417 0 -3.0 1e-06 
3.0 2.417 0 -3.0 1e-06 
0.05 2.418 0 -3.0 1e-06 
3.0 2.418 0 -3.0 1e-06 
0.05 2.419 0 -3.0 1e-06 
3.0 2.419 0 -3.0 1e-06 
0.05 2.42 0 -3.0 1e-06 
3.0 2.42 0 -3.0 1e-06 
0.05 2.421 0 -3.0 1e-06 
3.0 2.421 0 -3.0 1e-06 
0.05 2.422 0 -3.0 1e-06 
3.0 2.422 0 -3.0 1e-06 
0.05 2.423 0 -3.0 1e-06 
3.0 2.423 0 -3.0 1e-06 
0.05 2.424 0 -3.0 1e-06 
3.0 2.424 0 -3.0 1e-06 
0.05 2.425 0 -3.0 1e-06 
3.0 2.425 0 -3.0 1e-06 
0.05 2.426 0 -3.0 1e-06 
3.0 2.426 0 -3.0 1e-06 
0.05 2.427 0 -3.0 1e-06 
3.0 2.427 0 -3.0 1e-06 
0.05 2.428 0 -3.0 1e-06 
3.0 2.428 0 -3.0 1e-06 
0.05 2.429 0 -3.0 1e-06 
3.0 2.429 0 -3.0 1e-06 
0.05 2.43 0 -3.0 1e-06 
3.0 2.43 0 -3.0 1e-06 
0.05 2.431 0 -3.0 1e-06 
3.0 2.431 0 -3.0 1e-06 
0.05 2.432 0 -3.0 1e-06 
3.0 2.432 0 -3.0 1e-06 
0.05 2.433 0 -3.0 1e-06 
3.0 2.433 0 -3.0 1e-06 
0.05 2.434 0 -3.0 1e-06 
3.0 2.434 0 -3.0 1e-06 
0.05 2.435 0 -3.0 1e-06 
3.0 2.435 0 -3.0 1e-06 
0.05 2.436 0 -3.0 1e-06 
3.0 2.436 0 -3.0 1e-06 
0.05 2.437 0 -3.0 1e-06 
3.0 2.437 0 -3.0 1e-06 
0.05 2.438 0 -3.0 1e-06 
3.0 2.438 0 -3.0 1e-06 
0.05 2.439 0 -3.0 1e-06 
3.0 2.439 0 -3.0 1e-06 
0.05 2.44 0 -3.0 1e-06 
3.0 2.44 0 -3.0 1e-06 
0.05 2.441 0 -3.0 1e-06 
3.0 2.441 0 -3.0 1e-06 
0.05 2.442 0 -3.0 1e-06 
3.0 2.442 0 -3.0 1e-06 
0.05 2.443 0 -3.0 1e-06 
3.0 2.443 0 -3.0 1e-06 
0.05 2.444 0 -3.0 1e-06 
3.0 2.444 0 -3.0 1e-06 
0.05 2.445 0 -3.0 1e-06 
3.0 2.445 0 -3.0 1e-06 
0.05 2.446 0 -3.0 1e-06 
3.0 2.446 0 -3.0 1e-06 
0.05 2.447 0 -3.0 1e-06 
3.0 2.447 0 -3.0 1e-06 
0.05 2.448 0 -3.0 1e-06 
3.0 2.448 0 -3.0 1e-06 
0.05 2.449 0 -3.0 1e-06 
3.0 2.449 0 -3.0 1e-06 
0.05 2.45 0 -3.0 1e-06 
3.0 2.45 0 -3.0 1e-06 
0.05 2.451 0 -3.0 1e-06 
3.0 2.451 0 -3.0 1e-06 
0.05 2.452 0 -3.0 1e-06 
3.0 2.452 0 -3.0 1e-06 
0.05 2.453 0 -3.0 1e-06 
3.0 2.453 0 -3.0 1e-06 
0.05 2.454 0 -3.0 1e-06 
3.0 2.454 0 -3.0 1e-06 
0.05 2.455 0 -3.0 1e-06 
3.0 2.455 0 -3.0 1e-06 
0.05 2.456 0 -3.0 1e-06 
3.0 2.456 0 -3.0 1e-06 
0.05 2.457 0 -3.0 1e-06 
3.0 2.457 0 -3.0 1e-06 
0.05 2.458 0 -3.0 1e-06 
3.0 2.458 0 -3.0 1e-06 
0.05 2.459 0 -3.0 1e-06 
3.0 2.459 0 -3.0 1e-06 
0.05 2.46 0 -3.0 1e-06 
3.0 2.46 0 -3.0 1e-06 
0.05 2.461 0 -3.0 1e-06 
3.0 2.461 0 -3.0 1e-06 
0.05 2.462 0 -3.0 1e-06 
3.0 2.462 0 -3.0 1e-06 
0.05 2.463 0 -3.0 1e-06 
3.0 2.463 0 -3.0 1e-06 
0.05 2.464 0 -3.0 1e-06 
3.0 2.464 0 -3.0 1e-06 
0.05 2.465 0 -3.0 1e-06 
3.0 2.465 0 -3.0 1e-06 
0.05 2.466 0 -3.0 1e-06 
3.0 2.466 0 -3.0 1e-06 
0.05 2.467 0 -3.0 1e-06 
3.0 2.467 0 -3.0 1e-06 
0.05 2.468 0 -3.0 1e-06 
3.0 2.468 0 -3.0 1e-06 
0.05 2.469 0 -3.0 1e-06 
3.0 2.469 0 -3.0 1e-06 
0.05 2.47 0 -3.0 1e-06 
3.0 2.47 0 -3.0 1e-06 
0.05 2.471 0 -3.0 1e-06 
3.0 2.471 0 -3.0 1e-06 
0.05 2.472 0 -3.0 1e-06 
3.0 2.472 0 -3.0 1e-06 
0.05 2.473 0 -3.0 1e-06 
3.0 2.473 0 -3.0 1e-06 
0.05 2.474 0 -3.0 1e-06 
3.0 2.474 0 -3.0 1e-06 
0.05 2.475 0 -3.0 1e-06 
3.0 2.475 0 -3.0 1e-06 
0.05 2.476 0 -3.0 1e-06 
3.0 2.476 0 -3.0 1e-06 
0.05 2.477 0 -3.0 1e-06 
3.0 2.477 0 -3.0 1e-06 
0.05 2.478 0 -3.0 1e-06 
3.0 2.478 0 -3.0 1e-06 
0.05 2.479 0 -3.0 1e-06 
3.0 2.479 0 -3.0 1e-06 
0.05 2.48 0 -3.0 1e-06 
3.0 2.48 0 -3.0 1e-06 
0.05 2.481 0 -3.0 1e-06 
3.0 2.481 0 -3.0 1e-06 
0.05 2.482 0 -3.0 1e-06 
3.0 2.482 0 -3.0 1e-06 
0.05 2.483 0 -3.0 1e-06 
3.0 2.483 0 -3.0 1e-06 
0.05 2.484 0 -3.0 1e-06 
3.0 2.484 0 -3.0 1e-06 
0.05 2.485 0 -3.0 1e-06 
3.0 2.485 0 -3.0 1e-06 
0.05 2.486 0 -3.0 1e-06 
3.0 2.486 0 -3.0 1e-06 
0.05 2.487 0 -3.0 1e-06 
3.0 2.487 0 -3.0 1e-06 
0.05 2.488 0 -3.0 1e-06 
3.0 2.488 0 -3.0 1e-06 
0.05 2.489 0 -3.0 1e-06 
3.0 2.489 0 -3.0 1e-06 
0.05 2.49 0 -3.0 1e-06 
3.0 2.49 0 -3.0 1e-06 
0.05 2.491 0 -3.0 1e-06 
3.0 2.491 0 -3.0 1e-06 
0.05 2.492 0 -3.0 1e-06 
3.0 2.492 0 -3.0 1e-06 
0.05 2.493 0 -3.0 1e-06 
3.0 2.493 0 -3.0 1e-06 
0.05 2.494 0 -3.0 1e-06 
3.0 2.494 0 -3.0 1e-06 
0.05 2.495 0 -3.0 1e-06 
3.0 2.495 0 -3.0 1e-06 
0.05 2.496 0 -3.0 1e-06 
3.0 2.496 0 -3.0 1e-06 
0.05 2.497 0 -3.0 1e-06 
3.0 2.497 0 -3.0 1e-06 
0.05 2.498 0 -3.0 1e-06 
3.0 2.498 0 -3.0 1e-06 
0.05 2.499 0 -3.0 1e-06 
3.0 2.499 0 -3.0 1e-06 
0.05 2.5 0 -3.0 1e-06 
3.0 2.5 0 -3.0 1e-06 
0.05 2.501 0 -3.0 1e-06 
3.0 2.501 0 -3.0 1e-06 
0.05 2.502 0 -3.0 1e-06 
3.0 2.502 0 -3.0 1e-06 
0.05 2.503 0 -3.0 1e-06 
3.0 2.503 0 -3.0 1e-06 
0.05 2.504 0 -3.0 1e-06 
3.0 2.504 0 -3.0 1e-06 
0.05 2.505 0 -3.0 1e-06 
3.0 2.505 0 -3.0 1e-06 
0.05 2.506 0 -3.0 1e-06 
3.0 2.506 0 -3.0 1e-06 
0.05 2.507 0 -3.0 1e-06 
3.0 2.507 0 -3.0 1e-06 
0.05 2.508 0 -3.0 1e-06 
3.0 2.508 0 -3.0 1e-06 
0.05 2.509 0 -3.0 1e-06 
3.0 2.509 0 -3.0 1e-06 
0.05 2.51 0 -3.0 1e-06 
3.0 2.51 0 -3.0 1e-06 
0.05 2.511 0 -3.0 1e-06 
3.0 2.511 0 -3.0 1e-06 
0.05 2.512 0 -3.0 1e-06 
3.0 2.512 0 -3.0 1e-06 
0.05 2.513 0 -3.0 1e-06 
3.0 2.513 0 -3.0 1e-06 
0.05 2.514 0 -3.0 1e-06 
3.0 2.514 0 -3.0 1e-06 
0.05 2.515 0 -3.0 1e-06 
3.0 2.515 0 -3.0 1e-06 
0.05 2.516 0 -3.0 1e-06 
3.0 2.516 0 -3.0 1e-06 
0.05 2.517 0 -3.0 1e-06 
3.0 2.517 0 -3.0 1e-06 
0.05 2.518 0 -3.0 1e-06 
3.0 2.518 0 -3.0 1e-06 
0.05 2.519 0 -3.0 1e-06 
3.0 2.519 0 -3.0 1e-06 
0.05 2.52 0 -3.0 1e-06 
3.0 2.52 0 -3.0 1e-06 
0.05 2.521 0 -3.0 1e-06 
3.0 2.521 0 -3.0 1e-06 
0.05 2.522 0 -3.0 1e-06 
3.0 2.522 0 -3.0 1e-06 
0.05 2.523 0 -3.0 1e-06 
3.0 2.523 0 -3.0 1e-06 
0.05 2.524 0 -3.0 1e-06 
3.0 2.524 0 -3.0 1e-06 
0.05 2.525 0 -3.0 1e-06 
3.0 2.525 0 -3.0 1e-06 
0.05 2.526 0 -3.0 1e-06 
3.0 2.526 0 -3.0 1e-06 
0.05 2.527 0 -3.0 1e-06 
3.0 2.527 0 -3.0 1e-06 
0.05 2.528 0 -3.0 1e-06 
3.0 2.528 0 -3.0 1e-06 
0.05 2.529 0 -3.0 1e-06 
3.0 2.529 0 -3.0 1e-06 
0.05 2.53 0 -3.0 1e-06 
3.0 2.53 0 -3.0 1e-06 
0.05 2.531 0 -3.0 1e-06 
3.0 2.531 0 -3.0 1e-06 
0.05 2.532 0 -3.0 1e-06 
3.0 2.532 0 -3.0 1e-06 
0.05 2.533 0 -3.0 1e-06 
3.0 2.533 0 -3.0 1e-06 
0.05 2.534 0 -3.0 1e-06 
3.0 2.534 0 -3.0 1e-06 
0.05 2.535 0 -3.0 1e-06 
3.0 2.535 0 -3.0 1e-06 
0.05 2.536 0 -3.0 1e-06 
3.0 2.536 0 -3.0 1e-06 
0.05 2.537 0 -3.0 1e-06 
3.0 2.537 0 -3.0 1e-06 
0.05 2.538 0 -3.0 1e-06 
3.0 2.538 0 -3.0 1e-06 
0.05 2.539 0 -3.0 1e-06 
3.0 2.539 0 -3.0 1e-06 
0.05 2.54 0 -3.0 1e-06 
3.0 2.54 0 -3.0 1e-06 
0.05 2.541 0 -3.0 1e-06 
3.0 2.541 0 -3.0 1e-06 
0.05 2.542 0 -3.0 1e-06 
3.0 2.542 0 -3.0 1e-06 
0.05 2.543 0 -3.0 1e-06 
3.0 2.543 0 -3.0 1e-06 
0.05 2.544 0 -3.0 1e-06 
3.0 2.544 0 -3.0 1e-06 
0.05 2.545 0 -3.0 1e-06 
3.0 2.545 0 -3.0 1e-06 
0.05 2.546 0 -3.0 1e-06 
3.0 2.546 0 -3.0 1e-06 
0.05 2.547 0 -3.0 1e-06 
3.0 2.547 0 -3.0 1e-06 
0.05 2.548 0 -3.0 1e-06 
3.0 2.548 0 -3.0 1e-06 
0.05 2.549 0 -3.0 1e-06 
3.0 2.549 0 -3.0 1e-06 
0.05 2.55 0 -3.0 1e-06 
3.0 2.55 0 -3.0 1e-06 
0.05 2.551 0 -3.0 1e-06 
3.0 2.551 0 -3.0 1e-06 
0.05 2.552 0 -3.0 1e-06 
3.0 2.552 0 -3.0 1e-06 
0.05 2.553 0 -3.0 1e-06 
3.0 2.553 0 -3.0 1e-06 
0.05 2.554 0 -3.0 1e-06 
3.0 2.554 0 -3.0 1e-06 
0.05 2.555 0 -3.0 1e-06 
3.0 2.555 0 -3.0 1e-06 
0.05 2.556 0 -3.0 1e-06 
3.0 2.556 0 -3.0 1e-06 
0.05 2.557 0 -3.0 1e-06 
3.0 2.557 0 -3.0 1e-06 
0.05 2.558 0 -3.0 1e-06 
3.0 2.558 0 -3.0 1e-06 
0.05 2.559 0 -3.0 1e-06 
3.0 2.559 0 -3.0 1e-06 
0.05 2.56 0 -3.0 1e-06 
3.0 2.56 0 -3.0 1e-06 
0.05 2.561 0 -3.0 1e-06 
3.0 2.561 0 -3.0 1e-06 
0.05 2.562 0 -3.0 1e-06 
3.0 2.562 0 -3.0 1e-06 
0.05 2.563 0 -3.0 1e-06 
3.0 2.563 0 -3.0 1e-06 
0.05 2.564 0 -3.0 1e-06 
3.0 2.564 0 -3.0 1e-06 
0.05 2.565 0 -3.0 1e-06 
3.0 2.565 0 -3.0 1e-06 
0.05 2.566 0 -3.0 1e-06 
3.0 2.566 0 -3.0 1e-06 
0.05 2.567 0 -3.0 1e-06 
3.0 2.567 0 -3.0 1e-06 
0.05 2.568 0 -3.0 1e-06 
3.0 2.568 0 -3.0 1e-06 
0.05 2.569 0 -3.0 1e-06 
3.0 2.569 0 -3.0 1e-06 
0.05 2.57 0 -3.0 1e-06 
3.0 2.57 0 -3.0 1e-06 
0.05 2.571 0 -3.0 1e-06 
3.0 2.571 0 -3.0 1e-06 
0.05 2.572 0 -3.0 1e-06 
3.0 2.572 0 -3.0 1e-06 
0.05 2.573 0 -3.0 1e-06 
3.0 2.573 0 -3.0 1e-06 
0.05 2.574 0 -3.0 1e-06 
3.0 2.574 0 -3.0 1e-06 
0.05 2.575 0 -3.0 1e-06 
3.0 2.575 0 -3.0 1e-06 
0.05 2.576 0 -3.0 1e-06 
3.0 2.576 0 -3.0 1e-06 
0.05 2.577 0 -3.0 1e-06 
3.0 2.577 0 -3.0 1e-06 
0.05 2.578 0 -3.0 1e-06 
3.0 2.578 0 -3.0 1e-06 
0.05 2.579 0 -3.0 1e-06 
3.0 2.579 0 -3.0 1e-06 
0.05 2.58 0 -3.0 1e-06 
3.0 2.58 0 -3.0 1e-06 
0.05 2.581 0 -3.0 1e-06 
3.0 2.581 0 -3.0 1e-06 
0.05 2.582 0 -3.0 1e-06 
3.0 2.582 0 -3.0 1e-06 
0.05 2.583 0 -3.0 1e-06 
3.0 2.583 0 -3.0 1e-06 
0.05 2.584 0 -3.0 1e-06 
3.0 2.584 0 -3.0 1e-06 
0.05 2.585 0 -3.0 1e-06 
3.0 2.585 0 -3.0 1e-06 
0.05 2.586 0 -3.0 1e-06 
3.0 2.586 0 -3.0 1e-06 
0.05 2.587 0 -3.0 1e-06 
3.0 2.587 0 -3.0 1e-06 
0.05 2.588 0 -3.0 1e-06 
3.0 2.588 0 -3.0 1e-06 
0.05 2.589 0 -3.0 1e-06 
3.0 2.589 0 -3.0 1e-06 
0.05 2.59 0 -3.0 1e-06 
3.0 2.59 0 -3.0 1e-06 
0.05 2.591 0 -3.0 1e-06 
3.0 2.591 0 -3.0 1e-06 
0.05 2.592 0 -3.0 1e-06 
3.0 2.592 0 -3.0 1e-06 
0.05 2.593 0 -3.0 1e-06 
3.0 2.593 0 -3.0 1e-06 
0.05 2.594 0 -3.0 1e-06 
3.0 2.594 0 -3.0 1e-06 
0.05 2.595 0 -3.0 1e-06 
3.0 2.595 0 -3.0 1e-06 
0.05 2.596 0 -3.0 1e-06 
3.0 2.596 0 -3.0 1e-06 
0.05 2.597 0 -3.0 1e-06 
3.0 2.597 0 -3.0 1e-06 
0.05 2.598 0 -3.0 1e-06 
3.0 2.598 0 -3.0 1e-06 
0.05 2.599 0 -3.0 1e-06 
3.0 2.599 0 -3.0 1e-06 
0.05 2.6 0 -3.0 1e-06 
3.0 2.6 0 -3.0 1e-06 
0.05 2.601 0 -3.0 1e-06 
3.0 2.601 0 -3.0 1e-06 
0.05 2.602 0 -3.0 1e-06 
3.0 2.602 0 -3.0 1e-06 
0.05 2.603 0 -3.0 1e-06 
3.0 2.603 0 -3.0 1e-06 
0.05 2.604 0 -3.0 1e-06 
3.0 2.604 0 -3.0 1e-06 
0.05 2.605 0 -3.0 1e-06 
3.0 2.605 0 -3.0 1e-06 
0.05 2.606 0 -3.0 1e-06 
3.0 2.606 0 -3.0 1e-06 
0.05 2.607 0 -3.0 1e-06 
3.0 2.607 0 -3.0 1e-06 
0.05 2.608 0 -3.0 1e-06 
3.0 2.608 0 -3.0 1e-06 
0.05 2.609 0 -3.0 1e-06 
3.0 2.609 0 -3.0 1e-06 
0.05 2.61 0 -3.0 1e-06 
3.0 2.61 0 -3.0 1e-06 
0.05 2.611 0 -3.0 1e-06 
3.0 2.611 0 -3.0 1e-06 
0.05 2.612 0 -3.0 1e-06 
3.0 2.612 0 -3.0 1e-06 
0.05 2.613 0 -3.0 1e-06 
3.0 2.613 0 -3.0 1e-06 
0.05 2.614 0 -3.0 1e-06 
3.0 2.614 0 -3.0 1e-06 
0.05 2.615 0 -3.0 1e-06 
3.0 2.615 0 -3.0 1e-06 
0.05 2.616 0 -3.0 1e-06 
3.0 2.616 0 -3.0 1e-06 
0.05 2.617 0 -3.0 1e-06 
3.0 2.617 0 -3.0 1e-06 
0.05 2.618 0 -3.0 1e-06 
3.0 2.618 0 -3.0 1e-06 
0.05 2.619 0 -3.0 1e-06 
3.0 2.619 0 -3.0 1e-06 
0.05 2.62 0 -3.0 1e-06 
3.0 2.62 0 -3.0 1e-06 
0.05 2.621 0 -3.0 1e-06 
3.0 2.621 0 -3.0 1e-06 
0.05 2.622 0 -3.0 1e-06 
3.0 2.622 0 -3.0 1e-06 
0.05 2.623 0 -3.0 1e-06 
3.0 2.623 0 -3.0 1e-06 
0.05 2.624 0 -3.0 1e-06 
3.0 2.624 0 -3.0 1e-06 
0.05 2.625 0 -3.0 1e-06 
3.0 2.625 0 -3.0 1e-06 
0.05 2.626 0 -3.0 1e-06 
3.0 2.626 0 -3.0 1e-06 
0.05 2.627 0 -3.0 1e-06 
3.0 2.627 0 -3.0 1e-06 
0.05 2.628 0 -3.0 1e-06 
3.0 2.628 0 -3.0 1e-06 
0.05 2.629 0 -3.0 1e-06 
3.0 2.629 0 -3.0 1e-06 
0.05 2.63 0 -3.0 1e-06 
3.0 2.63 0 -3.0 1e-06 
0.05 2.631 0 -3.0 1e-06 
3.0 2.631 0 -3.0 1e-06 
0.05 2.632 0 -3.0 1e-06 
3.0 2.632 0 -3.0 1e-06 
0.05 2.633 0 -3.0 1e-06 
3.0 2.633 0 -3.0 1e-06 
0.05 2.634 0 -3.0 1e-06 
3.0 2.634 0 -3.0 1e-06 
0.05 2.635 0 -3.0 1e-06 
3.0 2.635 0 -3.0 1e-06 
0.05 2.636 0 -3.0 1e-06 
3.0 2.636 0 -3.0 1e-06 
0.05 2.637 0 -3.0 1e-06 
3.0 2.637 0 -3.0 1e-06 
0.05 2.638 0 -3.0 1e-06 
3.0 2.638 0 -3.0 1e-06 
0.05 2.639 0 -3.0 1e-06 
3.0 2.639 0 -3.0 1e-06 
0.05 2.64 0 -3.0 1e-06 
3.0 2.64 0 -3.0 1e-06 
0.05 2.641 0 -3.0 1e-06 
3.0 2.641 0 -3.0 1e-06 
0.05 2.642 0 -3.0 1e-06 
3.0 2.642 0 -3.0 1e-06 
0.05 2.643 0 -3.0 1e-06 
3.0 2.643 0 -3.0 1e-06 
0.05 2.644 0 -3.0 1e-06 
3.0 2.644 0 -3.0 1e-06 
0.05 2.645 0 -3.0 1e-06 
3.0 2.645 0 -3.0 1e-06 
0.05 2.646 0 -3.0 1e-06 
3.0 2.646 0 -3.0 1e-06 
0.05 2.647 0 -3.0 1e-06 
3.0 2.647 0 -3.0 1e-06 
0.05 2.648 0 -3.0 1e-06 
3.0 2.648 0 -3.0 1e-06 
0.05 2.649 0 -3.0 1e-06 
3.0 2.649 0 -3.0 1e-06 
0.05 2.65 0 -3.0 1e-06 
3.0 2.65 0 -3.0 1e-06 
0.05 2.651 0 -3.0 1e-06 
3.0 2.651 0 -3.0 1e-06 
0.05 2.652 0 -3.0 1e-06 
3.0 2.652 0 -3.0 1e-06 
0.05 2.653 0 -3.0 1e-06 
3.0 2.653 0 -3.0 1e-06 
0.05 2.654 0 -3.0 1e-06 
3.0 2.654 0 -3.0 1e-06 
0.05 2.655 0 -3.0 1e-06 
3.0 2.655 0 -3.0 1e-06 
0.05 2.656 0 -3.0 1e-06 
3.0 2.656 0 -3.0 1e-06 
0.05 2.657 0 -3.0 1e-06 
3.0 2.657 0 -3.0 1e-06 
0.05 2.658 0 -3.0 1e-06 
3.0 2.658 0 -3.0 1e-06 
0.05 2.659 0 -3.0 1e-06 
3.0 2.659 0 -3.0 1e-06 
0.05 2.66 0 -3.0 1e-06 
3.0 2.66 0 -3.0 1e-06 
0.05 2.661 0 -3.0 1e-06 
3.0 2.661 0 -3.0 1e-06 
0.05 2.662 0 -3.0 1e-06 
3.0 2.662 0 -3.0 1e-06 
0.05 2.663 0 -3.0 1e-06 
3.0 2.663 0 -3.0 1e-06 
0.05 2.664 0 -3.0 1e-06 
3.0 2.664 0 -3.0 1e-06 
0.05 2.665 0 -3.0 1e-06 
3.0 2.665 0 -3.0 1e-06 
0.05 2.666 0 -3.0 1e-06 
3.0 2.666 0 -3.0 1e-06 
0.05 2.667 0 -3.0 1e-06 
3.0 2.667 0 -3.0 1e-06 
0.05 2.668 0 -3.0 1e-06 
3.0 2.668 0 -3.0 1e-06 
0.05 2.669 0 -3.0 1e-06 
3.0 2.669 0 -3.0 1e-06 
0.05 2.67 0 -3.0 1e-06 
3.0 2.67 0 -3.0 1e-06 
0.05 2.671 0 -3.0 1e-06 
3.0 2.671 0 -3.0 1e-06 
0.05 2.672 0 -3.0 1e-06 
3.0 2.672 0 -3.0 1e-06 
0.05 2.673 0 -3.0 1e-06 
3.0 2.673 0 -3.0 1e-06 
0.05 2.674 0 -3.0 1e-06 
3.0 2.674 0 -3.0 1e-06 
0.05 2.675 0 -3.0 1e-06 
3.0 2.675 0 -3.0 1e-06 
0.05 2.676 0 -3.0 1e-06 
3.0 2.676 0 -3.0 1e-06 
0.05 2.677 0 -3.0 1e-06 
3.0 2.677 0 -3.0 1e-06 
0.05 2.678 0 -3.0 1e-06 
3.0 2.678 0 -3.0 1e-06 
0.05 2.679 0 -3.0 1e-06 
3.0 2.679 0 -3.0 1e-06 
0.05 2.68 0 -3.0 1e-06 
3.0 2.68 0 -3.0 1e-06 
0.05 2.681 0 -3.0 1e-06 
3.0 2.681 0 -3.0 1e-06 
0.05 2.682 0 -3.0 1e-06 
3.0 2.682 0 -3.0 1e-06 
0.05 2.683 0 -3.0 1e-06 
3.0 2.683 0 -3.0 1e-06 
0.05 2.684 0 -3.0 1e-06 
3.0 2.684 0 -3.0 1e-06 
0.05 2.685 0 -3.0 1e-06 
3.0 2.685 0 -3.0 1e-06 
0.05 2.686 0 -3.0 1e-06 
3.0 2.686 0 -3.0 1e-06 
0.05 2.687 0 -3.0 1e-06 
3.0 2.687 0 -3.0 1e-06 
0.05 2.688 0 -3.0 1e-06 
3.0 2.688 0 -3.0 1e-06 
0.05 2.689 0 -3.0 1e-06 
3.0 2.689 0 -3.0 1e-06 
0.05 2.69 0 -3.0 1e-06 
3.0 2.69 0 -3.0 1e-06 
0.05 2.691 0 -3.0 1e-06 
3.0 2.691 0 -3.0 1e-06 
0.05 2.692 0 -3.0 1e-06 
3.0 2.692 0 -3.0 1e-06 
0.05 2.693 0 -3.0 1e-06 
3.0 2.693 0 -3.0 1e-06 
0.05 2.694 0 -3.0 1e-06 
3.0 2.694 0 -3.0 1e-06 
0.05 2.695 0 -3.0 1e-06 
3.0 2.695 0 -3.0 1e-06 
0.05 2.696 0 -3.0 1e-06 
3.0 2.696 0 -3.0 1e-06 
0.05 2.697 0 -3.0 1e-06 
3.0 2.697 0 -3.0 1e-06 
0.05 2.698 0 -3.0 1e-06 
3.0 2.698 0 -3.0 1e-06 
0.05 2.699 0 -3.0 1e-06 
3.0 2.699 0 -3.0 1e-06 
0.05 2.7 0 -3.0 1e-06 
3.0 2.7 0 -3.0 1e-06 
0.05 2.701 0 -3.0 1e-06 
3.0 2.701 0 -3.0 1e-06 
0.05 2.702 0 -3.0 1e-06 
3.0 2.702 0 -3.0 1e-06 
0.05 2.703 0 -3.0 1e-06 
3.0 2.703 0 -3.0 1e-06 
0.05 2.704 0 -3.0 1e-06 
3.0 2.704 0 -3.0 1e-06 
0.05 2.705 0 -3.0 1e-06 
3.0 2.705 0 -3.0 1e-06 
0.05 2.706 0 -3.0 1e-06 
3.0 2.706 0 -3.0 1e-06 
0.05 2.707 0 -3.0 1e-06 
3.0 2.707 0 -3.0 1e-06 
0.05 2.708 0 -3.0 1e-06 
3.0 2.708 0 -3.0 1e-06 
0.05 2.709 0 -3.0 1e-06 
3.0 2.709 0 -3.0 1e-06 
0.05 2.71 0 -3.0 1e-06 
3.0 2.71 0 -3.0 1e-06 
0.05 2.711 0 -3.0 1e-06 
3.0 2.711 0 -3.0 1e-06 
0.05 2.712 0 -3.0 1e-06 
3.0 2.712 0 -3.0 1e-06 
0.05 2.713 0 -3.0 1e-06 
3.0 2.713 0 -3.0 1e-06 
0.05 2.714 0 -3.0 1e-06 
3.0 2.714 0 -3.0 1e-06 
0.05 2.715 0 -3.0 1e-06 
3.0 2.715 0 -3.0 1e-06 
0.05 2.716 0 -3.0 1e-06 
3.0 2.716 0 -3.0 1e-06 
0.05 2.717 0 -3.0 1e-06 
3.0 2.717 0 -3.0 1e-06 
0.05 2.718 0 -3.0 1e-06 
3.0 2.718 0 -3.0 1e-06 
0.05 2.719 0 -3.0 1e-06 
3.0 2.719 0 -3.0 1e-06 
0.05 2.72 0 -3.0 1e-06 
3.0 2.72 0 -3.0 1e-06 
0.05 2.721 0 -3.0 1e-06 
3.0 2.721 0 -3.0 1e-06 
0.05 2.722 0 -3.0 1e-06 
3.0 2.722 0 -3.0 1e-06 
0.05 2.723 0 -3.0 1e-06 
3.0 2.723 0 -3.0 1e-06 
0.05 2.724 0 -3.0 1e-06 
3.0 2.724 0 -3.0 1e-06 
0.05 2.725 0 -3.0 1e-06 
3.0 2.725 0 -3.0 1e-06 
0.05 2.726 0 -3.0 1e-06 
3.0 2.726 0 -3.0 1e-06 
0.05 2.727 0 -3.0 1e-06 
3.0 2.727 0 -3.0 1e-06 
0.05 2.728 0 -3.0 1e-06 
3.0 2.728 0 -3.0 1e-06 
0.05 2.729 0 -3.0 1e-06 
3.0 2.729 0 -3.0 1e-06 
0.05 2.73 0 -3.0 1e-06 
3.0 2.73 0 -3.0 1e-06 
0.05 2.731 0 -3.0 1e-06 
3.0 2.731 0 -3.0 1e-06 
0.05 2.732 0 -3.0 1e-06 
3.0 2.732 0 -3.0 1e-06 
0.05 2.733 0 -3.0 1e-06 
3.0 2.733 0 -3.0 1e-06 
0.05 2.734 0 -3.0 1e-06 
3.0 2.734 0 -3.0 1e-06 
0.05 2.735 0 -3.0 1e-06 
3.0 2.735 0 -3.0 1e-06 
0.05 2.736 0 -3.0 1e-06 
3.0 2.736 0 -3.0 1e-06 
0.05 2.737 0 -3.0 1e-06 
3.0 2.737 0 -3.0 1e-06 
0.05 2.738 0 -3.0 1e-06 
3.0 2.738 0 -3.0 1e-06 
0.05 2.739 0 -3.0 1e-06 
3.0 2.739 0 -3.0 1e-06 
0.05 2.74 0 -3.0 1e-06 
3.0 2.74 0 -3.0 1e-06 
0.05 2.741 0 -3.0 1e-06 
3.0 2.741 0 -3.0 1e-06 
0.05 2.742 0 -3.0 1e-06 
3.0 2.742 0 -3.0 1e-06 
0.05 2.743 0 -3.0 1e-06 
3.0 2.743 0 -3.0 1e-06 
0.05 2.744 0 -3.0 1e-06 
3.0 2.744 0 -3.0 1e-06 
0.05 2.745 0 -3.0 1e-06 
3.0 2.745 0 -3.0 1e-06 
0.05 2.746 0 -3.0 1e-06 
3.0 2.746 0 -3.0 1e-06 
0.05 2.747 0 -3.0 1e-06 
3.0 2.747 0 -3.0 1e-06 
0.05 2.748 0 -3.0 1e-06 
3.0 2.748 0 -3.0 1e-06 
0.05 2.749 0 -3.0 1e-06 
3.0 2.749 0 -3.0 1e-06 
0.05 2.75 0 -3.0 1e-06 
3.0 2.75 0 -3.0 1e-06 
0.05 2.751 0 -3.0 1e-06 
3.0 2.751 0 -3.0 1e-06 
0.05 2.752 0 -3.0 1e-06 
3.0 2.752 0 -3.0 1e-06 
0.05 2.753 0 -3.0 1e-06 
3.0 2.753 0 -3.0 1e-06 
0.05 2.754 0 -3.0 1e-06 
3.0 2.754 0 -3.0 1e-06 
0.05 2.755 0 -3.0 1e-06 
3.0 2.755 0 -3.0 1e-06 
0.05 2.756 0 -3.0 1e-06 
3.0 2.756 0 -3.0 1e-06 
0.05 2.757 0 -3.0 1e-06 
3.0 2.757 0 -3.0 1e-06 
0.05 2.758 0 -3.0 1e-06 
3.0 2.758 0 -3.0 1e-06 
0.05 2.759 0 -3.0 1e-06 
3.0 2.759 0 -3.0 1e-06 
0.05 2.76 0 -3.0 1e-06 
3.0 2.76 0 -3.0 1e-06 
0.05 2.761 0 -3.0 1e-06 
3.0 2.761 0 -3.0 1e-06 
0.05 2.762 0 -3.0 1e-06 
3.0 2.762 0 -3.0 1e-06 
0.05 2.763 0 -3.0 1e-06 
3.0 2.763 0 -3.0 1e-06 
0.05 2.764 0 -3.0 1e-06 
3.0 2.764 0 -3.0 1e-06 
0.05 2.765 0 -3.0 1e-06 
3.0 2.765 0 -3.0 1e-06 
0.05 2.766 0 -3.0 1e-06 
3.0 2.766 0 -3.0 1e-06 
0.05 2.767 0 -3.0 1e-06 
3.0 2.767 0 -3.0 1e-06 
0.05 2.768 0 -3.0 1e-06 
3.0 2.768 0 -3.0 1e-06 
0.05 2.769 0 -3.0 1e-06 
3.0 2.769 0 -3.0 1e-06 
0.05 2.77 0 -3.0 1e-06 
3.0 2.77 0 -3.0 1e-06 
0.05 2.771 0 -3.0 1e-06 
3.0 2.771 0 -3.0 1e-06 
0.05 2.772 0 -3.0 1e-06 
3.0 2.772 0 -3.0 1e-06 
0.05 2.773 0 -3.0 1e-06 
3.0 2.773 0 -3.0 1e-06 
0.05 2.774 0 -3.0 1e-06 
3.0 2.774 0 -3.0 1e-06 
0.05 2.775 0 -3.0 1e-06 
3.0 2.775 0 -3.0 1e-06 
0.05 2.776 0 -3.0 1e-06 
3.0 2.776 0 -3.0 1e-06 
0.05 2.777 0 -3.0 1e-06 
3.0 2.777 0 -3.0 1e-06 
0.05 2.778 0 -3.0 1e-06 
3.0 2.778 0 -3.0 1e-06 
0.05 2.779 0 -3.0 1e-06 
3.0 2.779 0 -3.0 1e-06 
0.05 2.78 0 -3.0 1e-06 
3.0 2.78 0 -3.0 1e-06 
0.05 2.781 0 -3.0 1e-06 
3.0 2.781 0 -3.0 1e-06 
0.05 2.782 0 -3.0 1e-06 
3.0 2.782 0 -3.0 1e-06 
0.05 2.783 0 -3.0 1e-06 
3.0 2.783 0 -3.0 1e-06 
0.05 2.784 0 -3.0 1e-06 
3.0 2.784 0 -3.0 1e-06 
0.05 2.785 0 -3.0 1e-06 
3.0 2.785 0 -3.0 1e-06 
0.05 2.786 0 -3.0 1e-06 
3.0 2.786 0 -3.0 1e-06 
0.05 2.787 0 -3.0 1e-06 
3.0 2.787 0 -3.0 1e-06 
0.05 2.788 0 -3.0 1e-06 
3.0 2.788 0 -3.0 1e-06 
0.05 2.789 0 -3.0 1e-06 
3.0 2.789 0 -3.0 1e-06 
0.05 2.79 0 -3.0 1e-06 
3.0 2.79 0 -3.0 1e-06 
0.05 2.791 0 -3.0 1e-06 
3.0 2.791 0 -3.0 1e-06 
0.05 2.792 0 -3.0 1e-06 
3.0 2.792 0 -3.0 1e-06 
0.05 2.793 0 -3.0 1e-06 
3.0 2.793 0 -3.0 1e-06 
0.05 2.794 0 -3.0 1e-06 
3.0 2.794 0 -3.0 1e-06 
0.05 2.795 0 -3.0 1e-06 
3.0 2.795 0 -3.0 1e-06 
0.05 2.796 0 -3.0 1e-06 
3.0 2.796 0 -3.0 1e-06 
0.05 2.797 0 -3.0 1e-06 
3.0 2.797 0 -3.0 1e-06 
0.05 2.798 0 -3.0 1e-06 
3.0 2.798 0 -3.0 1e-06 
0.05 2.799 0 -3.0 1e-06 
3.0 2.799 0 -3.0 1e-06 
0.05 2.8 0 -3.0 1e-06 
3.0 2.8 0 -3.0 1e-06 
0.05 2.801 0 -3.0 1e-06 
3.0 2.801 0 -3.0 1e-06 
0.05 2.802 0 -3.0 1e-06 
3.0 2.802 0 -3.0 1e-06 
0.05 2.803 0 -3.0 1e-06 
3.0 2.803 0 -3.0 1e-06 
0.05 2.804 0 -3.0 1e-06 
3.0 2.804 0 -3.0 1e-06 
0.05 2.805 0 -3.0 1e-06 
3.0 2.805 0 -3.0 1e-06 
0.05 2.806 0 -3.0 1e-06 
3.0 2.806 0 -3.0 1e-06 
0.05 2.807 0 -3.0 1e-06 
3.0 2.807 0 -3.0 1e-06 
0.05 2.808 0 -3.0 1e-06 
3.0 2.808 0 -3.0 1e-06 
0.05 2.809 0 -3.0 1e-06 
3.0 2.809 0 -3.0 1e-06 
0.05 2.81 0 -3.0 1e-06 
3.0 2.81 0 -3.0 1e-06 
0.05 2.811 0 -3.0 1e-06 
3.0 2.811 0 -3.0 1e-06 
0.05 2.812 0 -3.0 1e-06 
3.0 2.812 0 -3.0 1e-06 
0.05 2.813 0 -3.0 1e-06 
3.0 2.813 0 -3.0 1e-06 
0.05 2.814 0 -3.0 1e-06 
3.0 2.814 0 -3.0 1e-06 
0.05 2.815 0 -3.0 1e-06 
3.0 2.815 0 -3.0 1e-06 
0.05 2.816 0 -3.0 1e-06 
3.0 2.816 0 -3.0 1e-06 
0.05 2.817 0 -3.0 1e-06 
3.0 2.817 0 -3.0 1e-06 
0.05 2.818 0 -3.0 1e-06 
3.0 2.818 0 -3.0 1e-06 
0.05 2.819 0 -3.0 1e-06 
3.0 2.819 0 -3.0 1e-06 
0.05 2.82 0 -3.0 1e-06 
3.0 2.82 0 -3.0 1e-06 
0.05 2.821 0 -3.0 1e-06 
3.0 2.821 0 -3.0 1e-06 
0.05 2.822 0 -3.0 1e-06 
3.0 2.822 0 -3.0 1e-06 
0.05 2.823 0 -3.0 1e-06 
3.0 2.823 0 -3.0 1e-06 
0.05 2.824 0 -3.0 1e-06 
3.0 2.824 0 -3.0 1e-06 
0.05 2.825 0 -3.0 1e-06 
3.0 2.825 0 -3.0 1e-06 
0.05 2.826 0 -3.0 1e-06 
3.0 2.826 0 -3.0 1e-06 
0.05 2.827 0 -3.0 1e-06 
3.0 2.827 0 -3.0 1e-06 
0.05 2.828 0 -3.0 1e-06 
3.0 2.828 0 -3.0 1e-06 
0.05 2.829 0 -3.0 1e-06 
3.0 2.829 0 -3.0 1e-06 
0.05 2.83 0 -3.0 1e-06 
3.0 2.83 0 -3.0 1e-06 
0.05 2.831 0 -3.0 1e-06 
3.0 2.831 0 -3.0 1e-06 
0.05 2.832 0 -3.0 1e-06 
3.0 2.832 0 -3.0 1e-06 
0.05 2.833 0 -3.0 1e-06 
3.0 2.833 0 -3.0 1e-06 
0.05 2.834 0 -3.0 1e-06 
3.0 2.834 0 -3.0 1e-06 
0.05 2.835 0 -3.0 1e-06 
3.0 2.835 0 -3.0 1e-06 
0.05 2.836 0 -3.0 1e-06 
3.0 2.836 0 -3.0 1e-06 
0.05 2.837 0 -3.0 1e-06 
3.0 2.837 0 -3.0 1e-06 
0.05 2.838 0 -3.0 1e-06 
3.0 2.838 0 -3.0 1e-06 
0.05 2.839 0 -3.0 1e-06 
3.0 2.839 0 -3.0 1e-06 
0.05 2.84 0 -3.0 1e-06 
3.0 2.84 0 -3.0 1e-06 
0.05 2.841 0 -3.0 1e-06 
3.0 2.841 0 -3.0 1e-06 
0.05 2.842 0 -3.0 1e-06 
3.0 2.842 0 -3.0 1e-06 
0.05 2.843 0 -3.0 1e-06 
3.0 2.843 0 -3.0 1e-06 
0.05 2.844 0 -3.0 1e-06 
3.0 2.844 0 -3.0 1e-06 
0.05 2.845 0 -3.0 1e-06 
3.0 2.845 0 -3.0 1e-06 
0.05 2.846 0 -3.0 1e-06 
3.0 2.846 0 -3.0 1e-06 
0.05 2.847 0 -3.0 1e-06 
3.0 2.847 0 -3.0 1e-06 
0.05 2.848 0 -3.0 1e-06 
3.0 2.848 0 -3.0 1e-06 
0.05 2.849 0 -3.0 1e-06 
3.0 2.849 0 -3.0 1e-06 
0.05 2.85 0 -3.0 1e-06 
3.0 2.85 0 -3.0 1e-06 
0.05 2.851 0 -3.0 1e-06 
3.0 2.851 0 -3.0 1e-06 
0.05 2.852 0 -3.0 1e-06 
3.0 2.852 0 -3.0 1e-06 
0.05 2.853 0 -3.0 1e-06 
3.0 2.853 0 -3.0 1e-06 
0.05 2.854 0 -3.0 1e-06 
3.0 2.854 0 -3.0 1e-06 
0.05 2.855 0 -3.0 1e-06 
3.0 2.855 0 -3.0 1e-06 
0.05 2.856 0 -3.0 1e-06 
3.0 2.856 0 -3.0 1e-06 
0.05 2.857 0 -3.0 1e-06 
3.0 2.857 0 -3.0 1e-06 
0.05 2.858 0 -3.0 1e-06 
3.0 2.858 0 -3.0 1e-06 
0.05 2.859 0 -3.0 1e-06 
3.0 2.859 0 -3.0 1e-06 
0.05 2.86 0 -3.0 1e-06 
3.0 2.86 0 -3.0 1e-06 
0.05 2.861 0 -3.0 1e-06 
3.0 2.861 0 -3.0 1e-06 
0.05 2.862 0 -3.0 1e-06 
3.0 2.862 0 -3.0 1e-06 
0.05 2.863 0 -3.0 1e-06 
3.0 2.863 0 -3.0 1e-06 
0.05 2.864 0 -3.0 1e-06 
3.0 2.864 0 -3.0 1e-06 
0.05 2.865 0 -3.0 1e-06 
3.0 2.865 0 -3.0 1e-06 
0.05 2.866 0 -3.0 1e-06 
3.0 2.866 0 -3.0 1e-06 
0.05 2.867 0 -3.0 1e-06 
3.0 2.867 0 -3.0 1e-06 
0.05 2.868 0 -3.0 1e-06 
3.0 2.868 0 -3.0 1e-06 
0.05 2.869 0 -3.0 1e-06 
3.0 2.869 0 -3.0 1e-06 
0.05 2.87 0 -3.0 1e-06 
3.0 2.87 0 -3.0 1e-06 
0.05 2.871 0 -3.0 1e-06 
3.0 2.871 0 -3.0 1e-06 
0.05 2.872 0 -3.0 1e-06 
3.0 2.872 0 -3.0 1e-06 
0.05 2.873 0 -3.0 1e-06 
3.0 2.873 0 -3.0 1e-06 
0.05 2.874 0 -3.0 1e-06 
3.0 2.874 0 -3.0 1e-06 
0.05 2.875 0 -3.0 1e-06 
3.0 2.875 0 -3.0 1e-06 
0.05 2.876 0 -3.0 1e-06 
3.0 2.876 0 -3.0 1e-06 
0.05 2.877 0 -3.0 1e-06 
3.0 2.877 0 -3.0 1e-06 
0.05 2.878 0 -3.0 1e-06 
3.0 2.878 0 -3.0 1e-06 
0.05 2.879 0 -3.0 1e-06 
3.0 2.879 0 -3.0 1e-06 
0.05 2.88 0 -3.0 1e-06 
3.0 2.88 0 -3.0 1e-06 
0.05 2.881 0 -3.0 1e-06 
3.0 2.881 0 -3.0 1e-06 
0.05 2.882 0 -3.0 1e-06 
3.0 2.882 0 -3.0 1e-06 
0.05 2.883 0 -3.0 1e-06 
3.0 2.883 0 -3.0 1e-06 
0.05 2.884 0 -3.0 1e-06 
3.0 2.884 0 -3.0 1e-06 
0.05 2.885 0 -3.0 1e-06 
3.0 2.885 0 -3.0 1e-06 
0.05 2.886 0 -3.0 1e-06 
3.0 2.886 0 -3.0 1e-06 
0.05 2.887 0 -3.0 1e-06 
3.0 2.887 0 -3.0 1e-06 
0.05 2.888 0 -3.0 1e-06 
3.0 2.888 0 -3.0 1e-06 
0.05 2.889 0 -3.0 1e-06 
3.0 2.889 0 -3.0 1e-06 
0.05 2.89 0 -3.0 1e-06 
3.0 2.89 0 -3.0 1e-06 
0.05 2.891 0 -3.0 1e-06 
3.0 2.891 0 -3.0 1e-06 
0.05 2.892 0 -3.0 1e-06 
3.0 2.892 0 -3.0 1e-06 
0.05 2.893 0 -3.0 1e-06 
3.0 2.893 0 -3.0 1e-06 
0.05 2.894 0 -3.0 1e-06 
3.0 2.894 0 -3.0 1e-06 
0.05 2.895 0 -3.0 1e-06 
3.0 2.895 0 -3.0 1e-06 
0.05 2.896 0 -3.0 1e-06 
3.0 2.896 0 -3.0 1e-06 
0.05 2.897 0 -3.0 1e-06 
3.0 2.897 0 -3.0 1e-06 
0.05 2.898 0 -3.0 1e-06 
3.0 2.898 0 -3.0 1e-06 
0.05 2.899 0 -3.0 1e-06 
3.0 2.899 0 -3.0 1e-06 
0.05 2.9 0 -3.0 1e-06 
3.0 2.9 0 -3.0 1e-06 
0.05 2.901 0 -3.0 1e-06 
3.0 2.901 0 -3.0 1e-06 
0.05 2.902 0 -3.0 1e-06 
3.0 2.902 0 -3.0 1e-06 
0.05 2.903 0 -3.0 1e-06 
3.0 2.903 0 -3.0 1e-06 
0.05 2.904 0 -3.0 1e-06 
3.0 2.904 0 -3.0 1e-06 
0.05 2.905 0 -3.0 1e-06 
3.0 2.905 0 -3.0 1e-06 
0.05 2.906 0 -3.0 1e-06 
3.0 2.906 0 -3.0 1e-06 
0.05 2.907 0 -3.0 1e-06 
3.0 2.907 0 -3.0 1e-06 
0.05 2.908 0 -3.0 1e-06 
3.0 2.908 0 -3.0 1e-06 
0.05 2.909 0 -3.0 1e-06 
3.0 2.909 0 -3.0 1e-06 
0.05 2.91 0 -3.0 1e-06 
3.0 2.91 0 -3.0 1e-06 
0.05 2.911 0 -3.0 1e-06 
3.0 2.911 0 -3.0 1e-06 
0.05 2.912 0 -3.0 1e-06 
3.0 2.912 0 -3.0 1e-06 
0.05 2.913 0 -3.0 1e-06 
3.0 2.913 0 -3.0 1e-06 
0.05 2.914 0 -3.0 1e-06 
3.0 2.914 0 -3.0 1e-06 
0.05 2.915 0 -3.0 1e-06 
3.0 2.915 0 -3.0 1e-06 
0.05 2.916 0 -3.0 1e-06 
3.0 2.916 0 -3.0 1e-06 
0.05 2.917 0 -3.0 1e-06 
3.0 2.917 0 -3.0 1e-06 
0.05 2.918 0 -3.0 1e-06 
3.0 2.918 0 -3.0 1e-06 
0.05 2.919 0 -3.0 1e-06 
3.0 2.919 0 -3.0 1e-06 
0.05 2.92 0 -3.0 1e-06 
3.0 2.92 0 -3.0 1e-06 
0.05 2.921 0 -3.0 1e-06 
3.0 2.921 0 -3.0 1e-06 
0.05 2.922 0 -3.0 1e-06 
3.0 2.922 0 -3.0 1e-06 
0.05 2.923 0 -3.0 1e-06 
3.0 2.923 0 -3.0 1e-06 
0.05 2.924 0 -3.0 1e-06 
3.0 2.924 0 -3.0 1e-06 
0.05 2.925 0 -3.0 1e-06 
3.0 2.925 0 -3.0 1e-06 
0.05 2.926 0 -3.0 1e-06 
3.0 2.926 0 -3.0 1e-06 
0.05 2.927 0 -3.0 1e-06 
3.0 2.927 0 -3.0 1e-06 
0.05 2.928 0 -3.0 1e-06 
3.0 2.928 0 -3.0 1e-06 
0.05 2.929 0 -3.0 1e-06 
3.0 2.929 0 -3.0 1e-06 
0.05 2.93 0 -3.0 1e-06 
3.0 2.93 0 -3.0 1e-06 
0.05 2.931 0 -3.0 1e-06 
3.0 2.931 0 -3.0 1e-06 
0.05 2.932 0 -3.0 1e-06 
3.0 2.932 0 -3.0 1e-06 
0.05 2.933 0 -3.0 1e-06 
3.0 2.933 0 -3.0 1e-06 
0.05 2.934 0 -3.0 1e-06 
3.0 2.934 0 -3.0 1e-06 
0.05 2.935 0 -3.0 1e-06 
3.0 2.935 0 -3.0 1e-06 
0.05 2.936 0 -3.0 1e-06 
3.0 2.936 0 -3.0 1e-06 
0.05 2.937 0 -3.0 1e-06 
3.0 2.937 0 -3.0 1e-06 
0.05 2.938 0 -3.0 1e-06 
3.0 2.938 0 -3.0 1e-06 
0.05 2.939 0 -3.0 1e-06 
3.0 2.939 0 -3.0 1e-06 
0.05 2.94 0 -3.0 1e-06 
3.0 2.94 0 -3.0 1e-06 
0.05 2.941 0 -3.0 1e-06 
3.0 2.941 0 -3.0 1e-06 
0.05 2.942 0 -3.0 1e-06 
3.0 2.942 0 -3.0 1e-06 
0.05 2.943 0 -3.0 1e-06 
3.0 2.943 0 -3.0 1e-06 
0.05 2.944 0 -3.0 1e-06 
3.0 2.944 0 -3.0 1e-06 
0.05 2.945 0 -3.0 1e-06 
3.0 2.945 0 -3.0 1e-06 
0.05 2.946 0 -3.0 1e-06 
3.0 2.946 0 -3.0 1e-06 
0.05 2.947 0 -3.0 1e-06 
3.0 2.947 0 -3.0 1e-06 
0.05 2.948 0 -3.0 1e-06 
3.0 2.948 0 -3.0 1e-06 
0.05 2.949 0 -3.0 1e-06 
3.0 2.949 0 -3.0 1e-06 
0.05 2.95 0 -3.0 1e-06 
3.0 2.95 0 -3.0 1e-06 
0.05 2.951 0 -3.0 1e-06 
3.0 2.951 0 -3.0 1e-06 
0.05 2.952 0 -3.0 1e-06 
3.0 2.952 0 -3.0 1e-06 
0.05 2.953 0 -3.0 1e-06 
3.0 2.953 0 -3.0 1e-06 
0.05 2.954 0 -3.0 1e-06 
3.0 2.954 0 -3.0 1e-06 
0.05 2.955 0 -3.0 1e-06 
3.0 2.955 0 -3.0 1e-06 
0.05 2.956 0 -3.0 1e-06 
3.0 2.956 0 -3.0 1e-06 
0.05 2.957 0 -3.0 1e-06 
3.0 2.957 0 -3.0 1e-06 
0.05 2.958 0 -3.0 1e-06 
3.0 2.958 0 -3.0 1e-06 
0.05 2.959 0 -3.0 1e-06 
3.0 2.959 0 -3.0 1e-06 
0.05 2.96 0 -3.0 1e-06 
3.0 2.96 0 -3.0 1e-06 
0.05 2.961 0 -3.0 1e-06 
3.0 2.961 0 -3.0 1e-06 
0.05 2.962 0 -3.0 1e-06 
3.0 2.962 0 -3.0 1e-06 
0.05 2.963 0 -3.0 1e-06 
3.0 2.963 0 -3.0 1e-06 
0.05 2.964 0 -3.0 1e-06 
3.0 2.964 0 -3.0 1e-06 
0.05 2.965 0 -3.0 1e-06 
3.0 2.965 0 -3.0 1e-06 
0.05 2.966 0 -3.0 1e-06 
3.0 2.966 0 -3.0 1e-06 
0.05 2.967 0 -3.0 1e-06 
3.0 2.967 0 -3.0 1e-06 
0.05 2.968 0 -3.0 1e-06 
3.0 2.968 0 -3.0 1e-06 
0.05 2.969 0 -3.0 1e-06 
3.0 2.969 0 -3.0 1e-06 
0.05 2.97 0 -3.0 1e-06 
3.0 2.97 0 -3.0 1e-06 
0.05 2.971 0 -3.0 1e-06 
3.0 2.971 0 -3.0 1e-06 
0.05 2.972 0 -3.0 1e-06 
3.0 2.972 0 -3.0 1e-06 
0.05 2.973 0 -3.0 1e-06 
3.0 2.973 0 -3.0 1e-06 
0.05 2.974 0 -3.0 1e-06 
3.0 2.974 0 -3.0 1e-06 
0.05 2.975 0 -3.0 1e-06 
3.0 2.975 0 -3.0 1e-06 
0.05 2.976 0 -3.0 1e-06 
3.0 2.976 0 -3.0 1e-06 
0.05 2.977 0 -3.0 1e-06 
3.0 2.977 0 -3.0 1e-06 
0.05 2.978 0 -3.0 1e-06 
3.0 2.978 0 -3.0 1e-06 
0.05 2.979 0 -3.0 1e-06 
3.0 2.979 0 -3.0 1e-06 
0.05 2.98 0 -3.0 1e-06 
3.0 2.98 0 -3.0 1e-06 
0.05 2.981 0 -3.0 1e-06 
3.0 2.981 0 -3.0 1e-06 
0.05 2.982 0 -3.0 1e-06 
3.0 2.982 0 -3.0 1e-06 
0.05 2.983 0 -3.0 1e-06 
3.0 2.983 0 -3.0 1e-06 
0.05 2.984 0 -3.0 1e-06 
3.0 2.984 0 -3.0 1e-06 
0.05 2.985 0 -3.0 1e-06 
3.0 2.985 0 -3.0 1e-06 
0.05 2.986 0 -3.0 1e-06 
3.0 2.986 0 -3.0 1e-06 
0.05 2.987 0 -3.0 1e-06 
3.0 2.987 0 -3.0 1e-06 
0.05 2.988 0 -3.0 1e-06 
3.0 2.988 0 -3.0 1e-06 
0.05 2.989 0 -3.0 1e-06 
3.0 2.989 0 -3.0 1e-06 
0.05 2.99 0 -3.0 1e-06 
3.0 2.99 0 -3.0 1e-06 
0.05 2.991 0 -3.0 1e-06 
3.0 2.991 0 -3.0 1e-06 
0.05 2.992 0 -3.0 1e-06 
3.0 2.992 0 -3.0 1e-06 
0.05 2.993 0 -3.0 1e-06 
3.0 2.993 0 -3.0 1e-06 
0.05 2.994 0 -3.0 1e-06 
3.0 2.994 0 -3.0 1e-06 
0.05 2.995 0 -3.0 1e-06 
3.0 2.995 0 -3.0 1e-06 
0.05 2.996 0 -3.0 1e-06 
3.0 2.996 0 -3.0 1e-06 
0.05 2.997 0 -3.0 1e-06 
3.0 2.997 0 -3.0 1e-06 
0.05 2.998 0 -3.0 1e-06 
3.0 2.998 0 -3.0 1e-06 
0.05 2.999 0 -3.0 1e-06 
3.0 2.999 0 -3.0 1e-06 
0.05 3.0 0 -3.0 1e-06 
3.0 3.0 0 -3.0 1e-06 
0.05 3.001 0 -3.0 1e-06 
3.0 3.001 0 -3.0 1e-06 
0.05 3.002 0 -3.0 1e-06 
3.0 3.002 0 -3.0 1e-06 
0.05 3.003 0 -3.0 1e-06 
3.0 3.003 0 -3.0 1e-06 
0.05 3.004 0 -3.0 1e-06 
3.0 3.004 0 -3.0 1e-06 
0.05 3.005 0 -3.0 1e-06 
3.0 3.005 0 -3.0 1e-06 
0.05 3.006 0 -3.0 1e-06 
3.0 3.006 0 -3.0 1e-06 
0.05 3.007 0 -3.0 1e-06 
3.0 3.007 0 -3.0 1e-06 
0.05 3.008 0 -3.0 1e-06 
3.0 3.008 0 -3.0 1e-06 
0.05 3.009 0 -3.0 1e-06 
3.0 3.009 0 -3.0 1e-06 
0.05 3.01 0 -3.0 1e-06 
3.0 3.01 0 -3.0 1e-06 
0.05 3.011 0 -3.0 1e-06 
3.0 3.011 0 -3.0 1e-06 
0.05 3.012 0 -3.0 1e-06 
3.0 3.012 0 -3.0 1e-06 
0.05 3.013 0 -3.0 1e-06 
3.0 3.013 0 -3.0 1e-06 
0.05 3.014 0 -3.0 1e-06 
3.0 3.014 0 -3.0 1e-06 
0.05 3.015 0 -3.0 1e-06 
3.0 3.015 0 -3.0 1e-06 
0.05 3.016 0 -3.0 1e-06 
3.0 3.016 0 -3.0 1e-06 
0.05 3.017 0 -3.0 1e-06 
3.0 3.017 0 -3.0 1e-06 
0.05 3.018 0 -3.0 1e-06 
3.0 3.018 0 -3.0 1e-06 
0.05 3.019 0 -3.0 1e-06 
3.0 3.019 0 -3.0 1e-06 
0.05 3.02 0 -3.0 1e-06 
3.0 3.02 0 -3.0 1e-06 
0.05 3.021 0 -3.0 1e-06 
3.0 3.021 0 -3.0 1e-06 
0.05 3.022 0 -3.0 1e-06 
3.0 3.022 0 -3.0 1e-06 
0.05 3.023 0 -3.0 1e-06 
3.0 3.023 0 -3.0 1e-06 
0.05 3.024 0 -3.0 1e-06 
3.0 3.024 0 -3.0 1e-06 
0.05 3.025 0 -3.0 1e-06 
3.0 3.025 0 -3.0 1e-06 
0.05 3.026 0 -3.0 1e-06 
3.0 3.026 0 -3.0 1e-06 
0.05 3.027 0 -3.0 1e-06 
3.0 3.027 0 -3.0 1e-06 
0.05 3.028 0 -3.0 1e-06 
3.0 3.028 0 -3.0 1e-06 
0.05 3.029 0 -3.0 1e-06 
3.0 3.029 0 -3.0 1e-06 
0.05 3.03 0 -3.0 1e-06 
3.0 3.03 0 -3.0 1e-06 
0.05 3.031 0 -3.0 1e-06 
3.0 3.031 0 -3.0 1e-06 
0.05 3.032 0 -3.0 1e-06 
3.0 3.032 0 -3.0 1e-06 
0.05 3.033 0 -3.0 1e-06 
3.0 3.033 0 -3.0 1e-06 
0.05 3.034 0 -3.0 1e-06 
3.0 3.034 0 -3.0 1e-06 
0.05 3.035 0 -3.0 1e-06 
3.0 3.035 0 -3.0 1e-06 
0.05 3.036 0 -3.0 1e-06 
3.0 3.036 0 -3.0 1e-06 
0.05 3.037 0 -3.0 1e-06 
3.0 3.037 0 -3.0 1e-06 
0.05 3.038 0 -3.0 1e-06 
3.0 3.038 0 -3.0 1e-06 
0.05 3.039 0 -3.0 1e-06 
3.0 3.039 0 -3.0 1e-06 
0.05 3.04 0 -3.0 1e-06 
3.0 3.04 0 -3.0 1e-06 
0.05 3.041 0 -3.0 1e-06 
3.0 3.041 0 -3.0 1e-06 
0.05 3.042 0 -3.0 1e-06 
3.0 3.042 0 -3.0 1e-06 
0.05 3.043 0 -3.0 1e-06 
3.0 3.043 0 -3.0 1e-06 
0.05 3.044 0 -3.0 1e-06 
3.0 3.044 0 -3.0 1e-06 
0.05 3.045 0 -3.0 1e-06 
3.0 3.045 0 -3.0 1e-06 
0.05 3.046 0 -3.0 1e-06 
3.0 3.046 0 -3.0 1e-06 
0.05 3.047 0 -3.0 1e-06 
3.0 3.047 0 -3.0 1e-06 
0.05 3.048 0 -3.0 1e-06 
3.0 3.048 0 -3.0 1e-06 
0.05 3.049 0 -3.0 1e-06 
3.0 3.049 0 -3.0 1e-06 
0.05 3.05 0 -3.0 1e-06 
3.0 3.05 0 -3.0 1e-06 
0.05 3.051 0 -3.0 1e-06 
3.0 3.051 0 -3.0 1e-06 
0.05 3.052 0 -3.0 1e-06 
3.0 3.052 0 -3.0 1e-06 
0.05 3.053 0 -3.0 1e-06 
3.0 3.053 0 -3.0 1e-06 
0.05 3.054 0 -3.0 1e-06 
3.0 3.054 0 -3.0 1e-06 
0.05 3.055 0 -3.0 1e-06 
3.0 3.055 0 -3.0 1e-06 
0.05 3.056 0 -3.0 1e-06 
3.0 3.056 0 -3.0 1e-06 
0.05 3.057 0 -3.0 1e-06 
3.0 3.057 0 -3.0 1e-06 
0.05 3.058 0 -3.0 1e-06 
3.0 3.058 0 -3.0 1e-06 
0.05 3.059 0 -3.0 1e-06 
3.0 3.059 0 -3.0 1e-06 
0.05 3.06 0 -3.0 1e-06 
3.0 3.06 0 -3.0 1e-06 
0.05 3.061 0 -3.0 1e-06 
3.0 3.061 0 -3.0 1e-06 
0.05 3.062 0 -3.0 1e-06 
3.0 3.062 0 -3.0 1e-06 
0.05 3.063 0 -3.0 1e-06 
3.0 3.063 0 -3.0 1e-06 
0.05 3.064 0 -3.0 1e-06 
3.0 3.064 0 -3.0 1e-06 
0.05 3.065 0 -3.0 1e-06 
3.0 3.065 0 -3.0 1e-06 
0.05 3.066 0 -3.0 1e-06 
3.0 3.066 0 -3.0 1e-06 
0.05 3.067 0 -3.0 1e-06 
3.0 3.067 0 -3.0 1e-06 
0.05 3.068 0 -3.0 1e-06 
3.0 3.068 0 -3.0 1e-06 
0.05 3.069 0 -3.0 1e-06 
3.0 3.069 0 -3.0 1e-06 
0.05 3.07 0 -3.0 1e-06 
3.0 3.07 0 -3.0 1e-06 
0.05 3.071 0 -3.0 1e-06 
3.0 3.071 0 -3.0 1e-06 
0.05 3.072 0 -3.0 1e-06 
3.0 3.072 0 -3.0 1e-06 
0.05 3.073 0 -3.0 1e-06 
3.0 3.073 0 -3.0 1e-06 
0.05 3.074 0 -3.0 1e-06 
3.0 3.074 0 -3.0 1e-06 
0.05 3.075 0 -3.0 1e-06 
3.0 3.075 0 -3.0 1e-06 
0.05 3.076 0 -3.0 1e-06 
3.0 3.076 0 -3.0 1e-06 
0.05 3.077 0 -3.0 1e-06 
3.0 3.077 0 -3.0 1e-06 
0.05 3.078 0 -3.0 1e-06 
3.0 3.078 0 -3.0 1e-06 
0.05 3.079 0 -3.0 1e-06 
3.0 3.079 0 -3.0 1e-06 
0.05 3.08 0 -3.0 1e-06 
3.0 3.08 0 -3.0 1e-06 
0.05 3.081 0 -3.0 1e-06 
3.0 3.081 0 -3.0 1e-06 
0.05 3.082 0 -3.0 1e-06 
3.0 3.082 0 -3.0 1e-06 
0.05 3.083 0 -3.0 1e-06 
3.0 3.083 0 -3.0 1e-06 
0.05 3.084 0 -3.0 1e-06 
3.0 3.084 0 -3.0 1e-06 
0.05 3.085 0 -3.0 1e-06 
3.0 3.085 0 -3.0 1e-06 
0.05 3.086 0 -3.0 1e-06 
3.0 3.086 0 -3.0 1e-06 
0.05 3.087 0 -3.0 1e-06 
3.0 3.087 0 -3.0 1e-06 
0.05 3.088 0 -3.0 1e-06 
3.0 3.088 0 -3.0 1e-06 
0.05 3.089 0 -3.0 1e-06 
3.0 3.089 0 -3.0 1e-06 
0.05 3.09 0 -3.0 1e-06 
3.0 3.09 0 -3.0 1e-06 
0.05 3.091 0 -3.0 1e-06 
3.0 3.091 0 -3.0 1e-06 
0.05 3.092 0 -3.0 1e-06 
3.0 3.092 0 -3.0 1e-06 
0.05 3.093 0 -3.0 1e-06 
3.0 3.093 0 -3.0 1e-06 
0.05 3.094 0 -3.0 1e-06 
3.0 3.094 0 -3.0 1e-06 
0.05 3.095 0 -3.0 1e-06 
3.0 3.095 0 -3.0 1e-06 
0.05 3.096 0 -3.0 1e-06 
3.0 3.096 0 -3.0 1e-06 
0.05 3.097 0 -3.0 1e-06 
3.0 3.097 0 -3.0 1e-06 
0.05 3.098 0 -3.0 1e-06 
3.0 3.098 0 -3.0 1e-06 
0.05 3.099 0 -3.0 1e-06 
3.0 3.099 0 -3.0 1e-06 
0.05 3.1 0 -3.0 1e-06 
3.0 3.1 0 -3.0 1e-06 
0.05 3.101 0 -3.0 1e-06 
3.0 3.101 0 -3.0 1e-06 
0.05 3.102 0 -3.0 1e-06 
3.0 3.102 0 -3.0 1e-06 
0.05 3.103 0 -3.0 1e-06 
3.0 3.103 0 -3.0 1e-06 
0.05 3.104 0 -3.0 1e-06 
3.0 3.104 0 -3.0 1e-06 
0.05 3.105 0 -3.0 1e-06 
3.0 3.105 0 -3.0 1e-06 
0.05 3.106 0 -3.0 1e-06 
3.0 3.106 0 -3.0 1e-06 
0.05 3.107 0 -3.0 1e-06 
3.0 3.107 0 -3.0 1e-06 
0.05 3.108 0 -3.0 1e-06 
3.0 3.108 0 -3.0 1e-06 
0.05 3.109 0 -3.0 1e-06 
3.0 3.109 0 -3.0 1e-06 
0.05 3.11 0 -3.0 1e-06 
3.0 3.11 0 -3.0 1e-06 
0.05 3.111 0 -3.0 1e-06 
3.0 3.111 0 -3.0 1e-06 
0.05 3.112 0 -3.0 1e-06 
3.0 3.112 0 -3.0 1e-06 
0.05 3.113 0 -3.0 1e-06 
3.0 3.113 0 -3.0 1e-06 
0.05 3.114 0 -3.0 1e-06 
3.0 3.114 0 -3.0 1e-06 
0.05 3.115 0 -3.0 1e-06 
3.0 3.115 0 -3.0 1e-06 
0.05 3.116 0 -3.0 1e-06 
3.0 3.116 0 -3.0 1e-06 
0.05 3.117 0 -3.0 1e-06 
3.0 3.117 0 -3.0 1e-06 
0.05 3.118 0 -3.0 1e-06 
3.0 3.118 0 -3.0 1e-06 
0.05 3.119 0 -3.0 1e-06 
3.0 3.119 0 -3.0 1e-06 
0.05 3.12 0 -3.0 1e-06 
3.0 3.12 0 -3.0 1e-06 
0.05 3.121 0 -3.0 1e-06 
3.0 3.121 0 -3.0 1e-06 
0.05 3.122 0 -3.0 1e-06 
3.0 3.122 0 -3.0 1e-06 
0.05 3.123 0 -3.0 1e-06 
3.0 3.123 0 -3.0 1e-06 
0.05 3.124 0 -3.0 1e-06 
3.0 3.124 0 -3.0 1e-06 
0.05 3.125 0 -3.0 1e-06 
3.0 3.125 0 -3.0 1e-06 
0.05 3.126 0 -3.0 1e-06 
3.0 3.126 0 -3.0 1e-06 
0.05 3.127 0 -3.0 1e-06 
3.0 3.127 0 -3.0 1e-06 
0.05 3.128 0 -3.0 1e-06 
3.0 3.128 0 -3.0 1e-06 
0.05 3.129 0 -3.0 1e-06 
3.0 3.129 0 -3.0 1e-06 
0.05 3.13 0 -3.0 1e-06 
3.0 3.13 0 -3.0 1e-06 
0.05 3.131 0 -3.0 1e-06 
3.0 3.131 0 -3.0 1e-06 
0.05 3.132 0 -3.0 1e-06 
3.0 3.132 0 -3.0 1e-06 
0.05 3.133 0 -3.0 1e-06 
3.0 3.133 0 -3.0 1e-06 
0.05 3.134 0 -3.0 1e-06 
3.0 3.134 0 -3.0 1e-06 
0.05 3.135 0 -3.0 1e-06 
3.0 3.135 0 -3.0 1e-06 
0.05 3.136 0 -3.0 1e-06 
3.0 3.136 0 -3.0 1e-06 
0.05 3.137 0 -3.0 1e-06 
3.0 3.137 0 -3.0 1e-06 
0.05 3.138 0 -3.0 1e-06 
3.0 3.138 0 -3.0 1e-06 
0.05 3.139 0 -3.0 1e-06 
3.0 3.139 0 -3.0 1e-06 
0.05 3.14 0 -3.0 1e-06 
3.0 3.14 0 -3.0 1e-06 
0.05 3.141 0 -3.0 1e-06 
3.0 3.141 0 -3.0 1e-06 
0.05 3.142 0 -3.0 1e-06 
3.0 3.142 0 -3.0 1e-06 
0.05 3.143 0 -3.0 1e-06 
3.0 3.143 0 -3.0 1e-06 
0.05 3.144 0 -3.0 1e-06 
3.0 3.144 0 -3.0 1e-06 
0.05 3.145 0 -3.0 1e-06 
3.0 3.145 0 -3.0 1e-06 
0.05 3.146 0 -3.0 1e-06 
3.0 3.146 0 -3.0 1e-06 
0.05 3.147 0 -3.0 1e-06 
3.0 3.147 0 -3.0 1e-06 
0.05 3.148 0 -3.0 1e-06 
3.0 3.148 0 -3.0 1e-06 
0.05 3.149 0 -3.0 1e-06 
3.0 3.149 0 -3.0 1e-06 
0.05 3.15 0 -3.0 1e-06 
3.0 3.15 0 -3.0 1e-06 
0.05 3.151 0 -3.0 1e-06 
3.0 3.151 0 -3.0 1e-06 
0.05 3.152 0 -3.0 1e-06 
3.0 3.152 0 -3.0 1e-06 
0.05 3.153 0 -3.0 1e-06 
3.0 3.153 0 -3.0 1e-06 
0.05 3.154 0 -3.0 1e-06 
3.0 3.154 0 -3.0 1e-06 
0.05 3.155 0 -3.0 1e-06 
3.0 3.155 0 -3.0 1e-06 
0.05 3.156 0 -3.0 1e-06 
3.0 3.156 0 -3.0 1e-06 
0.05 3.157 0 -3.0 1e-06 
3.0 3.157 0 -3.0 1e-06 
0.05 3.158 0 -3.0 1e-06 
3.0 3.158 0 -3.0 1e-06 
0.05 3.159 0 -3.0 1e-06 
3.0 3.159 0 -3.0 1e-06 
0.05 3.16 0 -3.0 1e-06 
3.0 3.16 0 -3.0 1e-06 
0.05 3.161 0 -3.0 1e-06 
3.0 3.161 0 -3.0 1e-06 
0.05 3.162 0 -3.0 1e-06 
3.0 3.162 0 -3.0 1e-06 
0.05 3.163 0 -3.0 1e-06 
3.0 3.163 0 -3.0 1e-06 
0.05 3.164 0 -3.0 1e-06 
3.0 3.164 0 -3.0 1e-06 
0.05 3.165 0 -3.0 1e-06 
3.0 3.165 0 -3.0 1e-06 
0.05 3.166 0 -3.0 1e-06 
3.0 3.166 0 -3.0 1e-06 
0.05 3.167 0 -3.0 1e-06 
3.0 3.167 0 -3.0 1e-06 
0.05 3.168 0 -3.0 1e-06 
3.0 3.168 0 -3.0 1e-06 
0.05 3.169 0 -3.0 1e-06 
3.0 3.169 0 -3.0 1e-06 
0.05 3.17 0 -3.0 1e-06 
3.0 3.17 0 -3.0 1e-06 
0.05 3.171 0 -3.0 1e-06 
3.0 3.171 0 -3.0 1e-06 
0.05 3.172 0 -3.0 1e-06 
3.0 3.172 0 -3.0 1e-06 
0.05 3.173 0 -3.0 1e-06 
3.0 3.173 0 -3.0 1e-06 
0.05 3.174 0 -3.0 1e-06 
3.0 3.174 0 -3.0 1e-06 
0.05 3.175 0 -3.0 1e-06 
3.0 3.175 0 -3.0 1e-06 
0.05 3.176 0 -3.0 1e-06 
3.0 3.176 0 -3.0 1e-06 
0.05 3.177 0 -3.0 1e-06 
3.0 3.177 0 -3.0 1e-06 
0.05 3.178 0 -3.0 1e-06 
3.0 3.178 0 -3.0 1e-06 
0.05 3.179 0 -3.0 1e-06 
3.0 3.179 0 -3.0 1e-06 
0.05 3.18 0 -3.0 1e-06 
3.0 3.18 0 -3.0 1e-06 
0.05 3.181 0 -3.0 1e-06 
3.0 3.181 0 -3.0 1e-06 
0.05 3.182 0 -3.0 1e-06 
3.0 3.182 0 -3.0 1e-06 
0.05 3.183 0 -3.0 1e-06 
3.0 3.183 0 -3.0 1e-06 
0.05 3.184 0 -3.0 1e-06 
3.0 3.184 0 -3.0 1e-06 
0.05 3.185 0 -3.0 1e-06 
3.0 3.185 0 -3.0 1e-06 
0.05 3.186 0 -3.0 1e-06 
3.0 3.186 0 -3.0 1e-06 
0.05 3.187 0 -3.0 1e-06 
3.0 3.187 0 -3.0 1e-06 
0.05 3.188 0 -3.0 1e-06 
3.0 3.188 0 -3.0 1e-06 
0.05 3.189 0 -3.0 1e-06 
3.0 3.189 0 -3.0 1e-06 
0.05 3.19 0 -3.0 1e-06 
3.0 3.19 0 -3.0 1e-06 
0.05 3.191 0 -3.0 1e-06 
3.0 3.191 0 -3.0 1e-06 
0.05 3.192 0 -3.0 1e-06 
3.0 3.192 0 -3.0 1e-06 
0.05 3.193 0 -3.0 1e-06 
3.0 3.193 0 -3.0 1e-06 
0.05 3.194 0 -3.0 1e-06 
3.0 3.194 0 -3.0 1e-06 
0.05 3.195 0 -3.0 1e-06 
3.0 3.195 0 -3.0 1e-06 
0.05 3.196 0 -3.0 1e-06 
3.0 3.196 0 -3.0 1e-06 
0.05 3.197 0 -3.0 1e-06 
3.0 3.197 0 -3.0 1e-06 
0.05 3.198 0 -3.0 1e-06 
3.0 3.198 0 -3.0 1e-06 
0.05 3.199 0 -3.0 1e-06 
3.0 3.199 0 -3.0 1e-06 
0.05 3.2 0 -3.0 1e-06 
3.0 3.2 0 -3.0 1e-06 
0.05 3.201 0 -3.0 1e-06 
3.0 3.201 0 -3.0 1e-06 
0.05 3.202 0 -3.0 1e-06 
3.0 3.202 0 -3.0 1e-06 
0.05 3.203 0 -3.0 1e-06 
3.0 3.203 0 -3.0 1e-06 
0.05 3.204 0 -3.0 1e-06 
3.0 3.204 0 -3.0 1e-06 
0.05 3.205 0 -3.0 1e-06 
3.0 3.205 0 -3.0 1e-06 
0.05 3.206 0 -3.0 1e-06 
3.0 3.206 0 -3.0 1e-06 
0.05 3.207 0 -3.0 1e-06 
3.0 3.207 0 -3.0 1e-06 
0.05 3.208 0 -3.0 1e-06 
3.0 3.208 0 -3.0 1e-06 
0.05 3.209 0 -3.0 1e-06 
3.0 3.209 0 -3.0 1e-06 
0.05 3.21 0 -3.0 1e-06 
3.0 3.21 0 -3.0 1e-06 
0.05 3.211 0 -3.0 1e-06 
3.0 3.211 0 -3.0 1e-06 
0.05 3.212 0 -3.0 1e-06 
3.0 3.212 0 -3.0 1e-06 
0.05 3.213 0 -3.0 1e-06 
3.0 3.213 0 -3.0 1e-06 
0.05 3.214 0 -3.0 1e-06 
3.0 3.214 0 -3.0 1e-06 
0.05 3.215 0 -3.0 1e-06 
3.0 3.215 0 -3.0 1e-06 
0.05 3.216 0 -3.0 1e-06 
3.0 3.216 0 -3.0 1e-06 
0.05 3.217 0 -3.0 1e-06 
3.0 3.217 0 -3.0 1e-06 
0.05 3.218 0 -3.0 1e-06 
3.0 3.218 0 -3.0 1e-06 
0.05 3.219 0 -3.0 1e-06 
3.0 3.219 0 -3.0 1e-06 
0.05 3.22 0 -3.0 1e-06 
3.0 3.22 0 -3.0 1e-06 
0.05 3.221 0 -3.0 1e-06 
3.0 3.221 0 -3.0 1e-06 
0.05 3.222 0 -3.0 1e-06 
3.0 3.222 0 -3.0 1e-06 
0.05 3.223 0 -3.0 1e-06 
3.0 3.223 0 -3.0 1e-06 
0.05 3.224 0 -3.0 1e-06 
3.0 3.224 0 -3.0 1e-06 
0.05 3.225 0 -3.0 1e-06 
3.0 3.225 0 -3.0 1e-06 
0.05 3.226 0 -3.0 1e-06 
3.0 3.226 0 -3.0 1e-06 
0.05 3.227 0 -3.0 1e-06 
3.0 3.227 0 -3.0 1e-06 
0.05 3.228 0 -3.0 1e-06 
3.0 3.228 0 -3.0 1e-06 
0.05 3.229 0 -3.0 1e-06 
3.0 3.229 0 -3.0 1e-06 
0.05 3.23 0 -3.0 1e-06 
3.0 3.23 0 -3.0 1e-06 
0.05 3.231 0 -3.0 1e-06 
3.0 3.231 0 -3.0 1e-06 
0.05 3.232 0 -3.0 1e-06 
3.0 3.232 0 -3.0 1e-06 
0.05 3.233 0 -3.0 1e-06 
3.0 3.233 0 -3.0 1e-06 
0.05 3.234 0 -3.0 1e-06 
3.0 3.234 0 -3.0 1e-06 
0.05 3.235 0 -3.0 1e-06 
3.0 3.235 0 -3.0 1e-06 
0.05 3.236 0 -3.0 1e-06 
3.0 3.236 0 -3.0 1e-06 
0.05 3.237 0 -3.0 1e-06 
3.0 3.237 0 -3.0 1e-06 
0.05 3.238 0 -3.0 1e-06 
3.0 3.238 0 -3.0 1e-06 
0.05 3.239 0 -3.0 1e-06 
3.0 3.239 0 -3.0 1e-06 
0.05 3.24 0 -3.0 1e-06 
3.0 3.24 0 -3.0 1e-06 
0.05 3.241 0 -3.0 1e-06 
3.0 3.241 0 -3.0 1e-06 
0.05 3.242 0 -3.0 1e-06 
3.0 3.242 0 -3.0 1e-06 
0.05 3.243 0 -3.0 1e-06 
3.0 3.243 0 -3.0 1e-06 
0.05 3.244 0 -3.0 1e-06 
3.0 3.244 0 -3.0 1e-06 
0.05 3.245 0 -3.0 1e-06 
3.0 3.245 0 -3.0 1e-06 
0.05 3.246 0 -3.0 1e-06 
3.0 3.246 0 -3.0 1e-06 
0.05 3.247 0 -3.0 1e-06 
3.0 3.247 0 -3.0 1e-06 
0.05 3.248 0 -3.0 1e-06 
3.0 3.248 0 -3.0 1e-06 
0.05 3.249 0 -3.0 1e-06 
3.0 3.249 0 -3.0 1e-06 
0.05 3.25 0 -3.0 1e-06 
3.0 3.25 0 -3.0 1e-06 
0.05 3.251 0 -3.0 1e-06 
3.0 3.251 0 -3.0 1e-06 
0.05 3.252 0 -3.0 1e-06 
3.0 3.252 0 -3.0 1e-06 
0.05 3.253 0 -3.0 1e-06 
3.0 3.253 0 -3.0 1e-06 
0.05 3.254 0 -3.0 1e-06 
3.0 3.254 0 -3.0 1e-06 
0.05 3.255 0 -3.0 1e-06 
3.0 3.255 0 -3.0 1e-06 
0.05 3.256 0 -3.0 1e-06 
3.0 3.256 0 -3.0 1e-06 
0.05 3.257 0 -3.0 1e-06 
3.0 3.257 0 -3.0 1e-06 
0.05 3.258 0 -3.0 1e-06 
3.0 3.258 0 -3.0 1e-06 
0.05 3.259 0 -3.0 1e-06 
3.0 3.259 0 -3.0 1e-06 
0.05 3.26 0 -3.0 1e-06 
3.0 3.26 0 -3.0 1e-06 
0.05 3.261 0 -3.0 1e-06 
3.0 3.261 0 -3.0 1e-06 
0.05 3.262 0 -3.0 1e-06 
3.0 3.262 0 -3.0 1e-06 
0.05 3.263 0 -3.0 1e-06 
3.0 3.263 0 -3.0 1e-06 
0.05 3.264 0 -3.0 1e-06 
3.0 3.264 0 -3.0 1e-06 
0.05 3.265 0 -3.0 1e-06 
3.0 3.265 0 -3.0 1e-06 
0.05 3.266 0 -3.0 1e-06 
3.0 3.266 0 -3.0 1e-06 
0.05 3.267 0 -3.0 1e-06 
3.0 3.267 0 -3.0 1e-06 
0.05 3.268 0 -3.0 1e-06 
3.0 3.268 0 -3.0 1e-06 
0.05 3.269 0 -3.0 1e-06 
3.0 3.269 0 -3.0 1e-06 
0.05 3.27 0 -3.0 1e-06 
3.0 3.27 0 -3.0 1e-06 
0.05 3.271 0 -3.0 1e-06 
3.0 3.271 0 -3.0 1e-06 
0.05 3.272 0 -3.0 1e-06 
3.0 3.272 0 -3.0 1e-06 
0.05 3.273 0 -3.0 1e-06 
3.0 3.273 0 -3.0 1e-06 
0.05 3.274 0 -3.0 1e-06 
3.0 3.274 0 -3.0 1e-06 
0.05 3.275 0 -3.0 1e-06 
3.0 3.275 0 -3.0 1e-06 
0.05 3.276 0 -3.0 1e-06 
3.0 3.276 0 -3.0 1e-06 
0.05 3.277 0 -3.0 1e-06 
3.0 3.277 0 -3.0 1e-06 
0.05 3.278 0 -3.0 1e-06 
3.0 3.278 0 -3.0 1e-06 
0.05 3.279 0 -3.0 1e-06 
3.0 3.279 0 -3.0 1e-06 
0.05 3.28 0 -3.0 1e-06 
3.0 3.28 0 -3.0 1e-06 
0.05 3.281 0 -3.0 1e-06 
3.0 3.281 0 -3.0 1e-06 
0.05 3.282 0 -3.0 1e-06 
3.0 3.282 0 -3.0 1e-06 
0.05 3.283 0 -3.0 1e-06 
3.0 3.283 0 -3.0 1e-06 
0.05 3.284 0 -3.0 1e-06 
3.0 3.284 0 -3.0 1e-06 
0.05 3.285 0 -3.0 1e-06 
3.0 3.285 0 -3.0 1e-06 
0.05 3.286 0 -3.0 1e-06 
3.0 3.286 0 -3.0 1e-06 
0.05 3.287 0 -3.0 1e-06 
3.0 3.287 0 -3.0 1e-06 
0.05 3.288 0 -3.0 1e-06 
3.0 3.288 0 -3.0 1e-06 
0.05 3.289 0 -3.0 1e-06 
3.0 3.289 0 -3.0 1e-06 
0.05 3.29 0 -3.0 1e-06 
3.0 3.29 0 -3.0 1e-06 
0.05 3.291 0 -3.0 1e-06 
3.0 3.291 0 -3.0 1e-06 
0.05 3.292 0 -3.0 1e-06 
3.0 3.292 0 -3.0 1e-06 
0.05 3.293 0 -3.0 1e-06 
3.0 3.293 0 -3.0 1e-06 
0.05 3.294 0 -3.0 1e-06 
3.0 3.294 0 -3.0 1e-06 
0.05 3.295 0 -3.0 1e-06 
3.0 3.295 0 -3.0 1e-06 
0.05 3.296 0 -3.0 1e-06 
3.0 3.296 0 -3.0 1e-06 
0.05 3.297 0 -3.0 1e-06 
3.0 3.297 0 -3.0 1e-06 
0.05 3.298 0 -3.0 1e-06 
3.0 3.298 0 -3.0 1e-06 
0.05 3.299 0 -3.0 1e-06 
3.0 3.299 0 -3.0 1e-06 
0.05 3.3 0 -3.0 1e-06 
3.0 3.3 0 -3.0 1e-06 
0.05 3.301 0 -3.0 1e-06 
3.0 3.301 0 -3.0 1e-06 
0.05 3.302 0 -3.0 1e-06 
3.0 3.302 0 -3.0 1e-06 
0.05 3.303 0 -3.0 1e-06 
3.0 3.303 0 -3.0 1e-06 
0.05 3.304 0 -3.0 1e-06 
3.0 3.304 0 -3.0 1e-06 
0.05 3.305 0 -3.0 1e-06 
3.0 3.305 0 -3.0 1e-06 
0.05 3.306 0 -3.0 1e-06 
3.0 3.306 0 -3.0 1e-06 
0.05 3.307 0 -3.0 1e-06 
3.0 3.307 0 -3.0 1e-06 
0.05 3.308 0 -3.0 1e-06 
3.0 3.308 0 -3.0 1e-06 
0.05 3.309 0 -3.0 1e-06 
3.0 3.309 0 -3.0 1e-06 
0.05 3.31 0 -3.0 1e-06 
3.0 3.31 0 -3.0 1e-06 
0.05 3.311 0 -3.0 1e-06 
3.0 3.311 0 -3.0 1e-06 
0.05 3.312 0 -3.0 1e-06 
3.0 3.312 0 -3.0 1e-06 
0.05 3.313 0 -3.0 1e-06 
3.0 3.313 0 -3.0 1e-06 
0.05 3.314 0 -3.0 1e-06 
3.0 3.314 0 -3.0 1e-06 
0.05 3.315 0 -3.0 1e-06 
3.0 3.315 0 -3.0 1e-06 
0.05 3.316 0 -3.0 1e-06 
3.0 3.316 0 -3.0 1e-06 
0.05 3.317 0 -3.0 1e-06 
3.0 3.317 0 -3.0 1e-06 
0.05 3.318 0 -3.0 1e-06 
3.0 3.318 0 -3.0 1e-06 
0.05 3.319 0 -3.0 1e-06 
3.0 3.319 0 -3.0 1e-06 
0.05 3.32 0 -3.0 1e-06 
3.0 3.32 0 -3.0 1e-06 
0.05 3.321 0 -3.0 1e-06 
3.0 3.321 0 -3.0 1e-06 
0.05 3.322 0 -3.0 1e-06 
3.0 3.322 0 -3.0 1e-06 
0.05 3.323 0 -3.0 1e-06 
3.0 3.323 0 -3.0 1e-06 
0.05 3.324 0 -3.0 1e-06 
3.0 3.324 0 -3.0 1e-06 
0.05 3.325 0 -3.0 1e-06 
3.0 3.325 0 -3.0 1e-06 
0.05 3.326 0 -3.0 1e-06 
3.0 3.326 0 -3.0 1e-06 
0.05 3.327 0 -3.0 1e-06 
3.0 3.327 0 -3.0 1e-06 
0.05 3.328 0 -3.0 1e-06 
3.0 3.328 0 -3.0 1e-06 
0.05 3.329 0 -3.0 1e-06 
3.0 3.329 0 -3.0 1e-06 
0.05 3.33 0 -3.0 1e-06 
3.0 3.33 0 -3.0 1e-06 
0.05 3.331 0 -3.0 1e-06 
3.0 3.331 0 -3.0 1e-06 
0.05 3.332 0 -3.0 1e-06 
3.0 3.332 0 -3.0 1e-06 
0.05 3.333 0 -3.0 1e-06 
3.0 3.333 0 -3.0 1e-06 
0.05 3.334 0 -3.0 1e-06 
3.0 3.334 0 -3.0 1e-06 
0.05 3.335 0 -3.0 1e-06 
3.0 3.335 0 -3.0 1e-06 
0.05 3.336 0 -3.0 1e-06 
3.0 3.336 0 -3.0 1e-06 
0.05 3.337 0 -3.0 1e-06 
3.0 3.337 0 -3.0 1e-06 
0.05 3.338 0 -3.0 1e-06 
3.0 3.338 0 -3.0 1e-06 
0.05 3.339 0 -3.0 1e-06 
3.0 3.339 0 -3.0 1e-06 
0.05 3.34 0 -3.0 1e-06 
3.0 3.34 0 -3.0 1e-06 
0.05 3.341 0 -3.0 1e-06 
3.0 3.341 0 -3.0 1e-06 
0.05 3.342 0 -3.0 1e-06 
3.0 3.342 0 -3.0 1e-06 
0.05 3.343 0 -3.0 1e-06 
3.0 3.343 0 -3.0 1e-06 
0.05 3.344 0 -3.0 1e-06 
3.0 3.344 0 -3.0 1e-06 
0.05 3.345 0 -3.0 1e-06 
3.0 3.345 0 -3.0 1e-06 
0.05 3.346 0 -3.0 1e-06 
3.0 3.346 0 -3.0 1e-06 
0.05 3.347 0 -3.0 1e-06 
3.0 3.347 0 -3.0 1e-06 
0.05 3.348 0 -3.0 1e-06 
3.0 3.348 0 -3.0 1e-06 
0.05 3.349 0 -3.0 1e-06 
3.0 3.349 0 -3.0 1e-06 
0.05 3.35 0 -3.0 1e-06 
3.0 3.35 0 -3.0 1e-06 
0.05 3.351 0 -3.0 1e-06 
3.0 3.351 0 -3.0 1e-06 
0.05 3.352 0 -3.0 1e-06 
3.0 3.352 0 -3.0 1e-06 
0.05 3.353 0 -3.0 1e-06 
3.0 3.353 0 -3.0 1e-06 
0.05 3.354 0 -3.0 1e-06 
3.0 3.354 0 -3.0 1e-06 
0.05 3.355 0 -3.0 1e-06 
3.0 3.355 0 -3.0 1e-06 
0.05 3.356 0 -3.0 1e-06 
3.0 3.356 0 -3.0 1e-06 
0.05 3.357 0 -3.0 1e-06 
3.0 3.357 0 -3.0 1e-06 
0.05 3.358 0 -3.0 1e-06 
3.0 3.358 0 -3.0 1e-06 
0.05 3.359 0 -3.0 1e-06 
3.0 3.359 0 -3.0 1e-06 
0.05 3.36 0 -3.0 1e-06 
3.0 3.36 0 -3.0 1e-06 
0.05 3.361 0 -3.0 1e-06 
3.0 3.361 0 -3.0 1e-06 
0.05 3.362 0 -3.0 1e-06 
3.0 3.362 0 -3.0 1e-06 
0.05 3.363 0 -3.0 1e-06 
3.0 3.363 0 -3.0 1e-06 
0.05 3.364 0 -3.0 1e-06 
3.0 3.364 0 -3.0 1e-06 
0.05 3.365 0 -3.0 1e-06 
3.0 3.365 0 -3.0 1e-06 
0.05 3.366 0 -3.0 1e-06 
3.0 3.366 0 -3.0 1e-06 
0.05 3.367 0 -3.0 1e-06 
3.0 3.367 0 -3.0 1e-06 
0.05 3.368 0 -3.0 1e-06 
3.0 3.368 0 -3.0 1e-06 
0.05 3.369 0 -3.0 1e-06 
3.0 3.369 0 -3.0 1e-06 
0.05 3.37 0 -3.0 1e-06 
3.0 3.37 0 -3.0 1e-06 
0.05 3.371 0 -3.0 1e-06 
3.0 3.371 0 -3.0 1e-06 
0.05 3.372 0 -3.0 1e-06 
3.0 3.372 0 -3.0 1e-06 
0.05 3.373 0 -3.0 1e-06 
3.0 3.373 0 -3.0 1e-06 
0.05 3.374 0 -3.0 1e-06 
3.0 3.374 0 -3.0 1e-06 
0.05 3.375 0 -3.0 1e-06 
3.0 3.375 0 -3.0 1e-06 
0.05 3.376 0 -3.0 1e-06 
3.0 3.376 0 -3.0 1e-06 
0.05 3.377 0 -3.0 1e-06 
3.0 3.377 0 -3.0 1e-06 
0.05 3.378 0 -3.0 1e-06 
3.0 3.378 0 -3.0 1e-06 
0.05 3.379 0 -3.0 1e-06 
3.0 3.379 0 -3.0 1e-06 
0.05 3.38 0 -3.0 1e-06 
3.0 3.38 0 -3.0 1e-06 
0.05 3.381 0 -3.0 1e-06 
3.0 3.381 0 -3.0 1e-06 
0.05 3.382 0 -3.0 1e-06 
3.0 3.382 0 -3.0 1e-06 
0.05 3.383 0 -3.0 1e-06 
3.0 3.383 0 -3.0 1e-06 
0.05 3.384 0 -3.0 1e-06 
3.0 3.384 0 -3.0 1e-06 
0.05 3.385 0 -3.0 1e-06 
3.0 3.385 0 -3.0 1e-06 
0.05 3.386 0 -3.0 1e-06 
3.0 3.386 0 -3.0 1e-06 
0.05 3.387 0 -3.0 1e-06 
3.0 3.387 0 -3.0 1e-06 
0.05 3.388 0 -3.0 1e-06 
3.0 3.388 0 -3.0 1e-06 
0.05 3.389 0 -3.0 1e-06 
3.0 3.389 0 -3.0 1e-06 
0.05 3.39 0 -3.0 1e-06 
3.0 3.39 0 -3.0 1e-06 
0.05 3.391 0 -3.0 1e-06 
3.0 3.391 0 -3.0 1e-06 
0.05 3.392 0 -3.0 1e-06 
3.0 3.392 0 -3.0 1e-06 
0.05 3.393 0 -3.0 1e-06 
3.0 3.393 0 -3.0 1e-06 
0.05 3.394 0 -3.0 1e-06 
3.0 3.394 0 -3.0 1e-06 
0.05 3.395 0 -3.0 1e-06 
3.0 3.395 0 -3.0 1e-06 
0.05 3.396 0 -3.0 1e-06 
3.0 3.396 0 -3.0 1e-06 
0.05 3.397 0 -3.0 1e-06 
3.0 3.397 0 -3.0 1e-06 
0.05 3.398 0 -3.0 1e-06 
3.0 3.398 0 -3.0 1e-06 
0.05 3.399 0 -3.0 1e-06 
3.0 3.399 0 -3.0 1e-06 
0.05 3.4 0 -3.0 1e-06 
3.0 3.4 0 -3.0 1e-06 
0.05 3.401 0 -3.0 1e-06 
3.0 3.401 0 -3.0 1e-06 
0.05 3.402 0 -3.0 1e-06 
3.0 3.402 0 -3.0 1e-06 
0.05 3.403 0 -3.0 1e-06 
3.0 3.403 0 -3.0 1e-06 
0.05 3.404 0 -3.0 1e-06 
3.0 3.404 0 -3.0 1e-06 
0.05 3.405 0 -3.0 1e-06 
3.0 3.405 0 -3.0 1e-06 
0.05 3.406 0 -3.0 1e-06 
3.0 3.406 0 -3.0 1e-06 
0.05 3.407 0 -3.0 1e-06 
3.0 3.407 0 -3.0 1e-06 
0.05 3.408 0 -3.0 1e-06 
3.0 3.408 0 -3.0 1e-06 
0.05 3.409 0 -3.0 1e-06 
3.0 3.409 0 -3.0 1e-06 
0.05 3.41 0 -3.0 1e-06 
3.0 3.41 0 -3.0 1e-06 
0.05 3.411 0 -3.0 1e-06 
3.0 3.411 0 -3.0 1e-06 
0.05 3.412 0 -3.0 1e-06 
3.0 3.412 0 -3.0 1e-06 
0.05 3.413 0 -3.0 1e-06 
3.0 3.413 0 -3.0 1e-06 
0.05 3.414 0 -3.0 1e-06 
3.0 3.414 0 -3.0 1e-06 
0.05 3.415 0 -3.0 1e-06 
3.0 3.415 0 -3.0 1e-06 
0.05 3.416 0 -3.0 1e-06 
3.0 3.416 0 -3.0 1e-06 
0.05 3.417 0 -3.0 1e-06 
3.0 3.417 0 -3.0 1e-06 
0.05 3.418 0 -3.0 1e-06 
3.0 3.418 0 -3.0 1e-06 
0.05 3.419 0 -3.0 1e-06 
3.0 3.419 0 -3.0 1e-06 
0.05 3.42 0 -3.0 1e-06 
3.0 3.42 0 -3.0 1e-06 
0.05 3.421 0 -3.0 1e-06 
3.0 3.421 0 -3.0 1e-06 
0.05 3.422 0 -3.0 1e-06 
3.0 3.422 0 -3.0 1e-06 
0.05 3.423 0 -3.0 1e-06 
3.0 3.423 0 -3.0 1e-06 
0.05 3.424 0 -3.0 1e-06 
3.0 3.424 0 -3.0 1e-06 
0.05 3.425 0 -3.0 1e-06 
3.0 3.425 0 -3.0 1e-06 
0.05 3.426 0 -3.0 1e-06 
3.0 3.426 0 -3.0 1e-06 
0.05 3.427 0 -3.0 1e-06 
3.0 3.427 0 -3.0 1e-06 
0.05 3.428 0 -3.0 1e-06 
3.0 3.428 0 -3.0 1e-06 
0.05 3.429 0 -3.0 1e-06 
3.0 3.429 0 -3.0 1e-06 
0.05 3.43 0 -3.0 1e-06 
3.0 3.43 0 -3.0 1e-06 
0.05 3.431 0 -3.0 1e-06 
3.0 3.431 0 -3.0 1e-06 
0.05 3.432 0 -3.0 1e-06 
3.0 3.432 0 -3.0 1e-06 
0.05 3.433 0 -3.0 1e-06 
3.0 3.433 0 -3.0 1e-06 
0.05 3.434 0 -3.0 1e-06 
3.0 3.434 0 -3.0 1e-06 
0.05 3.435 0 -3.0 1e-06 
3.0 3.435 0 -3.0 1e-06 
0.05 3.436 0 -3.0 1e-06 
3.0 3.436 0 -3.0 1e-06 
0.05 3.437 0 -3.0 1e-06 
3.0 3.437 0 -3.0 1e-06 
0.05 3.438 0 -3.0 1e-06 
3.0 3.438 0 -3.0 1e-06 
0.05 3.439 0 -3.0 1e-06 
3.0 3.439 0 -3.0 1e-06 
0.05 3.44 0 -3.0 1e-06 
3.0 3.44 0 -3.0 1e-06 
0.05 3.441 0 -3.0 1e-06 
3.0 3.441 0 -3.0 1e-06 
0.05 3.442 0 -3.0 1e-06 
3.0 3.442 0 -3.0 1e-06 
0.05 3.443 0 -3.0 1e-06 
3.0 3.443 0 -3.0 1e-06 
0.05 3.444 0 -3.0 1e-06 
3.0 3.444 0 -3.0 1e-06 
0.05 3.445 0 -3.0 1e-06 
3.0 3.445 0 -3.0 1e-06 
0.05 3.446 0 -3.0 1e-06 
3.0 3.446 0 -3.0 1e-06 
0.05 3.447 0 -3.0 1e-06 
3.0 3.447 0 -3.0 1e-06 
0.05 3.448 0 -3.0 1e-06 
3.0 3.448 0 -3.0 1e-06 
0.05 3.449 0 -3.0 1e-06 
3.0 3.449 0 -3.0 1e-06 
0.05 3.45 0 -3.0 1e-06 
3.0 3.45 0 -3.0 1e-06 
0.05 3.451 0 -3.0 1e-06 
3.0 3.451 0 -3.0 1e-06 
0.05 3.452 0 -3.0 1e-06 
3.0 3.452 0 -3.0 1e-06 
0.05 3.453 0 -3.0 1e-06 
3.0 3.453 0 -3.0 1e-06 
0.05 3.454 0 -3.0 1e-06 
3.0 3.454 0 -3.0 1e-06 
0.05 3.455 0 -3.0 1e-06 
3.0 3.455 0 -3.0 1e-06 
0.05 3.456 0 -3.0 1e-06 
3.0 3.456 0 -3.0 1e-06 
0.05 3.457 0 -3.0 1e-06 
3.0 3.457 0 -3.0 1e-06 
0.05 3.458 0 -3.0 1e-06 
3.0 3.458 0 -3.0 1e-06 
0.05 3.459 0 -3.0 1e-06 
3.0 3.459 0 -3.0 1e-06 
0.05 3.46 0 -3.0 1e-06 
3.0 3.46 0 -3.0 1e-06 
0.05 3.461 0 -3.0 1e-06 
3.0 3.461 0 -3.0 1e-06 
0.05 3.462 0 -3.0 1e-06 
3.0 3.462 0 -3.0 1e-06 
0.05 3.463 0 -3.0 1e-06 
3.0 3.463 0 -3.0 1e-06 
0.05 3.464 0 -3.0 1e-06 
3.0 3.464 0 -3.0 1e-06 
0.05 3.465 0 -3.0 1e-06 
3.0 3.465 0 -3.0 1e-06 
0.05 3.466 0 -3.0 1e-06 
3.0 3.466 0 -3.0 1e-06 
0.05 3.467 0 -3.0 1e-06 
3.0 3.467 0 -3.0 1e-06 
0.05 3.468 0 -3.0 1e-06 
3.0 3.468 0 -3.0 1e-06 
0.05 3.469 0 -3.0 1e-06 
3.0 3.469 0 -3.0 1e-06 
0.05 3.47 0 -3.0 1e-06 
3.0 3.47 0 -3.0 1e-06 
0.05 3.471 0 -3.0 1e-06 
3.0 3.471 0 -3.0 1e-06 
0.05 3.472 0 -3.0 1e-06 
3.0 3.472 0 -3.0 1e-06 
0.05 3.473 0 -3.0 1e-06 
3.0 3.473 0 -3.0 1e-06 
0.05 3.474 0 -3.0 1e-06 
3.0 3.474 0 -3.0 1e-06 
0.05 3.475 0 -3.0 1e-06 
3.0 3.475 0 -3.0 1e-06 
0.05 3.476 0 -3.0 1e-06 
3.0 3.476 0 -3.0 1e-06 
0.05 3.477 0 -3.0 1e-06 
3.0 3.477 0 -3.0 1e-06 
0.05 3.478 0 -3.0 1e-06 
3.0 3.478 0 -3.0 1e-06 
0.05 3.479 0 -3.0 1e-06 
3.0 3.479 0 -3.0 1e-06 
0.05 3.48 0 -3.0 1e-06 
3.0 3.48 0 -3.0 1e-06 
0.05 3.481 0 -3.0 1e-06 
3.0 3.481 0 -3.0 1e-06 
0.05 3.482 0 -3.0 1e-06 
3.0 3.482 0 -3.0 1e-06 
0.05 3.483 0 -3.0 1e-06 
3.0 3.483 0 -3.0 1e-06 
0.05 3.484 0 -3.0 1e-06 
3.0 3.484 0 -3.0 1e-06 
0.05 3.485 0 -3.0 1e-06 
3.0 3.485 0 -3.0 1e-06 
0.05 3.486 0 -3.0 1e-06 
3.0 3.486 0 -3.0 1e-06 
0.05 3.487 0 -3.0 1e-06 
3.0 3.487 0 -3.0 1e-06 
0.05 3.488 0 -3.0 1e-06 
3.0 3.488 0 -3.0 1e-06 
0.05 3.489 0 -3.0 1e-06 
3.0 3.489 0 -3.0 1e-06 
0.05 3.49 0 -3.0 1e-06 
3.0 3.49 0 -3.0 1e-06 
0.05 3.491 0 -3.0 1e-06 
3.0 3.491 0 -3.0 1e-06 
0.05 3.492 0 -3.0 1e-06 
3.0 3.492 0 -3.0 1e-06 
0.05 3.493 0 -3.0 1e-06 
3.0 3.493 0 -3.0 1e-06 
0.05 3.494 0 -3.0 1e-06 
3.0 3.494 0 -3.0 1e-06 
0.05 3.495 0 -3.0 1e-06 
3.0 3.495 0 -3.0 1e-06 
0.05 3.496 0 -3.0 1e-06 
3.0 3.496 0 -3.0 1e-06 
0.05 3.497 0 -3.0 1e-06 
3.0 3.497 0 -3.0 1e-06 
0.05 3.498 0 -3.0 1e-06 
3.0 3.498 0 -3.0 1e-06 
0.05 3.499 0 -3.0 1e-06 
3.0 3.499 0 -3.0 1e-06 
0.05 3.5 0 -3.0 1e-06 
3.0 3.5 0 -3.0 1e-06 
0.05 3.501 0 -3.0 1e-06 
3.0 3.501 0 -3.0 1e-06 
0.05 3.502 0 -3.0 1e-06 
3.0 3.502 0 -3.0 1e-06 
0.05 3.503 0 -3.0 1e-06 
3.0 3.503 0 -3.0 1e-06 
0.05 3.504 0 -3.0 1e-06 
3.0 3.504 0 -3.0 1e-06 
0.05 3.505 0 -3.0 1e-06 
3.0 3.505 0 -3.0 1e-06 
0.05 3.506 0 -3.0 1e-06 
3.0 3.506 0 -3.0 1e-06 
0.05 3.507 0 -3.0 1e-06 
3.0 3.507 0 -3.0 1e-06 
0.05 3.508 0 -3.0 1e-06 
3.0 3.508 0 -3.0 1e-06 
0.05 3.509 0 -3.0 1e-06 
3.0 3.509 0 -3.0 1e-06 
0.05 3.51 0 -3.0 1e-06 
3.0 3.51 0 -3.0 1e-06 
0.05 3.511 0 -3.0 1e-06 
3.0 3.511 0 -3.0 1e-06 
0.05 3.512 0 -3.0 1e-06 
3.0 3.512 0 -3.0 1e-06 
0.05 3.513 0 -3.0 1e-06 
3.0 3.513 0 -3.0 1e-06 
0.05 3.514 0 -3.0 1e-06 
3.0 3.514 0 -3.0 1e-06 
0.05 3.515 0 -3.0 1e-06 
3.0 3.515 0 -3.0 1e-06 
0.05 3.516 0 -3.0 1e-06 
3.0 3.516 0 -3.0 1e-06 
0.05 3.517 0 -3.0 1e-06 
3.0 3.517 0 -3.0 1e-06 
0.05 3.518 0 -3.0 1e-06 
3.0 3.518 0 -3.0 1e-06 
0.05 3.519 0 -3.0 1e-06 
3.0 3.519 0 -3.0 1e-06 
0.05 3.52 0 -3.0 1e-06 
3.0 3.52 0 -3.0 1e-06 
0.05 3.521 0 -3.0 1e-06 
3.0 3.521 0 -3.0 1e-06 
0.05 3.522 0 -3.0 1e-06 
3.0 3.522 0 -3.0 1e-06 
0.05 3.523 0 -3.0 1e-06 
3.0 3.523 0 -3.0 1e-06 
0.05 3.524 0 -3.0 1e-06 
3.0 3.524 0 -3.0 1e-06 
0.05 3.525 0 -3.0 1e-06 
3.0 3.525 0 -3.0 1e-06 
0.05 3.526 0 -3.0 1e-06 
3.0 3.526 0 -3.0 1e-06 
0.05 3.527 0 -3.0 1e-06 
3.0 3.527 0 -3.0 1e-06 
0.05 3.528 0 -3.0 1e-06 
3.0 3.528 0 -3.0 1e-06 
0.05 3.529 0 -3.0 1e-06 
3.0 3.529 0 -3.0 1e-06 
0.05 3.53 0 -3.0 1e-06 
3.0 3.53 0 -3.0 1e-06 
0.05 3.531 0 -3.0 1e-06 
3.0 3.531 0 -3.0 1e-06 
0.05 3.532 0 -3.0 1e-06 
3.0 3.532 0 -3.0 1e-06 
0.05 3.533 0 -3.0 1e-06 
3.0 3.533 0 -3.0 1e-06 
0.05 3.534 0 -3.0 1e-06 
3.0 3.534 0 -3.0 1e-06 
0.05 3.535 0 -3.0 1e-06 
3.0 3.535 0 -3.0 1e-06 
0.05 3.536 0 -3.0 1e-06 
3.0 3.536 0 -3.0 1e-06 
0.05 3.537 0 -3.0 1e-06 
3.0 3.537 0 -3.0 1e-06 
0.05 3.538 0 -3.0 1e-06 
3.0 3.538 0 -3.0 1e-06 
0.05 3.539 0 -3.0 1e-06 
3.0 3.539 0 -3.0 1e-06 
0.05 3.54 0 -3.0 1e-06 
3.0 3.54 0 -3.0 1e-06 
0.05 3.541 0 -3.0 1e-06 
3.0 3.541 0 -3.0 1e-06 
0.05 3.542 0 -3.0 1e-06 
3.0 3.542 0 -3.0 1e-06 
0.05 3.543 0 -3.0 1e-06 
3.0 3.543 0 -3.0 1e-06 
0.05 3.544 0 -3.0 1e-06 
3.0 3.544 0 -3.0 1e-06 
0.05 3.545 0 -3.0 1e-06 
3.0 3.545 0 -3.0 1e-06 
0.05 3.546 0 -3.0 1e-06 
3.0 3.546 0 -3.0 1e-06 
0.05 3.547 0 -3.0 1e-06 
3.0 3.547 0 -3.0 1e-06 
0.05 3.548 0 -3.0 1e-06 
3.0 3.548 0 -3.0 1e-06 
0.05 3.549 0 -3.0 1e-06 
3.0 3.549 0 -3.0 1e-06 
0.05 3.55 0 -3.0 1e-06 
3.0 3.55 0 -3.0 1e-06 
0.05 3.551 0 -3.0 1e-06 
3.0 3.551 0 -3.0 1e-06 
0.05 3.552 0 -3.0 1e-06 
3.0 3.552 0 -3.0 1e-06 
0.05 3.553 0 -3.0 1e-06 
3.0 3.553 0 -3.0 1e-06 
0.05 3.554 0 -3.0 1e-06 
3.0 3.554 0 -3.0 1e-06 
0.05 3.555 0 -3.0 1e-06 
3.0 3.555 0 -3.0 1e-06 
0.05 3.556 0 -3.0 1e-06 
3.0 3.556 0 -3.0 1e-06 
0.05 3.557 0 -3.0 1e-06 
3.0 3.557 0 -3.0 1e-06 
0.05 3.558 0 -3.0 1e-06 
3.0 3.558 0 -3.0 1e-06 
0.05 3.559 0 -3.0 1e-06 
3.0 3.559 0 -3.0 1e-06 
0.05 3.56 0 -3.0 1e-06 
3.0 3.56 0 -3.0 1e-06 
0.05 3.561 0 -3.0 1e-06 
3.0 3.561 0 -3.0 1e-06 
0.05 3.562 0 -3.0 1e-06 
3.0 3.562 0 -3.0 1e-06 
0.05 3.563 0 -3.0 1e-06 
3.0 3.563 0 -3.0 1e-06 
0.05 3.564 0 -3.0 1e-06 
3.0 3.564 0 -3.0 1e-06 
0.05 3.565 0 -3.0 1e-06 
3.0 3.565 0 -3.0 1e-06 
0.05 3.566 0 -3.0 1e-06 
3.0 3.566 0 -3.0 1e-06 
0.05 3.567 0 -3.0 1e-06 
3.0 3.567 0 -3.0 1e-06 
0.05 3.568 0 -3.0 1e-06 
3.0 3.568 0 -3.0 1e-06 
0.05 3.569 0 -3.0 1e-06 
3.0 3.569 0 -3.0 1e-06 
0.05 3.57 0 -3.0 1e-06 
3.0 3.57 0 -3.0 1e-06 
0.05 3.571 0 -3.0 1e-06 
3.0 3.571 0 -3.0 1e-06 
0.05 3.572 0 -3.0 1e-06 
3.0 3.572 0 -3.0 1e-06 
0.05 3.573 0 -3.0 1e-06 
3.0 3.573 0 -3.0 1e-06 
0.05 3.574 0 -3.0 1e-06 
3.0 3.574 0 -3.0 1e-06 
0.05 3.575 0 -3.0 1e-06 
3.0 3.575 0 -3.0 1e-06 
0.05 3.576 0 -3.0 1e-06 
3.0 3.576 0 -3.0 1e-06 
0.05 3.577 0 -3.0 1e-06 
3.0 3.577 0 -3.0 1e-06 
0.05 3.578 0 -3.0 1e-06 
3.0 3.578 0 -3.0 1e-06 
0.05 3.579 0 -3.0 1e-06 
3.0 3.579 0 -3.0 1e-06 
0.05 3.58 0 -3.0 1e-06 
3.0 3.58 0 -3.0 1e-06 
0.05 3.581 0 -3.0 1e-06 
3.0 3.581 0 -3.0 1e-06 
0.05 3.582 0 -3.0 1e-06 
3.0 3.582 0 -3.0 1e-06 
0.05 3.583 0 -3.0 1e-06 
3.0 3.583 0 -3.0 1e-06 
0.05 3.584 0 -3.0 1e-06 
3.0 3.584 0 -3.0 1e-06 
0.05 3.585 0 -3.0 1e-06 
3.0 3.585 0 -3.0 1e-06 
0.05 3.586 0 -3.0 1e-06 
3.0 3.586 0 -3.0 1e-06 
0.05 3.587 0 -3.0 1e-06 
3.0 3.587 0 -3.0 1e-06 
0.05 3.588 0 -3.0 1e-06 
3.0 3.588 0 -3.0 1e-06 
0.05 3.589 0 -3.0 1e-06 
3.0 3.589 0 -3.0 1e-06 
0.05 3.59 0 -3.0 1e-06 
3.0 3.59 0 -3.0 1e-06 
0.05 3.591 0 -3.0 1e-06 
3.0 3.591 0 -3.0 1e-06 
0.05 3.592 0 -3.0 1e-06 
3.0 3.592 0 -3.0 1e-06 
0.05 3.593 0 -3.0 1e-06 
3.0 3.593 0 -3.0 1e-06 
0.05 3.594 0 -3.0 1e-06 
3.0 3.594 0 -3.0 1e-06 
0.05 3.595 0 -3.0 1e-06 
3.0 3.595 0 -3.0 1e-06 
0.05 3.596 0 -3.0 1e-06 
3.0 3.596 0 -3.0 1e-06 
0.05 3.597 0 -3.0 1e-06 
3.0 3.597 0 -3.0 1e-06 
0.05 3.598 0 -3.0 1e-06 
3.0 3.598 0 -3.0 1e-06 
0.05 3.599 0 -3.0 1e-06 
3.0 3.599 0 -3.0 1e-06 
0.05 3.6 0 -3.0 1e-06 
3.0 3.6 0 -3.0 1e-06 
0.05 3.601 0 -3.0 1e-06 
3.0 3.601 0 -3.0 1e-06 
0.05 3.602 0 -3.0 1e-06 
3.0 3.602 0 -3.0 1e-06 
0.05 3.603 0 -3.0 1e-06 
3.0 3.603 0 -3.0 1e-06 
0.05 3.604 0 -3.0 1e-06 
3.0 3.604 0 -3.0 1e-06 
0.05 3.605 0 -3.0 1e-06 
3.0 3.605 0 -3.0 1e-06 
0.05 3.606 0 -3.0 1e-06 
3.0 3.606 0 -3.0 1e-06 
0.05 3.607 0 -3.0 1e-06 
3.0 3.607 0 -3.0 1e-06 
0.05 3.608 0 -3.0 1e-06 
3.0 3.608 0 -3.0 1e-06 
0.05 3.609 0 -3.0 1e-06 
3.0 3.609 0 -3.0 1e-06 
0.05 3.61 0 -3.0 1e-06 
3.0 3.61 0 -3.0 1e-06 
0.05 3.611 0 -3.0 1e-06 
3.0 3.611 0 -3.0 1e-06 
0.05 3.612 0 -3.0 1e-06 
3.0 3.612 0 -3.0 1e-06 
0.05 3.613 0 -3.0 1e-06 
3.0 3.613 0 -3.0 1e-06 
0.05 3.614 0 -3.0 1e-06 
3.0 3.614 0 -3.0 1e-06 
0.05 3.615 0 -3.0 1e-06 
3.0 3.615 0 -3.0 1e-06 
0.05 3.616 0 -3.0 1e-06 
3.0 3.616 0 -3.0 1e-06 
0.05 3.617 0 -3.0 1e-06 
3.0 3.617 0 -3.0 1e-06 
0.05 3.618 0 -3.0 1e-06 
3.0 3.618 0 -3.0 1e-06 
0.05 3.619 0 -3.0 1e-06 
3.0 3.619 0 -3.0 1e-06 
0.05 3.62 0 -3.0 1e-06 
3.0 3.62 0 -3.0 1e-06 
0.05 3.621 0 -3.0 1e-06 
3.0 3.621 0 -3.0 1e-06 
0.05 3.622 0 -3.0 1e-06 
3.0 3.622 0 -3.0 1e-06 
0.05 3.623 0 -3.0 1e-06 
3.0 3.623 0 -3.0 1e-06 
0.05 3.624 0 -3.0 1e-06 
3.0 3.624 0 -3.0 1e-06 
0.05 3.625 0 -3.0 1e-06 
3.0 3.625 0 -3.0 1e-06 
0.05 3.626 0 -3.0 1e-06 
3.0 3.626 0 -3.0 1e-06 
0.05 3.627 0 -3.0 1e-06 
3.0 3.627 0 -3.0 1e-06 
0.05 3.628 0 -3.0 1e-06 
3.0 3.628 0 -3.0 1e-06 
0.05 3.629 0 -3.0 1e-06 
3.0 3.629 0 -3.0 1e-06 
0.05 3.63 0 -3.0 1e-06 
3.0 3.63 0 -3.0 1e-06 
0.05 3.631 0 -3.0 1e-06 
3.0 3.631 0 -3.0 1e-06 
0.05 3.632 0 -3.0 1e-06 
3.0 3.632 0 -3.0 1e-06 
0.05 3.633 0 -3.0 1e-06 
3.0 3.633 0 -3.0 1e-06 
0.05 3.634 0 -3.0 1e-06 
3.0 3.634 0 -3.0 1e-06 
0.05 3.635 0 -3.0 1e-06 
3.0 3.635 0 -3.0 1e-06 
0.05 3.636 0 -3.0 1e-06 
3.0 3.636 0 -3.0 1e-06 
0.05 3.637 0 -3.0 1e-06 
3.0 3.637 0 -3.0 1e-06 
0.05 3.638 0 -3.0 1e-06 
3.0 3.638 0 -3.0 1e-06 
0.05 3.639 0 -3.0 1e-06 
3.0 3.639 0 -3.0 1e-06 
0.05 3.64 0 -3.0 1e-06 
3.0 3.64 0 -3.0 1e-06 
0.05 3.641 0 -3.0 1e-06 
3.0 3.641 0 -3.0 1e-06 
0.05 3.642 0 -3.0 1e-06 
3.0 3.642 0 -3.0 1e-06 
0.05 3.643 0 -3.0 1e-06 
3.0 3.643 0 -3.0 1e-06 
0.05 3.644 0 -3.0 1e-06 
3.0 3.644 0 -3.0 1e-06 
0.05 3.645 0 -3.0 1e-06 
3.0 3.645 0 -3.0 1e-06 
0.05 3.646 0 -3.0 1e-06 
3.0 3.646 0 -3.0 1e-06 
0.05 3.647 0 -3.0 1e-06 
3.0 3.647 0 -3.0 1e-06 
0.05 3.648 0 -3.0 1e-06 
3.0 3.648 0 -3.0 1e-06 
0.05 3.649 0 -3.0 1e-06 
3.0 3.649 0 -3.0 1e-06 
0.05 3.65 0 -3.0 1e-06 
3.0 3.65 0 -3.0 1e-06 
0.05 3.651 0 -3.0 1e-06 
3.0 3.651 0 -3.0 1e-06 
0.05 3.652 0 -3.0 1e-06 
3.0 3.652 0 -3.0 1e-06 
0.05 3.653 0 -3.0 1e-06 
3.0 3.653 0 -3.0 1e-06 
0.05 3.654 0 -3.0 1e-06 
3.0 3.654 0 -3.0 1e-06 
0.05 3.655 0 -3.0 1e-06 
3.0 3.655 0 -3.0 1e-06 
0.05 3.656 0 -3.0 1e-06 
3.0 3.656 0 -3.0 1e-06 
0.05 3.657 0 -3.0 1e-06 
3.0 3.657 0 -3.0 1e-06 
0.05 3.658 0 -3.0 1e-06 
3.0 3.658 0 -3.0 1e-06 
0.05 3.659 0 -3.0 1e-06 
3.0 3.659 0 -3.0 1e-06 
0.05 3.66 0 -3.0 1e-06 
3.0 3.66 0 -3.0 1e-06 
0.05 3.661 0 -3.0 1e-06 
3.0 3.661 0 -3.0 1e-06 
0.05 3.662 0 -3.0 1e-06 
3.0 3.662 0 -3.0 1e-06 
0.05 3.663 0 -3.0 1e-06 
3.0 3.663 0 -3.0 1e-06 
0.05 3.664 0 -3.0 1e-06 
3.0 3.664 0 -3.0 1e-06 
0.05 3.665 0 -3.0 1e-06 
3.0 3.665 0 -3.0 1e-06 
0.05 3.666 0 -3.0 1e-06 
3.0 3.666 0 -3.0 1e-06 
0.05 3.667 0 -3.0 1e-06 
3.0 3.667 0 -3.0 1e-06 
0.05 3.668 0 -3.0 1e-06 
3.0 3.668 0 -3.0 1e-06 
0.05 3.669 0 -3.0 1e-06 
3.0 3.669 0 -3.0 1e-06 
0.05 3.67 0 -3.0 1e-06 
3.0 3.67 0 -3.0 1e-06 
0.05 3.671 0 -3.0 1e-06 
3.0 3.671 0 -3.0 1e-06 
0.05 3.672 0 -3.0 1e-06 
3.0 3.672 0 -3.0 1e-06 
0.05 3.673 0 -3.0 1e-06 
3.0 3.673 0 -3.0 1e-06 
0.05 3.674 0 -3.0 1e-06 
3.0 3.674 0 -3.0 1e-06 
0.05 3.675 0 -3.0 1e-06 
3.0 3.675 0 -3.0 1e-06 
0.05 3.676 0 -3.0 1e-06 
3.0 3.676 0 -3.0 1e-06 
0.05 3.677 0 -3.0 1e-06 
3.0 3.677 0 -3.0 1e-06 
0.05 3.678 0 -3.0 1e-06 
3.0 3.678 0 -3.0 1e-06 
0.05 3.679 0 -3.0 1e-06 
3.0 3.679 0 -3.0 1e-06 
0.05 3.68 0 -3.0 1e-06 
3.0 3.68 0 -3.0 1e-06 
0.05 3.681 0 -3.0 1e-06 
3.0 3.681 0 -3.0 1e-06 
0.05 3.682 0 -3.0 1e-06 
3.0 3.682 0 -3.0 1e-06 
0.05 3.683 0 -3.0 1e-06 
3.0 3.683 0 -3.0 1e-06 
0.05 3.684 0 -3.0 1e-06 
3.0 3.684 0 -3.0 1e-06 
0.05 3.685 0 -3.0 1e-06 
3.0 3.685 0 -3.0 1e-06 
0.05 3.686 0 -3.0 1e-06 
3.0 3.686 0 -3.0 1e-06 
0.05 3.687 0 -3.0 1e-06 
3.0 3.687 0 -3.0 1e-06 
0.05 3.688 0 -3.0 1e-06 
3.0 3.688 0 -3.0 1e-06 
0.05 3.689 0 -3.0 1e-06 
3.0 3.689 0 -3.0 1e-06 
0.05 3.69 0 -3.0 1e-06 
3.0 3.69 0 -3.0 1e-06 
0.05 3.691 0 -3.0 1e-06 
3.0 3.691 0 -3.0 1e-06 
0.05 3.692 0 -3.0 1e-06 
3.0 3.692 0 -3.0 1e-06 
0.05 3.693 0 -3.0 1e-06 
3.0 3.693 0 -3.0 1e-06 
0.05 3.694 0 -3.0 1e-06 
3.0 3.694 0 -3.0 1e-06 
0.05 3.695 0 -3.0 1e-06 
3.0 3.695 0 -3.0 1e-06 
0.05 3.696 0 -3.0 1e-06 
3.0 3.696 0 -3.0 1e-06 
0.05 3.697 0 -3.0 1e-06 
3.0 3.697 0 -3.0 1e-06 
0.05 3.698 0 -3.0 1e-06 
3.0 3.698 0 -3.0 1e-06 
0.05 3.699 0 -3.0 1e-06 
3.0 3.699 0 -3.0 1e-06 
0.05 3.7 0 -3.0 1e-06 
3.0 3.7 0 -3.0 1e-06 
0.05 3.701 0 -3.0 1e-06 
3.0 3.701 0 -3.0 1e-06 
0.05 3.702 0 -3.0 1e-06 
3.0 3.702 0 -3.0 1e-06 
0.05 3.703 0 -3.0 1e-06 
3.0 3.703 0 -3.0 1e-06 
0.05 3.704 0 -3.0 1e-06 
3.0 3.704 0 -3.0 1e-06 
0.05 3.705 0 -3.0 1e-06 
3.0 3.705 0 -3.0 1e-06 
0.05 3.706 0 -3.0 1e-06 
3.0 3.706 0 -3.0 1e-06 
0.05 3.707 0 -3.0 1e-06 
3.0 3.707 0 -3.0 1e-06 
0.05 3.708 0 -3.0 1e-06 
3.0 3.708 0 -3.0 1e-06 
0.05 3.709 0 -3.0 1e-06 
3.0 3.709 0 -3.0 1e-06 
0.05 3.71 0 -3.0 1e-06 
3.0 3.71 0 -3.0 1e-06 
0.05 3.711 0 -3.0 1e-06 
3.0 3.711 0 -3.0 1e-06 
0.05 3.712 0 -3.0 1e-06 
3.0 3.712 0 -3.0 1e-06 
0.05 3.713 0 -3.0 1e-06 
3.0 3.713 0 -3.0 1e-06 
0.05 3.714 0 -3.0 1e-06 
3.0 3.714 0 -3.0 1e-06 
0.05 3.715 0 -3.0 1e-06 
3.0 3.715 0 -3.0 1e-06 
0.05 3.716 0 -3.0 1e-06 
3.0 3.716 0 -3.0 1e-06 
0.05 3.717 0 -3.0 1e-06 
3.0 3.717 0 -3.0 1e-06 
0.05 3.718 0 -3.0 1e-06 
3.0 3.718 0 -3.0 1e-06 
0.05 3.719 0 -3.0 1e-06 
3.0 3.719 0 -3.0 1e-06 
0.05 3.72 0 -3.0 1e-06 
3.0 3.72 0 -3.0 1e-06 
0.05 3.721 0 -3.0 1e-06 
3.0 3.721 0 -3.0 1e-06 
0.05 3.722 0 -3.0 1e-06 
3.0 3.722 0 -3.0 1e-06 
0.05 3.723 0 -3.0 1e-06 
3.0 3.723 0 -3.0 1e-06 
0.05 3.724 0 -3.0 1e-06 
3.0 3.724 0 -3.0 1e-06 
0.05 3.725 0 -3.0 1e-06 
3.0 3.725 0 -3.0 1e-06 
0.05 3.726 0 -3.0 1e-06 
3.0 3.726 0 -3.0 1e-06 
0.05 3.727 0 -3.0 1e-06 
3.0 3.727 0 -3.0 1e-06 
0.05 3.728 0 -3.0 1e-06 
3.0 3.728 0 -3.0 1e-06 
0.05 3.729 0 -3.0 1e-06 
3.0 3.729 0 -3.0 1e-06 
0.05 3.73 0 -3.0 1e-06 
3.0 3.73 0 -3.0 1e-06 
0.05 3.731 0 -3.0 1e-06 
3.0 3.731 0 -3.0 1e-06 
0.05 3.732 0 -3.0 1e-06 
3.0 3.732 0 -3.0 1e-06 
0.05 3.733 0 -3.0 1e-06 
3.0 3.733 0 -3.0 1e-06 
0.05 3.734 0 -3.0 1e-06 
3.0 3.734 0 -3.0 1e-06 
0.05 3.735 0 -3.0 1e-06 
3.0 3.735 0 -3.0 1e-06 
0.05 3.736 0 -3.0 1e-06 
3.0 3.736 0 -3.0 1e-06 
0.05 3.737 0 -3.0 1e-06 
3.0 3.737 0 -3.0 1e-06 
0.05 3.738 0 -3.0 1e-06 
3.0 3.738 0 -3.0 1e-06 
0.05 3.739 0 -3.0 1e-06 
3.0 3.739 0 -3.0 1e-06 
0.05 3.74 0 -3.0 1e-06 
3.0 3.74 0 -3.0 1e-06 
0.05 3.741 0 -3.0 1e-06 
3.0 3.741 0 -3.0 1e-06 
0.05 3.742 0 -3.0 1e-06 
3.0 3.742 0 -3.0 1e-06 
0.05 3.743 0 -3.0 1e-06 
3.0 3.743 0 -3.0 1e-06 
0.05 3.744 0 -3.0 1e-06 
3.0 3.744 0 -3.0 1e-06 
0.05 3.745 0 -3.0 1e-06 
3.0 3.745 0 -3.0 1e-06 
0.05 3.746 0 -3.0 1e-06 
3.0 3.746 0 -3.0 1e-06 
0.05 3.747 0 -3.0 1e-06 
3.0 3.747 0 -3.0 1e-06 
0.05 3.748 0 -3.0 1e-06 
3.0 3.748 0 -3.0 1e-06 
0.05 3.749 0 -3.0 1e-06 
3.0 3.749 0 -3.0 1e-06 
0.05 3.75 0 -3.0 1e-06 
3.0 3.75 0 -3.0 1e-06 
0.05 3.751 0 -3.0 1e-06 
3.0 3.751 0 -3.0 1e-06 
0.05 3.752 0 -3.0 1e-06 
3.0 3.752 0 -3.0 1e-06 
0.05 3.753 0 -3.0 1e-06 
3.0 3.753 0 -3.0 1e-06 
0.05 3.754 0 -3.0 1e-06 
3.0 3.754 0 -3.0 1e-06 
0.05 3.755 0 -3.0 1e-06 
3.0 3.755 0 -3.0 1e-06 
0.05 3.756 0 -3.0 1e-06 
3.0 3.756 0 -3.0 1e-06 
0.05 3.757 0 -3.0 1e-06 
3.0 3.757 0 -3.0 1e-06 
0.05 3.758 0 -3.0 1e-06 
3.0 3.758 0 -3.0 1e-06 
0.05 3.759 0 -3.0 1e-06 
3.0 3.759 0 -3.0 1e-06 
0.05 3.76 0 -3.0 1e-06 
3.0 3.76 0 -3.0 1e-06 
0.05 3.761 0 -3.0 1e-06 
3.0 3.761 0 -3.0 1e-06 
0.05 3.762 0 -3.0 1e-06 
3.0 3.762 0 -3.0 1e-06 
0.05 3.763 0 -3.0 1e-06 
3.0 3.763 0 -3.0 1e-06 
0.05 3.764 0 -3.0 1e-06 
3.0 3.764 0 -3.0 1e-06 
0.05 3.765 0 -3.0 1e-06 
3.0 3.765 0 -3.0 1e-06 
0.05 3.766 0 -3.0 1e-06 
3.0 3.766 0 -3.0 1e-06 
0.05 3.767 0 -3.0 1e-06 
3.0 3.767 0 -3.0 1e-06 
0.05 3.768 0 -3.0 1e-06 
3.0 3.768 0 -3.0 1e-06 
0.05 3.769 0 -3.0 1e-06 
3.0 3.769 0 -3.0 1e-06 
0.05 3.77 0 -3.0 1e-06 
3.0 3.77 0 -3.0 1e-06 
0.05 3.771 0 -3.0 1e-06 
3.0 3.771 0 -3.0 1e-06 
0.05 3.772 0 -3.0 1e-06 
3.0 3.772 0 -3.0 1e-06 
0.05 3.773 0 -3.0 1e-06 
3.0 3.773 0 -3.0 1e-06 
0.05 3.774 0 -3.0 1e-06 
3.0 3.774 0 -3.0 1e-06 
0.05 3.775 0 -3.0 1e-06 
3.0 3.775 0 -3.0 1e-06 
0.05 3.776 0 -3.0 1e-06 
3.0 3.776 0 -3.0 1e-06 
0.05 3.777 0 -3.0 1e-06 
3.0 3.777 0 -3.0 1e-06 
0.05 3.778 0 -3.0 1e-06 
3.0 3.778 0 -3.0 1e-06 
0.05 3.779 0 -3.0 1e-06 
3.0 3.779 0 -3.0 1e-06 
0.05 3.78 0 -3.0 1e-06 
3.0 3.78 0 -3.0 1e-06 
0.05 3.781 0 -3.0 1e-06 
3.0 3.781 0 -3.0 1e-06 
0.05 3.782 0 -3.0 1e-06 
3.0 3.782 0 -3.0 1e-06 
0.05 3.783 0 -3.0 1e-06 
3.0 3.783 0 -3.0 1e-06 
0.05 3.784 0 -3.0 1e-06 
3.0 3.784 0 -3.0 1e-06 
0.05 3.785 0 -3.0 1e-06 
3.0 3.785 0 -3.0 1e-06 
0.05 3.786 0 -3.0 1e-06 
3.0 3.786 0 -3.0 1e-06 
0.05 3.787 0 -3.0 1e-06 
3.0 3.787 0 -3.0 1e-06 
0.05 3.788 0 -3.0 1e-06 
3.0 3.788 0 -3.0 1e-06 
0.05 3.789 0 -3.0 1e-06 
3.0 3.789 0 -3.0 1e-06 
0.05 3.79 0 -3.0 1e-06 
3.0 3.79 0 -3.0 1e-06 
0.05 3.791 0 -3.0 1e-06 
3.0 3.791 0 -3.0 1e-06 
0.05 3.792 0 -3.0 1e-06 
3.0 3.792 0 -3.0 1e-06 
0.05 3.793 0 -3.0 1e-06 
3.0 3.793 0 -3.0 1e-06 
0.05 3.794 0 -3.0 1e-06 
3.0 3.794 0 -3.0 1e-06 
0.05 3.795 0 -3.0 1e-06 
3.0 3.795 0 -3.0 1e-06 
0.05 3.796 0 -3.0 1e-06 
3.0 3.796 0 -3.0 1e-06 
0.05 3.797 0 -3.0 1e-06 
3.0 3.797 0 -3.0 1e-06 
0.05 3.798 0 -3.0 1e-06 
3.0 3.798 0 -3.0 1e-06 
0.05 3.799 0 -3.0 1e-06 
3.0 3.799 0 -3.0 1e-06 
0.05 3.8 0 -3.0 1e-06 
3.0 3.8 0 -3.0 1e-06 
0.05 3.801 0 -3.0 1e-06 
3.0 3.801 0 -3.0 1e-06 
0.05 3.802 0 -3.0 1e-06 
3.0 3.802 0 -3.0 1e-06 
0.05 3.803 0 -3.0 1e-06 
3.0 3.803 0 -3.0 1e-06 
0.05 3.804 0 -3.0 1e-06 
3.0 3.804 0 -3.0 1e-06 
0.05 3.805 0 -3.0 1e-06 
3.0 3.805 0 -3.0 1e-06 
0.05 3.806 0 -3.0 1e-06 
3.0 3.806 0 -3.0 1e-06 
0.05 3.807 0 -3.0 1e-06 
3.0 3.807 0 -3.0 1e-06 
0.05 3.808 0 -3.0 1e-06 
3.0 3.808 0 -3.0 1e-06 
0.05 3.809 0 -3.0 1e-06 
3.0 3.809 0 -3.0 1e-06 
0.05 3.81 0 -3.0 1e-06 
3.0 3.81 0 -3.0 1e-06 
0.05 3.811 0 -3.0 1e-06 
3.0 3.811 0 -3.0 1e-06 
0.05 3.812 0 -3.0 1e-06 
3.0 3.812 0 -3.0 1e-06 
0.05 3.813 0 -3.0 1e-06 
3.0 3.813 0 -3.0 1e-06 
0.05 3.814 0 -3.0 1e-06 
3.0 3.814 0 -3.0 1e-06 
0.05 3.815 0 -3.0 1e-06 
3.0 3.815 0 -3.0 1e-06 
0.05 3.816 0 -3.0 1e-06 
3.0 3.816 0 -3.0 1e-06 
0.05 3.817 0 -3.0 1e-06 
3.0 3.817 0 -3.0 1e-06 
0.05 3.818 0 -3.0 1e-06 
3.0 3.818 0 -3.0 1e-06 
0.05 3.819 0 -3.0 1e-06 
3.0 3.819 0 -3.0 1e-06 
0.05 3.82 0 -3.0 1e-06 
3.0 3.82 0 -3.0 1e-06 
0.05 3.821 0 -3.0 1e-06 
3.0 3.821 0 -3.0 1e-06 
0.05 3.822 0 -3.0 1e-06 
3.0 3.822 0 -3.0 1e-06 
0.05 3.823 0 -3.0 1e-06 
3.0 3.823 0 -3.0 1e-06 
0.05 3.824 0 -3.0 1e-06 
3.0 3.824 0 -3.0 1e-06 
0.05 3.825 0 -3.0 1e-06 
3.0 3.825 0 -3.0 1e-06 
0.05 3.826 0 -3.0 1e-06 
3.0 3.826 0 -3.0 1e-06 
0.05 3.827 0 -3.0 1e-06 
3.0 3.827 0 -3.0 1e-06 
0.05 3.828 0 -3.0 1e-06 
3.0 3.828 0 -3.0 1e-06 
0.05 3.829 0 -3.0 1e-06 
3.0 3.829 0 -3.0 1e-06 
0.05 3.83 0 -3.0 1e-06 
3.0 3.83 0 -3.0 1e-06 
0.05 3.831 0 -3.0 1e-06 
3.0 3.831 0 -3.0 1e-06 
0.05 3.832 0 -3.0 1e-06 
3.0 3.832 0 -3.0 1e-06 
0.05 3.833 0 -3.0 1e-06 
3.0 3.833 0 -3.0 1e-06 
0.05 3.834 0 -3.0 1e-06 
3.0 3.834 0 -3.0 1e-06 
0.05 3.835 0 -3.0 1e-06 
3.0 3.835 0 -3.0 1e-06 
0.05 3.836 0 -3.0 1e-06 
3.0 3.836 0 -3.0 1e-06 
0.05 3.837 0 -3.0 1e-06 
3.0 3.837 0 -3.0 1e-06 
0.05 3.838 0 -3.0 1e-06 
3.0 3.838 0 -3.0 1e-06 
0.05 3.839 0 -3.0 1e-06 
3.0 3.839 0 -3.0 1e-06 
0.05 3.84 0 -3.0 1e-06 
3.0 3.84 0 -3.0 1e-06 
0.05 3.841 0 -3.0 1e-06 
3.0 3.841 0 -3.0 1e-06 
0.05 3.842 0 -3.0 1e-06 
3.0 3.842 0 -3.0 1e-06 
0.05 3.843 0 -3.0 1e-06 
3.0 3.843 0 -3.0 1e-06 
0.05 3.844 0 -3.0 1e-06 
3.0 3.844 0 -3.0 1e-06 
0.05 3.845 0 -3.0 1e-06 
3.0 3.845 0 -3.0 1e-06 
0.05 3.846 0 -3.0 1e-06 
3.0 3.846 0 -3.0 1e-06 
0.05 3.847 0 -3.0 1e-06 
3.0 3.847 0 -3.0 1e-06 
0.05 3.848 0 -3.0 1e-06 
3.0 3.848 0 -3.0 1e-06 
0.05 3.849 0 -3.0 1e-06 
3.0 3.849 0 -3.0 1e-06 
0.05 3.85 0 -3.0 1e-06 
3.0 3.85 0 -3.0 1e-06 
0.05 3.851 0 -3.0 1e-06 
3.0 3.851 0 -3.0 1e-06 
0.05 3.852 0 -3.0 1e-06 
3.0 3.852 0 -3.0 1e-06 
0.05 3.853 0 -3.0 1e-06 
3.0 3.853 0 -3.0 1e-06 
0.05 3.854 0 -3.0 1e-06 
3.0 3.854 0 -3.0 1e-06 
0.05 3.855 0 -3.0 1e-06 
3.0 3.855 0 -3.0 1e-06 
0.05 3.856 0 -3.0 1e-06 
3.0 3.856 0 -3.0 1e-06 
0.05 3.857 0 -3.0 1e-06 
3.0 3.857 0 -3.0 1e-06 
0.05 3.858 0 -3.0 1e-06 
3.0 3.858 0 -3.0 1e-06 
0.05 3.859 0 -3.0 1e-06 
3.0 3.859 0 -3.0 1e-06 
0.05 3.86 0 -3.0 1e-06 
3.0 3.86 0 -3.0 1e-06 
0.05 3.861 0 -3.0 1e-06 
3.0 3.861 0 -3.0 1e-06 
0.05 3.862 0 -3.0 1e-06 
3.0 3.862 0 -3.0 1e-06 
0.05 3.863 0 -3.0 1e-06 
3.0 3.863 0 -3.0 1e-06 
0.05 3.864 0 -3.0 1e-06 
3.0 3.864 0 -3.0 1e-06 
0.05 3.865 0 -3.0 1e-06 
3.0 3.865 0 -3.0 1e-06 
0.05 3.866 0 -3.0 1e-06 
3.0 3.866 0 -3.0 1e-06 
0.05 3.867 0 -3.0 1e-06 
3.0 3.867 0 -3.0 1e-06 
0.05 3.868 0 -3.0 1e-06 
3.0 3.868 0 -3.0 1e-06 
0.05 3.869 0 -3.0 1e-06 
3.0 3.869 0 -3.0 1e-06 
0.05 3.87 0 -3.0 1e-06 
3.0 3.87 0 -3.0 1e-06 
0.05 3.871 0 -3.0 1e-06 
3.0 3.871 0 -3.0 1e-06 
0.05 3.872 0 -3.0 1e-06 
3.0 3.872 0 -3.0 1e-06 
0.05 3.873 0 -3.0 1e-06 
3.0 3.873 0 -3.0 1e-06 
0.05 3.874 0 -3.0 1e-06 
3.0 3.874 0 -3.0 1e-06 
0.05 3.875 0 -3.0 1e-06 
3.0 3.875 0 -3.0 1e-06 
0.05 3.876 0 -3.0 1e-06 
3.0 3.876 0 -3.0 1e-06 
0.05 3.877 0 -3.0 1e-06 
3.0 3.877 0 -3.0 1e-06 
0.05 3.878 0 -3.0 1e-06 
3.0 3.878 0 -3.0 1e-06 
0.05 3.879 0 -3.0 1e-06 
3.0 3.879 0 -3.0 1e-06 
0.05 3.88 0 -3.0 1e-06 
3.0 3.88 0 -3.0 1e-06 
0.05 3.881 0 -3.0 1e-06 
3.0 3.881 0 -3.0 1e-06 
0.05 3.882 0 -3.0 1e-06 
3.0 3.882 0 -3.0 1e-06 
0.05 3.883 0 -3.0 1e-06 
3.0 3.883 0 -3.0 1e-06 
0.05 3.884 0 -3.0 1e-06 
3.0 3.884 0 -3.0 1e-06 
0.05 3.885 0 -3.0 1e-06 
3.0 3.885 0 -3.0 1e-06 
0.05 3.886 0 -3.0 1e-06 
3.0 3.886 0 -3.0 1e-06 
0.05 3.887 0 -3.0 1e-06 
3.0 3.887 0 -3.0 1e-06 
0.05 3.888 0 -3.0 1e-06 
3.0 3.888 0 -3.0 1e-06 
0.05 3.889 0 -3.0 1e-06 
3.0 3.889 0 -3.0 1e-06 
0.05 3.89 0 -3.0 1e-06 
3.0 3.89 0 -3.0 1e-06 
0.05 3.891 0 -3.0 1e-06 
3.0 3.891 0 -3.0 1e-06 
0.05 3.892 0 -3.0 1e-06 
3.0 3.892 0 -3.0 1e-06 
0.05 3.893 0 -3.0 1e-06 
3.0 3.893 0 -3.0 1e-06 
0.05 3.894 0 -3.0 1e-06 
3.0 3.894 0 -3.0 1e-06 
0.05 3.895 0 -3.0 1e-06 
3.0 3.895 0 -3.0 1e-06 
0.05 3.896 0 -3.0 1e-06 
3.0 3.896 0 -3.0 1e-06 
0.05 3.897 0 -3.0 1e-06 
3.0 3.897 0 -3.0 1e-06 
0.05 3.898 0 -3.0 1e-06 
3.0 3.898 0 -3.0 1e-06 
0.05 3.899 0 -3.0 1e-06 
3.0 3.899 0 -3.0 1e-06 
0.05 3.9 0 -3.0 1e-06 
3.0 3.9 0 -3.0 1e-06 
0.05 3.901 0 -3.0 1e-06 
3.0 3.901 0 -3.0 1e-06 
0.05 3.902 0 -3.0 1e-06 
3.0 3.902 0 -3.0 1e-06 
0.05 3.903 0 -3.0 1e-06 
3.0 3.903 0 -3.0 1e-06 
0.05 3.904 0 -3.0 1e-06 
3.0 3.904 0 -3.0 1e-06 
0.05 3.905 0 -3.0 1e-06 
3.0 3.905 0 -3.0 1e-06 
0.05 3.906 0 -3.0 1e-06 
3.0 3.906 0 -3.0 1e-06 
0.05 3.907 0 -3.0 1e-06 
3.0 3.907 0 -3.0 1e-06 
0.05 3.908 0 -3.0 1e-06 
3.0 3.908 0 -3.0 1e-06 
0.05 3.909 0 -3.0 1e-06 
3.0 3.909 0 -3.0 1e-06 
0.05 3.91 0 -3.0 1e-06 
3.0 3.91 0 -3.0 1e-06 
0.05 3.911 0 -3.0 1e-06 
3.0 3.911 0 -3.0 1e-06 
0.05 3.912 0 -3.0 1e-06 
3.0 3.912 0 -3.0 1e-06 
0.05 3.913 0 -3.0 1e-06 
3.0 3.913 0 -3.0 1e-06 
0.05 3.914 0 -3.0 1e-06 
3.0 3.914 0 -3.0 1e-06 
0.05 3.915 0 -3.0 1e-06 
3.0 3.915 0 -3.0 1e-06 
0.05 3.916 0 -3.0 1e-06 
3.0 3.916 0 -3.0 1e-06 
0.05 3.917 0 -3.0 1e-06 
3.0 3.917 0 -3.0 1e-06 
0.05 3.918 0 -3.0 1e-06 
3.0 3.918 0 -3.0 1e-06 
0.05 3.919 0 -3.0 1e-06 
3.0 3.919 0 -3.0 1e-06 
0.05 3.92 0 -3.0 1e-06 
3.0 3.92 0 -3.0 1e-06 
0.05 3.921 0 -3.0 1e-06 
3.0 3.921 0 -3.0 1e-06 
0.05 3.922 0 -3.0 1e-06 
3.0 3.922 0 -3.0 1e-06 
0.05 3.923 0 -3.0 1e-06 
3.0 3.923 0 -3.0 1e-06 
0.05 3.924 0 -3.0 1e-06 
3.0 3.924 0 -3.0 1e-06 
0.05 3.925 0 -3.0 1e-06 
3.0 3.925 0 -3.0 1e-06 
0.05 3.926 0 -3.0 1e-06 
3.0 3.926 0 -3.0 1e-06 
0.05 3.927 0 -3.0 1e-06 
3.0 3.927 0 -3.0 1e-06 
0.05 3.928 0 -3.0 1e-06 
3.0 3.928 0 -3.0 1e-06 
0.05 3.929 0 -3.0 1e-06 
3.0 3.929 0 -3.0 1e-06 
0.05 3.93 0 -3.0 1e-06 
3.0 3.93 0 -3.0 1e-06 
0.05 3.931 0 -3.0 1e-06 
3.0 3.931 0 -3.0 1e-06 
0.05 3.932 0 -3.0 1e-06 
3.0 3.932 0 -3.0 1e-06 
0.05 3.933 0 -3.0 1e-06 
3.0 3.933 0 -3.0 1e-06 
0.05 3.934 0 -3.0 1e-06 
3.0 3.934 0 -3.0 1e-06 
0.05 3.935 0 -3.0 1e-06 
3.0 3.935 0 -3.0 1e-06 
0.05 3.936 0 -3.0 1e-06 
3.0 3.936 0 -3.0 1e-06 
0.05 3.937 0 -3.0 1e-06 
3.0 3.937 0 -3.0 1e-06 
0.05 3.938 0 -3.0 1e-06 
3.0 3.938 0 -3.0 1e-06 
0.05 3.939 0 -3.0 1e-06 
3.0 3.939 0 -3.0 1e-06 
0.05 3.94 0 -3.0 1e-06 
3.0 3.94 0 -3.0 1e-06 
0.05 3.941 0 -3.0 1e-06 
3.0 3.941 0 -3.0 1e-06 
0.05 3.942 0 -3.0 1e-06 
3.0 3.942 0 -3.0 1e-06 
0.05 3.943 0 -3.0 1e-06 
3.0 3.943 0 -3.0 1e-06 
0.05 3.944 0 -3.0 1e-06 
3.0 3.944 0 -3.0 1e-06 
0.05 3.945 0 -3.0 1e-06 
3.0 3.945 0 -3.0 1e-06 
0.05 3.946 0 -3.0 1e-06 
3.0 3.946 0 -3.0 1e-06 
0.05 3.947 0 -3.0 1e-06 
3.0 3.947 0 -3.0 1e-06 
0.05 3.948 0 -3.0 1e-06 
3.0 3.948 0 -3.0 1e-06 
0.05 3.949 0 -3.0 1e-06 
3.0 3.949 0 -3.0 1e-06 
0.05 3.95 0 -3.0 1e-06 
3.0 3.95 0 -3.0 1e-06 
0.05 3.951 0 -3.0 1e-06 
3.0 3.951 0 -3.0 1e-06 
0.05 3.952 0 -3.0 1e-06 
3.0 3.952 0 -3.0 1e-06 
0.05 3.953 0 -3.0 1e-06 
3.0 3.953 0 -3.0 1e-06 
0.05 3.954 0 -3.0 1e-06 
3.0 3.954 0 -3.0 1e-06 
0.05 3.955 0 -3.0 1e-06 
3.0 3.955 0 -3.0 1e-06 
0.05 3.956 0 -3.0 1e-06 
3.0 3.956 0 -3.0 1e-06 
0.05 3.957 0 -3.0 1e-06 
3.0 3.957 0 -3.0 1e-06 
0.05 3.958 0 -3.0 1e-06 
3.0 3.958 0 -3.0 1e-06 
0.05 3.959 0 -3.0 1e-06 
3.0 3.959 0 -3.0 1e-06 
0.05 3.96 0 -3.0 1e-06 
3.0 3.96 0 -3.0 1e-06 
0.05 3.961 0 -3.0 1e-06 
3.0 3.961 0 -3.0 1e-06 
0.05 3.962 0 -3.0 1e-06 
3.0 3.962 0 -3.0 1e-06 
0.05 3.963 0 -3.0 1e-06 
3.0 3.963 0 -3.0 1e-06 
0.05 3.964 0 -3.0 1e-06 
3.0 3.964 0 -3.0 1e-06 
0.05 3.965 0 -3.0 1e-06 
3.0 3.965 0 -3.0 1e-06 
0.05 3.966 0 -3.0 1e-06 
3.0 3.966 0 -3.0 1e-06 
0.05 3.967 0 -3.0 1e-06 
3.0 3.967 0 -3.0 1e-06 
0.05 3.968 0 -3.0 1e-06 
3.0 3.968 0 -3.0 1e-06 
0.05 3.969 0 -3.0 1e-06 
3.0 3.969 0 -3.0 1e-06 
0.05 3.97 0 -3.0 1e-06 
3.0 3.97 0 -3.0 1e-06 
0.05 3.971 0 -3.0 1e-06 
3.0 3.971 0 -3.0 1e-06 
0.05 3.972 0 -3.0 1e-06 
3.0 3.972 0 -3.0 1e-06 
0.05 3.973 0 -3.0 1e-06 
3.0 3.973 0 -3.0 1e-06 
0.05 3.974 0 -3.0 1e-06 
3.0 3.974 0 -3.0 1e-06 
0.05 3.975 0 -3.0 1e-06 
3.0 3.975 0 -3.0 1e-06 
0.05 3.976 0 -3.0 1e-06 
3.0 3.976 0 -3.0 1e-06 
0.05 3.977 0 -3.0 1e-06 
3.0 3.977 0 -3.0 1e-06 
0.05 3.978 0 -3.0 1e-06 
3.0 3.978 0 -3.0 1e-06 
0.05 3.979 0 -3.0 1e-06 
3.0 3.979 0 -3.0 1e-06 
0.05 3.98 0 -3.0 1e-06 
3.0 3.98 0 -3.0 1e-06 
0.05 3.981 0 -3.0 1e-06 
3.0 3.981 0 -3.0 1e-06 
0.05 3.982 0 -3.0 1e-06 
3.0 3.982 0 -3.0 1e-06 
0.05 3.983 0 -3.0 1e-06 
3.0 3.983 0 -3.0 1e-06 
0.05 3.984 0 -3.0 1e-06 
3.0 3.984 0 -3.0 1e-06 
0.05 3.985 0 -3.0 1e-06 
3.0 3.985 0 -3.0 1e-06 
0.05 3.986 0 -3.0 1e-06 
3.0 3.986 0 -3.0 1e-06 
0.05 3.987 0 -3.0 1e-06 
3.0 3.987 0 -3.0 1e-06 
0.05 3.988 0 -3.0 1e-06 
3.0 3.988 0 -3.0 1e-06 
0.05 3.989 0 -3.0 1e-06 
3.0 3.989 0 -3.0 1e-06 
0.05 3.99 0 -3.0 1e-06 
3.0 3.99 0 -3.0 1e-06 
0.05 3.991 0 -3.0 1e-06 
3.0 3.991 0 -3.0 1e-06 
0.05 3.992 0 -3.0 1e-06 
3.0 3.992 0 -3.0 1e-06 
0.05 3.993 0 -3.0 1e-06 
3.0 3.993 0 -3.0 1e-06 
0.05 3.994 0 -3.0 1e-06 
3.0 3.994 0 -3.0 1e-06 
0.05 3.995 0 -3.0 1e-06 
3.0 3.995 0 -3.0 1e-06 
0.05 3.996 0 -3.0 1e-06 
3.0 3.996 0 -3.0 1e-06 
0.05 3.997 0 -3.0 1e-06 
3.0 3.997 0 -3.0 1e-06 
0.05 3.998 0 -3.0 1e-06 
3.0 3.998 0 -3.0 1e-06 
0.05 3.999 0 -3.0 1e-06 
3.0 3.999 0 -3.0 1e-06 
0.05 4.0 0 -3.0 1e-06 
3.0 4.0 0 -3.0 1e-06 
0.05 4.001 0 -3.0 1e-06 
3.0 4.001 0 -3.0 1e-06 
0.05 4.002 0 -3.0 1e-06 
3.0 4.002 0 -3.0 1e-06 
0.05 4.003 0 -3.0 1e-06 
3.0 4.003 0 -3.0 1e-06 
0.05 4.004 0 -3.0 1e-06 
3.0 4.004 0 -3.0 1e-06 
0.05 4.005 0 -3.0 1e-06 
3.0 4.005 0 -3.0 1e-06 
0.05 4.006 0 -3.0 1e-06 
3.0 4.006 0 -3.0 1e-06 
0.05 4.007 0 -3.0 1e-06 
3.0 4.007 0 -3.0 1e-06 
0.05 4.008 0 -3.0 1e-06 
3.0 4.008 0 -3.0 1e-06 
0.05 4.009 0 -3.0 1e-06 
3.0 4.009 0 -3.0 1e-06 
0.05 4.01 0 -3.0 1e-06 
3.0 4.01 0 -3.0 1e-06 
0.05 4.011 0 -3.0 1e-06 
3.0 4.011 0 -3.0 1e-06 
0.05 4.012 0 -3.0 1e-06 
3.0 4.012 0 -3.0 1e-06 
0.05 4.013 0 -3.0 1e-06 
3.0 4.013 0 -3.0 1e-06 
0.05 4.014 0 -3.0 1e-06 
3.0 4.014 0 -3.0 1e-06 
0.05 4.015 0 -3.0 1e-06 
3.0 4.015 0 -3.0 1e-06 
0.05 4.016 0 -3.0 1e-06 
3.0 4.016 0 -3.0 1e-06 
0.05 4.017 0 -3.0 1e-06 
3.0 4.017 0 -3.0 1e-06 
0.05 4.018 0 -3.0 1e-06 
3.0 4.018 0 -3.0 1e-06 
0.05 4.019 0 -3.0 1e-06 
3.0 4.019 0 -3.0 1e-06 
0.05 4.02 0 -3.0 1e-06 
3.0 4.02 0 -3.0 1e-06 
0.05 4.021 0 -3.0 1e-06 
3.0 4.021 0 -3.0 1e-06 
0.05 4.022 0 -3.0 1e-06 
3.0 4.022 0 -3.0 1e-06 
0.05 4.023 0 -3.0 1e-06 
3.0 4.023 0 -3.0 1e-06 
0.05 4.024 0 -3.0 1e-06 
3.0 4.024 0 -3.0 1e-06 
0.05 4.025 0 -3.0 1e-06 
3.0 4.025 0 -3.0 1e-06 
0.05 4.026 0 -3.0 1e-06 
3.0 4.026 0 -3.0 1e-06 
0.05 4.027 0 -3.0 1e-06 
3.0 4.027 0 -3.0 1e-06 
0.05 4.028 0 -3.0 1e-06 
3.0 4.028 0 -3.0 1e-06 
0.05 4.029 0 -3.0 1e-06 
3.0 4.029 0 -3.0 1e-06 
0.05 4.03 0 -3.0 1e-06 
3.0 4.03 0 -3.0 1e-06 
0.05 4.031 0 -3.0 1e-06 
3.0 4.031 0 -3.0 1e-06 
0.05 4.032 0 -3.0 1e-06 
3.0 4.032 0 -3.0 1e-06 
0.05 4.033 0 -3.0 1e-06 
3.0 4.033 0 -3.0 1e-06 
0.05 4.034 0 -3.0 1e-06 
3.0 4.034 0 -3.0 1e-06 
0.05 4.035 0 -3.0 1e-06 
3.0 4.035 0 -3.0 1e-06 
0.05 4.036 0 -3.0 1e-06 
3.0 4.036 0 -3.0 1e-06 
0.05 4.037 0 -3.0 1e-06 
3.0 4.037 0 -3.0 1e-06 
0.05 4.038 0 -3.0 1e-06 
3.0 4.038 0 -3.0 1e-06 
0.05 4.039 0 -3.0 1e-06 
3.0 4.039 0 -3.0 1e-06 
0.05 4.04 0 -3.0 1e-06 
3.0 4.04 0 -3.0 1e-06 
0.05 4.041 0 -3.0 1e-06 
3.0 4.041 0 -3.0 1e-06 
0.05 4.042 0 -3.0 1e-06 
3.0 4.042 0 -3.0 1e-06 
0.05 4.043 0 -3.0 1e-06 
3.0 4.043 0 -3.0 1e-06 
0.05 4.044 0 -3.0 1e-06 
3.0 4.044 0 -3.0 1e-06 
0.05 4.045 0 -3.0 1e-06 
3.0 4.045 0 -3.0 1e-06 
0.05 4.046 0 -3.0 1e-06 
3.0 4.046 0 -3.0 1e-06 
0.05 4.047 0 -3.0 1e-06 
3.0 4.047 0 -3.0 1e-06 
0.05 4.048 0 -3.0 1e-06 
3.0 4.048 0 -3.0 1e-06 
0.05 4.049 0 -3.0 1e-06 
3.0 4.049 0 -3.0 1e-06 
0.05 4.05 0 -3.0 1e-06 
3.0 4.05 0 -3.0 1e-06 
0.05 4.051 0 -3.0 1e-06 
3.0 4.051 0 -3.0 1e-06 
0.05 4.052 0 -3.0 1e-06 
3.0 4.052 0 -3.0 1e-06 
0.05 4.053 0 -3.0 1e-06 
3.0 4.053 0 -3.0 1e-06 
0.05 4.054 0 -3.0 1e-06 
3.0 4.054 0 -3.0 1e-06 
0.05 4.055 0 -3.0 1e-06 
3.0 4.055 0 -3.0 1e-06 
0.05 4.056 0 -3.0 1e-06 
3.0 4.056 0 -3.0 1e-06 
0.05 4.057 0 -3.0 1e-06 
3.0 4.057 0 -3.0 1e-06 
0.05 4.058 0 -3.0 1e-06 
3.0 4.058 0 -3.0 1e-06 
0.05 4.059 0 -3.0 1e-06 
3.0 4.059 0 -3.0 1e-06 
0.05 4.06 0 -3.0 1e-06 
3.0 4.06 0 -3.0 1e-06 
0.05 4.061 0 -3.0 1e-06 
3.0 4.061 0 -3.0 1e-06 
0.05 4.062 0 -3.0 1e-06 
3.0 4.062 0 -3.0 1e-06 
0.05 4.063 0 -3.0 1e-06 
3.0 4.063 0 -3.0 1e-06 
0.05 4.064 0 -3.0 1e-06 
3.0 4.064 0 -3.0 1e-06 
0.05 4.065 0 -3.0 1e-06 
3.0 4.065 0 -3.0 1e-06 
0.05 4.066 0 -3.0 1e-06 
3.0 4.066 0 -3.0 1e-06 
0.05 4.067 0 -3.0 1e-06 
3.0 4.067 0 -3.0 1e-06 
0.05 4.068 0 -3.0 1e-06 
3.0 4.068 0 -3.0 1e-06 
0.05 4.069 0 -3.0 1e-06 
3.0 4.069 0 -3.0 1e-06 
0.05 4.07 0 -3.0 1e-06 
3.0 4.07 0 -3.0 1e-06 
0.05 4.071 0 -3.0 1e-06 
3.0 4.071 0 -3.0 1e-06 
0.05 4.072 0 -3.0 1e-06 
3.0 4.072 0 -3.0 1e-06 
0.05 4.073 0 -3.0 1e-06 
3.0 4.073 0 -3.0 1e-06 
0.05 4.074 0 -3.0 1e-06 
3.0 4.074 0 -3.0 1e-06 
0.05 4.075 0 -3.0 1e-06 
3.0 4.075 0 -3.0 1e-06 
0.05 4.076 0 -3.0 1e-06 
3.0 4.076 0 -3.0 1e-06 
0.05 4.077 0 -3.0 1e-06 
3.0 4.077 0 -3.0 1e-06 
0.05 4.078 0 -3.0 1e-06 
3.0 4.078 0 -3.0 1e-06 
0.05 4.079 0 -3.0 1e-06 
3.0 4.079 0 -3.0 1e-06 
0.05 4.08 0 -3.0 1e-06 
3.0 4.08 0 -3.0 1e-06 
0.05 4.081 0 -3.0 1e-06 
3.0 4.081 0 -3.0 1e-06 
0.05 4.082 0 -3.0 1e-06 
3.0 4.082 0 -3.0 1e-06 
0.05 4.083 0 -3.0 1e-06 
3.0 4.083 0 -3.0 1e-06 
0.05 4.084 0 -3.0 1e-06 
3.0 4.084 0 -3.0 1e-06 
0.05 4.085 0 -3.0 1e-06 
3.0 4.085 0 -3.0 1e-06 
0.05 4.086 0 -3.0 1e-06 
3.0 4.086 0 -3.0 1e-06 
0.05 4.087 0 -3.0 1e-06 
3.0 4.087 0 -3.0 1e-06 
0.05 4.088 0 -3.0 1e-06 
3.0 4.088 0 -3.0 1e-06 
0.05 4.089 0 -3.0 1e-06 
3.0 4.089 0 -3.0 1e-06 
0.05 4.09 0 -3.0 1e-06 
3.0 4.09 0 -3.0 1e-06 
0.05 4.091 0 -3.0 1e-06 
3.0 4.091 0 -3.0 1e-06 
0.05 4.092 0 -3.0 1e-06 
3.0 4.092 0 -3.0 1e-06 
0.05 4.093 0 -3.0 1e-06 
3.0 4.093 0 -3.0 1e-06 
0.05 4.094 0 -3.0 1e-06 
3.0 4.094 0 -3.0 1e-06 
0.05 4.095 0 -3.0 1e-06 
3.0 4.095 0 -3.0 1e-06 
0.05 4.096 0 -3.0 1e-06 
3.0 4.096 0 -3.0 1e-06 
0.05 4.097 0 -3.0 1e-06 
3.0 4.097 0 -3.0 1e-06 
0.05 4.098 0 -3.0 1e-06 
3.0 4.098 0 -3.0 1e-06 
0.05 4.099 0 -3.0 1e-06 
3.0 4.099 0 -3.0 1e-06 
0.05 4.1 0 -3.0 1e-06 
3.0 4.1 0 -3.0 1e-06 
0.05 4.101 0 -3.0 1e-06 
3.0 4.101 0 -3.0 1e-06 
0.05 4.102 0 -3.0 1e-06 
3.0 4.102 0 -3.0 1e-06 
0.05 4.103 0 -3.0 1e-06 
3.0 4.103 0 -3.0 1e-06 
0.05 4.104 0 -3.0 1e-06 
3.0 4.104 0 -3.0 1e-06 
0.05 4.105 0 -3.0 1e-06 
3.0 4.105 0 -3.0 1e-06 
0.05 4.106 0 -3.0 1e-06 
3.0 4.106 0 -3.0 1e-06 
0.05 4.107 0 -3.0 1e-06 
3.0 4.107 0 -3.0 1e-06 
0.05 4.108 0 -3.0 1e-06 
3.0 4.108 0 -3.0 1e-06 
0.05 4.109 0 -3.0 1e-06 
3.0 4.109 0 -3.0 1e-06 
0.05 4.11 0 -3.0 1e-06 
3.0 4.11 0 -3.0 1e-06 
0.05 4.111 0 -3.0 1e-06 
3.0 4.111 0 -3.0 1e-06 
0.05 4.112 0 -3.0 1e-06 
3.0 4.112 0 -3.0 1e-06 
0.05 4.113 0 -3.0 1e-06 
3.0 4.113 0 -3.0 1e-06 
0.05 4.114 0 -3.0 1e-06 
3.0 4.114 0 -3.0 1e-06 
0.05 4.115 0 -3.0 1e-06 
3.0 4.115 0 -3.0 1e-06 
0.05 4.116 0 -3.0 1e-06 
3.0 4.116 0 -3.0 1e-06 
0.05 4.117 0 -3.0 1e-06 
3.0 4.117 0 -3.0 1e-06 
0.05 4.118 0 -3.0 1e-06 
3.0 4.118 0 -3.0 1e-06 
0.05 4.119 0 -3.0 1e-06 
3.0 4.119 0 -3.0 1e-06 
0.05 4.12 0 -3.0 1e-06 
3.0 4.12 0 -3.0 1e-06 
0.05 4.121 0 -3.0 1e-06 
3.0 4.121 0 -3.0 1e-06 
0.05 4.122 0 -3.0 1e-06 
3.0 4.122 0 -3.0 1e-06 
0.05 4.123 0 -3.0 1e-06 
3.0 4.123 0 -3.0 1e-06 
0.05 4.124 0 -3.0 1e-06 
3.0 4.124 0 -3.0 1e-06 
0.05 4.125 0 -3.0 1e-06 
3.0 4.125 0 -3.0 1e-06 
0.05 4.126 0 -3.0 1e-06 
3.0 4.126 0 -3.0 1e-06 
0.05 4.127 0 -3.0 1e-06 
3.0 4.127 0 -3.0 1e-06 
0.05 4.128 0 -3.0 1e-06 
3.0 4.128 0 -3.0 1e-06 
0.05 4.129 0 -3.0 1e-06 
3.0 4.129 0 -3.0 1e-06 
0.05 4.13 0 -3.0 1e-06 
3.0 4.13 0 -3.0 1e-06 
0.05 4.131 0 -3.0 1e-06 
3.0 4.131 0 -3.0 1e-06 
0.05 4.132 0 -3.0 1e-06 
3.0 4.132 0 -3.0 1e-06 
0.05 4.133 0 -3.0 1e-06 
3.0 4.133 0 -3.0 1e-06 
0.05 4.134 0 -3.0 1e-06 
3.0 4.134 0 -3.0 1e-06 
0.05 4.135 0 -3.0 1e-06 
3.0 4.135 0 -3.0 1e-06 
0.05 4.136 0 -3.0 1e-06 
3.0 4.136 0 -3.0 1e-06 
0.05 4.137 0 -3.0 1e-06 
3.0 4.137 0 -3.0 1e-06 
0.05 4.138 0 -3.0 1e-06 
3.0 4.138 0 -3.0 1e-06 
0.05 4.139 0 -3.0 1e-06 
3.0 4.139 0 -3.0 1e-06 
0.05 4.14 0 -3.0 1e-06 
3.0 4.14 0 -3.0 1e-06 
0.05 4.141 0 -3.0 1e-06 
3.0 4.141 0 -3.0 1e-06 
0.05 4.142 0 -3.0 1e-06 
3.0 4.142 0 -3.0 1e-06 
0.05 4.143 0 -3.0 1e-06 
3.0 4.143 0 -3.0 1e-06 
0.05 4.144 0 -3.0 1e-06 
3.0 4.144 0 -3.0 1e-06 
0.05 4.145 0 -3.0 1e-06 
3.0 4.145 0 -3.0 1e-06 
0.05 4.146 0 -3.0 1e-06 
3.0 4.146 0 -3.0 1e-06 
0.05 4.147 0 -3.0 1e-06 
3.0 4.147 0 -3.0 1e-06 
0.05 4.148 0 -3.0 1e-06 
3.0 4.148 0 -3.0 1e-06 
0.05 4.149 0 -3.0 1e-06 
3.0 4.149 0 -3.0 1e-06 
0.05 4.15 0 -3.0 1e-06 
3.0 4.15 0 -3.0 1e-06 
0.05 4.151 0 -3.0 1e-06 
3.0 4.151 0 -3.0 1e-06 
0.05 4.152 0 -3.0 1e-06 
3.0 4.152 0 -3.0 1e-06 
0.05 4.153 0 -3.0 1e-06 
3.0 4.153 0 -3.0 1e-06 
0.05 4.154 0 -3.0 1e-06 
3.0 4.154 0 -3.0 1e-06 
0.05 4.155 0 -3.0 1e-06 
3.0 4.155 0 -3.0 1e-06 
0.05 4.156 0 -3.0 1e-06 
3.0 4.156 0 -3.0 1e-06 
0.05 4.157 0 -3.0 1e-06 
3.0 4.157 0 -3.0 1e-06 
0.05 4.158 0 -3.0 1e-06 
3.0 4.158 0 -3.0 1e-06 
0.05 4.159 0 -3.0 1e-06 
3.0 4.159 0 -3.0 1e-06 
0.05 4.16 0 -3.0 1e-06 
3.0 4.16 0 -3.0 1e-06 
0.05 4.161 0 -3.0 1e-06 
3.0 4.161 0 -3.0 1e-06 
0.05 4.162 0 -3.0 1e-06 
3.0 4.162 0 -3.0 1e-06 
0.05 4.163 0 -3.0 1e-06 
3.0 4.163 0 -3.0 1e-06 
0.05 4.164 0 -3.0 1e-06 
3.0 4.164 0 -3.0 1e-06 
0.05 4.165 0 -3.0 1e-06 
3.0 4.165 0 -3.0 1e-06 
0.05 4.166 0 -3.0 1e-06 
3.0 4.166 0 -3.0 1e-06 
0.05 4.167 0 -3.0 1e-06 
3.0 4.167 0 -3.0 1e-06 
0.05 4.168 0 -3.0 1e-06 
3.0 4.168 0 -3.0 1e-06 
0.05 4.169 0 -3.0 1e-06 
3.0 4.169 0 -3.0 1e-06 
0.05 4.17 0 -3.0 1e-06 
3.0 4.17 0 -3.0 1e-06 
0.05 4.171 0 -3.0 1e-06 
3.0 4.171 0 -3.0 1e-06 
0.05 4.172 0 -3.0 1e-06 
3.0 4.172 0 -3.0 1e-06 
0.05 4.173 0 -3.0 1e-06 
3.0 4.173 0 -3.0 1e-06 
0.05 4.174 0 -3.0 1e-06 
3.0 4.174 0 -3.0 1e-06 
0.05 4.175 0 -3.0 1e-06 
3.0 4.175 0 -3.0 1e-06 
0.05 4.176 0 -3.0 1e-06 
3.0 4.176 0 -3.0 1e-06 
0.05 4.177 0 -3.0 1e-06 
3.0 4.177 0 -3.0 1e-06 
0.05 4.178 0 -3.0 1e-06 
3.0 4.178 0 -3.0 1e-06 
0.05 4.179 0 -3.0 1e-06 
3.0 4.179 0 -3.0 1e-06 
0.05 4.18 0 -3.0 1e-06 
3.0 4.18 0 -3.0 1e-06 
0.05 4.181 0 -3.0 1e-06 
3.0 4.181 0 -3.0 1e-06 
0.05 4.182 0 -3.0 1e-06 
3.0 4.182 0 -3.0 1e-06 
0.05 4.183 0 -3.0 1e-06 
3.0 4.183 0 -3.0 1e-06 
0.05 4.184 0 -3.0 1e-06 
3.0 4.184 0 -3.0 1e-06 
0.05 4.185 0 -3.0 1e-06 
3.0 4.185 0 -3.0 1e-06 
0.05 4.186 0 -3.0 1e-06 
3.0 4.186 0 -3.0 1e-06 
0.05 4.187 0 -3.0 1e-06 
3.0 4.187 0 -3.0 1e-06 
0.05 4.188 0 -3.0 1e-06 
3.0 4.188 0 -3.0 1e-06 
0.05 4.189 0 -3.0 1e-06 
3.0 4.189 0 -3.0 1e-06 
0.05 4.19 0 -3.0 1e-06 
3.0 4.19 0 -3.0 1e-06 
0.05 4.191 0 -3.0 1e-06 
3.0 4.191 0 -3.0 1e-06 
0.05 4.192 0 -3.0 1e-06 
3.0 4.192 0 -3.0 1e-06 
0.05 4.193 0 -3.0 1e-06 
3.0 4.193 0 -3.0 1e-06 
0.05 4.194 0 -3.0 1e-06 
3.0 4.194 0 -3.0 1e-06 
0.05 4.195 0 -3.0 1e-06 
3.0 4.195 0 -3.0 1e-06 
0.05 4.196 0 -3.0 1e-06 
3.0 4.196 0 -3.0 1e-06 
0.05 4.197 0 -3.0 1e-06 
3.0 4.197 0 -3.0 1e-06 
0.05 4.198 0 -3.0 1e-06 
3.0 4.198 0 -3.0 1e-06 
0.05 4.199 0 -3.0 1e-06 
3.0 4.199 0 -3.0 1e-06 
0.05 4.2 0 -3.0 1e-06 
3.0 4.2 0 -3.0 1e-06 
0.05 4.201 0 -3.0 1e-06 
3.0 4.201 0 -3.0 1e-06 
0.05 4.202 0 -3.0 1e-06 
3.0 4.202 0 -3.0 1e-06 
0.05 4.203 0 -3.0 1e-06 
3.0 4.203 0 -3.0 1e-06 
0.05 4.204 0 -3.0 1e-06 
3.0 4.204 0 -3.0 1e-06 
0.05 4.205 0 -3.0 1e-06 
3.0 4.205 0 -3.0 1e-06 
0.05 4.206 0 -3.0 1e-06 
3.0 4.206 0 -3.0 1e-06 
0.05 4.207 0 -3.0 1e-06 
3.0 4.207 0 -3.0 1e-06 
0.05 4.208 0 -3.0 1e-06 
3.0 4.208 0 -3.0 1e-06 
0.05 4.209 0 -3.0 1e-06 
3.0 4.209 0 -3.0 1e-06 
0.05 4.21 0 -3.0 1e-06 
3.0 4.21 0 -3.0 1e-06 
0.05 4.211 0 -3.0 1e-06 
3.0 4.211 0 -3.0 1e-06 
0.05 4.212 0 -3.0 1e-06 
3.0 4.212 0 -3.0 1e-06 
0.05 4.213 0 -3.0 1e-06 
3.0 4.213 0 -3.0 1e-06 
0.05 4.214 0 -3.0 1e-06 
3.0 4.214 0 -3.0 1e-06 
0.05 4.215 0 -3.0 1e-06 
3.0 4.215 0 -3.0 1e-06 
0.05 4.216 0 -3.0 1e-06 
3.0 4.216 0 -3.0 1e-06 
0.05 4.217 0 -3.0 1e-06 
3.0 4.217 0 -3.0 1e-06 
0.05 4.218 0 -3.0 1e-06 
3.0 4.218 0 -3.0 1e-06 
0.05 4.219 0 -3.0 1e-06 
3.0 4.219 0 -3.0 1e-06 
0.05 4.22 0 -3.0 1e-06 
3.0 4.22 0 -3.0 1e-06 
0.05 4.221 0 -3.0 1e-06 
3.0 4.221 0 -3.0 1e-06 
0.05 4.222 0 -3.0 1e-06 
3.0 4.222 0 -3.0 1e-06 
0.05 4.223 0 -3.0 1e-06 
3.0 4.223 0 -3.0 1e-06 
0.05 4.224 0 -3.0 1e-06 
3.0 4.224 0 -3.0 1e-06 
0.05 4.225 0 -3.0 1e-06 
3.0 4.225 0 -3.0 1e-06 
0.05 4.226 0 -3.0 1e-06 
3.0 4.226 0 -3.0 1e-06 
0.05 4.227 0 -3.0 1e-06 
3.0 4.227 0 -3.0 1e-06 
0.05 4.228 0 -3.0 1e-06 
3.0 4.228 0 -3.0 1e-06 
0.05 4.229 0 -3.0 1e-06 
3.0 4.229 0 -3.0 1e-06 
0.05 4.23 0 -3.0 1e-06 
3.0 4.23 0 -3.0 1e-06 
0.05 4.231 0 -3.0 1e-06 
3.0 4.231 0 -3.0 1e-06 
0.05 4.232 0 -3.0 1e-06 
3.0 4.232 0 -3.0 1e-06 
0.05 4.233 0 -3.0 1e-06 
3.0 4.233 0 -3.0 1e-06 
0.05 4.234 0 -3.0 1e-06 
3.0 4.234 0 -3.0 1e-06 
0.05 4.235 0 -3.0 1e-06 
3.0 4.235 0 -3.0 1e-06 
0.05 4.236 0 -3.0 1e-06 
3.0 4.236 0 -3.0 1e-06 
0.05 4.237 0 -3.0 1e-06 
3.0 4.237 0 -3.0 1e-06 
0.05 4.238 0 -3.0 1e-06 
3.0 4.238 0 -3.0 1e-06 
0.05 4.239 0 -3.0 1e-06 
3.0 4.239 0 -3.0 1e-06 
0.05 4.24 0 -3.0 1e-06 
3.0 4.24 0 -3.0 1e-06 
0.05 4.241 0 -3.0 1e-06 
3.0 4.241 0 -3.0 1e-06 
0.05 4.242 0 -3.0 1e-06 
3.0 4.242 0 -3.0 1e-06 
0.05 4.243 0 -3.0 1e-06 
3.0 4.243 0 -3.0 1e-06 
0.05 4.244 0 -3.0 1e-06 
3.0 4.244 0 -3.0 1e-06 
0.05 4.245 0 -3.0 1e-06 
3.0 4.245 0 -3.0 1e-06 
0.05 4.246 0 -3.0 1e-06 
3.0 4.246 0 -3.0 1e-06 
0.05 4.247 0 -3.0 1e-06 
3.0 4.247 0 -3.0 1e-06 
0.05 4.248 0 -3.0 1e-06 
3.0 4.248 0 -3.0 1e-06 
0.05 4.249 0 -3.0 1e-06 
3.0 4.249 0 -3.0 1e-06 
0.05 4.25 0 -3.0 1e-06 
3.0 4.25 0 -3.0 1e-06 
0.05 4.251 0 -3.0 1e-06 
3.0 4.251 0 -3.0 1e-06 
0.05 4.252 0 -3.0 1e-06 
3.0 4.252 0 -3.0 1e-06 
0.05 4.253 0 -3.0 1e-06 
3.0 4.253 0 -3.0 1e-06 
0.05 4.254 0 -3.0 1e-06 
3.0 4.254 0 -3.0 1e-06 
0.05 4.255 0 -3.0 1e-06 
3.0 4.255 0 -3.0 1e-06 
0.05 4.256 0 -3.0 1e-06 
3.0 4.256 0 -3.0 1e-06 
0.05 4.257 0 -3.0 1e-06 
3.0 4.257 0 -3.0 1e-06 
0.05 4.258 0 -3.0 1e-06 
3.0 4.258 0 -3.0 1e-06 
0.05 4.259 0 -3.0 1e-06 
3.0 4.259 0 -3.0 1e-06 
0.05 4.26 0 -3.0 1e-06 
3.0 4.26 0 -3.0 1e-06 
0.05 4.261 0 -3.0 1e-06 
3.0 4.261 0 -3.0 1e-06 
0.05 4.262 0 -3.0 1e-06 
3.0 4.262 0 -3.0 1e-06 
0.05 4.263 0 -3.0 1e-06 
3.0 4.263 0 -3.0 1e-06 
0.05 4.264 0 -3.0 1e-06 
3.0 4.264 0 -3.0 1e-06 
0.05 4.265 0 -3.0 1e-06 
3.0 4.265 0 -3.0 1e-06 
0.05 4.266 0 -3.0 1e-06 
3.0 4.266 0 -3.0 1e-06 
0.05 4.267 0 -3.0 1e-06 
3.0 4.267 0 -3.0 1e-06 
0.05 4.268 0 -3.0 1e-06 
3.0 4.268 0 -3.0 1e-06 
0.05 4.269 0 -3.0 1e-06 
3.0 4.269 0 -3.0 1e-06 
0.05 4.27 0 -3.0 1e-06 
3.0 4.27 0 -3.0 1e-06 
0.05 4.271 0 -3.0 1e-06 
3.0 4.271 0 -3.0 1e-06 
0.05 4.272 0 -3.0 1e-06 
3.0 4.272 0 -3.0 1e-06 
0.05 4.273 0 -3.0 1e-06 
3.0 4.273 0 -3.0 1e-06 
0.05 4.274 0 -3.0 1e-06 
3.0 4.274 0 -3.0 1e-06 
0.05 4.275 0 -3.0 1e-06 
3.0 4.275 0 -3.0 1e-06 
0.05 4.276 0 -3.0 1e-06 
3.0 4.276 0 -3.0 1e-06 
0.05 4.277 0 -3.0 1e-06 
3.0 4.277 0 -3.0 1e-06 
0.05 4.278 0 -3.0 1e-06 
3.0 4.278 0 -3.0 1e-06 
0.05 4.279 0 -3.0 1e-06 
3.0 4.279 0 -3.0 1e-06 
0.05 4.28 0 -3.0 1e-06 
3.0 4.28 0 -3.0 1e-06 
0.05 4.281 0 -3.0 1e-06 
3.0 4.281 0 -3.0 1e-06 
0.05 4.282 0 -3.0 1e-06 
3.0 4.282 0 -3.0 1e-06 
0.05 4.283 0 -3.0 1e-06 
3.0 4.283 0 -3.0 1e-06 
0.05 4.284 0 -3.0 1e-06 
3.0 4.284 0 -3.0 1e-06 
0.05 4.285 0 -3.0 1e-06 
3.0 4.285 0 -3.0 1e-06 
0.05 4.286 0 -3.0 1e-06 
3.0 4.286 0 -3.0 1e-06 
0.05 4.287 0 -3.0 1e-06 
3.0 4.287 0 -3.0 1e-06 
0.05 4.288 0 -3.0 1e-06 
3.0 4.288 0 -3.0 1e-06 
0.05 4.289 0 -3.0 1e-06 
3.0 4.289 0 -3.0 1e-06 
0.05 4.29 0 -3.0 1e-06 
3.0 4.29 0 -3.0 1e-06 
0.05 4.291 0 -3.0 1e-06 
3.0 4.291 0 -3.0 1e-06 
0.05 4.292 0 -3.0 1e-06 
3.0 4.292 0 -3.0 1e-06 
0.05 4.293 0 -3.0 1e-06 
3.0 4.293 0 -3.0 1e-06 
0.05 4.294 0 -3.0 1e-06 
3.0 4.294 0 -3.0 1e-06 
0.05 4.295 0 -3.0 1e-06 
3.0 4.295 0 -3.0 1e-06 
0.05 4.296 0 -3.0 1e-06 
3.0 4.296 0 -3.0 1e-06 
0.05 4.297 0 -3.0 1e-06 
3.0 4.297 0 -3.0 1e-06 
0.05 4.298 0 -3.0 1e-06 
3.0 4.298 0 -3.0 1e-06 
0.05 4.299 0 -3.0 1e-06 
3.0 4.299 0 -3.0 1e-06 
0.05 4.3 0 -3.0 1e-06 
3.0 4.3 0 -3.0 1e-06 
0.05 4.301 0 -3.0 1e-06 
3.0 4.301 0 -3.0 1e-06 
0.05 4.302 0 -3.0 1e-06 
3.0 4.302 0 -3.0 1e-06 
0.05 4.303 0 -3.0 1e-06 
3.0 4.303 0 -3.0 1e-06 
0.05 4.304 0 -3.0 1e-06 
3.0 4.304 0 -3.0 1e-06 
0.05 4.305 0 -3.0 1e-06 
3.0 4.305 0 -3.0 1e-06 
0.05 4.306 0 -3.0 1e-06 
3.0 4.306 0 -3.0 1e-06 
0.05 4.307 0 -3.0 1e-06 
3.0 4.307 0 -3.0 1e-06 
0.05 4.308 0 -3.0 1e-06 
3.0 4.308 0 -3.0 1e-06 
0.05 4.309 0 -3.0 1e-06 
3.0 4.309 0 -3.0 1e-06 
0.05 4.31 0 -3.0 1e-06 
3.0 4.31 0 -3.0 1e-06 
0.05 4.311 0 -3.0 1e-06 
3.0 4.311 0 -3.0 1e-06 
0.05 4.312 0 -3.0 1e-06 
3.0 4.312 0 -3.0 1e-06 
0.05 4.313 0 -3.0 1e-06 
3.0 4.313 0 -3.0 1e-06 
0.05 4.314 0 -3.0 1e-06 
3.0 4.314 0 -3.0 1e-06 
0.05 4.315 0 -3.0 1e-06 
3.0 4.315 0 -3.0 1e-06 
0.05 4.316 0 -3.0 1e-06 
3.0 4.316 0 -3.0 1e-06 
0.05 4.317 0 -3.0 1e-06 
3.0 4.317 0 -3.0 1e-06 
0.05 4.318 0 -3.0 1e-06 
3.0 4.318 0 -3.0 1e-06 
0.05 4.319 0 -3.0 1e-06 
3.0 4.319 0 -3.0 1e-06 
0.05 4.32 0 -3.0 1e-06 
3.0 4.32 0 -3.0 1e-06 
0.05 4.321 0 -3.0 1e-06 
3.0 4.321 0 -3.0 1e-06 
0.05 4.322 0 -3.0 1e-06 
3.0 4.322 0 -3.0 1e-06 
0.05 4.323 0 -3.0 1e-06 
3.0 4.323 0 -3.0 1e-06 
0.05 4.324 0 -3.0 1e-06 
3.0 4.324 0 -3.0 1e-06 
0.05 4.325 0 -3.0 1e-06 
3.0 4.325 0 -3.0 1e-06 
0.05 4.326 0 -3.0 1e-06 
3.0 4.326 0 -3.0 1e-06 
0.05 4.327 0 -3.0 1e-06 
3.0 4.327 0 -3.0 1e-06 
0.05 4.328 0 -3.0 1e-06 
3.0 4.328 0 -3.0 1e-06 
0.05 4.329 0 -3.0 1e-06 
3.0 4.329 0 -3.0 1e-06 
0.05 4.33 0 -3.0 1e-06 
3.0 4.33 0 -3.0 1e-06 
0.05 4.331 0 -3.0 1e-06 
3.0 4.331 0 -3.0 1e-06 
0.05 4.332 0 -3.0 1e-06 
3.0 4.332 0 -3.0 1e-06 
0.05 4.333 0 -3.0 1e-06 
3.0 4.333 0 -3.0 1e-06 
0.05 4.334 0 -3.0 1e-06 
3.0 4.334 0 -3.0 1e-06 
0.05 4.335 0 -3.0 1e-06 
3.0 4.335 0 -3.0 1e-06 
0.05 4.336 0 -3.0 1e-06 
3.0 4.336 0 -3.0 1e-06 
0.05 4.337 0 -3.0 1e-06 
3.0 4.337 0 -3.0 1e-06 
0.05 4.338 0 -3.0 1e-06 
3.0 4.338 0 -3.0 1e-06 
0.05 4.339 0 -3.0 1e-06 
3.0 4.339 0 -3.0 1e-06 
0.05 4.34 0 -3.0 1e-06 
3.0 4.34 0 -3.0 1e-06 
0.05 4.341 0 -3.0 1e-06 
3.0 4.341 0 -3.0 1e-06 
0.05 4.342 0 -3.0 1e-06 
3.0 4.342 0 -3.0 1e-06 
0.05 4.343 0 -3.0 1e-06 
3.0 4.343 0 -3.0 1e-06 
0.05 4.344 0 -3.0 1e-06 
3.0 4.344 0 -3.0 1e-06 
0.05 4.345 0 -3.0 1e-06 
3.0 4.345 0 -3.0 1e-06 
0.05 4.346 0 -3.0 1e-06 
3.0 4.346 0 -3.0 1e-06 
0.05 4.347 0 -3.0 1e-06 
3.0 4.347 0 -3.0 1e-06 
0.05 4.348 0 -3.0 1e-06 
3.0 4.348 0 -3.0 1e-06 
0.05 4.349 0 -3.0 1e-06 
3.0 4.349 0 -3.0 1e-06 
0.05 4.35 0 -3.0 1e-06 
3.0 4.35 0 -3.0 1e-06 
0.05 4.351 0 -3.0 1e-06 
3.0 4.351 0 -3.0 1e-06 
0.05 4.352 0 -3.0 1e-06 
3.0 4.352 0 -3.0 1e-06 
0.05 4.353 0 -3.0 1e-06 
3.0 4.353 0 -3.0 1e-06 
0.05 4.354 0 -3.0 1e-06 
3.0 4.354 0 -3.0 1e-06 
0.05 4.355 0 -3.0 1e-06 
3.0 4.355 0 -3.0 1e-06 
0.05 4.356 0 -3.0 1e-06 
3.0 4.356 0 -3.0 1e-06 
0.05 4.357 0 -3.0 1e-06 
3.0 4.357 0 -3.0 1e-06 
0.05 4.358 0 -3.0 1e-06 
3.0 4.358 0 -3.0 1e-06 
0.05 4.359 0 -3.0 1e-06 
3.0 4.359 0 -3.0 1e-06 
0.05 4.36 0 -3.0 1e-06 
3.0 4.36 0 -3.0 1e-06 
0.05 4.361 0 -3.0 1e-06 
3.0 4.361 0 -3.0 1e-06 
0.05 4.362 0 -3.0 1e-06 
3.0 4.362 0 -3.0 1e-06 
0.05 4.363 0 -3.0 1e-06 
3.0 4.363 0 -3.0 1e-06 
0.05 4.364 0 -3.0 1e-06 
3.0 4.364 0 -3.0 1e-06 
0.05 4.365 0 -3.0 1e-06 
3.0 4.365 0 -3.0 1e-06 
0.05 4.366 0 -3.0 1e-06 
3.0 4.366 0 -3.0 1e-06 
0.05 4.367 0 -3.0 1e-06 
3.0 4.367 0 -3.0 1e-06 
0.05 4.368 0 -3.0 1e-06 
3.0 4.368 0 -3.0 1e-06 
0.05 4.369 0 -3.0 1e-06 
3.0 4.369 0 -3.0 1e-06 
0.05 4.37 0 -3.0 1e-06 
3.0 4.37 0 -3.0 1e-06 
0.05 4.371 0 -3.0 1e-06 
3.0 4.371 0 -3.0 1e-06 
0.05 4.372 0 -3.0 1e-06 
3.0 4.372 0 -3.0 1e-06 
0.05 4.373 0 -3.0 1e-06 
3.0 4.373 0 -3.0 1e-06 
0.05 4.374 0 -3.0 1e-06 
3.0 4.374 0 -3.0 1e-06 
0.05 4.375 0 -3.0 1e-06 
3.0 4.375 0 -3.0 1e-06 
0.05 4.376 0 -3.0 1e-06 
3.0 4.376 0 -3.0 1e-06 
0.05 4.377 0 -3.0 1e-06 
3.0 4.377 0 -3.0 1e-06 
0.05 4.378 0 -3.0 1e-06 
3.0 4.378 0 -3.0 1e-06 
0.05 4.379 0 -3.0 1e-06 
3.0 4.379 0 -3.0 1e-06 
0.05 4.38 0 -3.0 1e-06 
3.0 4.38 0 -3.0 1e-06 
0.05 4.381 0 -3.0 1e-06 
3.0 4.381 0 -3.0 1e-06 
0.05 4.382 0 -3.0 1e-06 
3.0 4.382 0 -3.0 1e-06 
0.05 4.383 0 -3.0 1e-06 
3.0 4.383 0 -3.0 1e-06 
0.05 4.384 0 -3.0 1e-06 
3.0 4.384 0 -3.0 1e-06 
0.05 4.385 0 -3.0 1e-06 
3.0 4.385 0 -3.0 1e-06 
0.05 4.386 0 -3.0 1e-06 
3.0 4.386 0 -3.0 1e-06 
0.05 4.387 0 -3.0 1e-06 
3.0 4.387 0 -3.0 1e-06 
0.05 4.388 0 -3.0 1e-06 
3.0 4.388 0 -3.0 1e-06 
0.05 4.389 0 -3.0 1e-06 
3.0 4.389 0 -3.0 1e-06 
0.05 4.39 0 -3.0 1e-06 
3.0 4.39 0 -3.0 1e-06 
0.05 4.391 0 -3.0 1e-06 
3.0 4.391 0 -3.0 1e-06 
0.05 4.392 0 -3.0 1e-06 
3.0 4.392 0 -3.0 1e-06 
0.05 4.393 0 -3.0 1e-06 
3.0 4.393 0 -3.0 1e-06 
0.05 4.394 0 -3.0 1e-06 
3.0 4.394 0 -3.0 1e-06 
0.05 4.395 0 -3.0 1e-06 
3.0 4.395 0 -3.0 1e-06 
0.05 4.396 0 -3.0 1e-06 
3.0 4.396 0 -3.0 1e-06 
0.05 4.397 0 -3.0 1e-06 
3.0 4.397 0 -3.0 1e-06 
0.05 4.398 0 -3.0 1e-06 
3.0 4.398 0 -3.0 1e-06 
0.05 4.399 0 -3.0 1e-06 
3.0 4.399 0 -3.0 1e-06 
0.05 4.4 0 -3.0 1e-06 
3.0 4.4 0 -3.0 1e-06 
0.05 4.401 0 -3.0 1e-06 
3.0 4.401 0 -3.0 1e-06 
0.05 4.402 0 -3.0 1e-06 
3.0 4.402 0 -3.0 1e-06 
0.05 4.403 0 -3.0 1e-06 
3.0 4.403 0 -3.0 1e-06 
0.05 4.404 0 -3.0 1e-06 
3.0 4.404 0 -3.0 1e-06 
0.05 4.405 0 -3.0 1e-06 
3.0 4.405 0 -3.0 1e-06 
0.05 4.406 0 -3.0 1e-06 
3.0 4.406 0 -3.0 1e-06 
0.05 4.407 0 -3.0 1e-06 
3.0 4.407 0 -3.0 1e-06 
0.05 4.408 0 -3.0 1e-06 
3.0 4.408 0 -3.0 1e-06 
0.05 4.409 0 -3.0 1e-06 
3.0 4.409 0 -3.0 1e-06 
0.05 4.41 0 -3.0 1e-06 
3.0 4.41 0 -3.0 1e-06 
0.05 4.411 0 -3.0 1e-06 
3.0 4.411 0 -3.0 1e-06 
0.05 4.412 0 -3.0 1e-06 
3.0 4.412 0 -3.0 1e-06 
0.05 4.413 0 -3.0 1e-06 
3.0 4.413 0 -3.0 1e-06 
0.05 4.414 0 -3.0 1e-06 
3.0 4.414 0 -3.0 1e-06 
0.05 4.415 0 -3.0 1e-06 
3.0 4.415 0 -3.0 1e-06 
0.05 4.416 0 -3.0 1e-06 
3.0 4.416 0 -3.0 1e-06 
0.05 4.417 0 -3.0 1e-06 
3.0 4.417 0 -3.0 1e-06 
0.05 4.418 0 -3.0 1e-06 
3.0 4.418 0 -3.0 1e-06 
0.05 4.419 0 -3.0 1e-06 
3.0 4.419 0 -3.0 1e-06 
0.05 4.42 0 -3.0 1e-06 
3.0 4.42 0 -3.0 1e-06 
0.05 4.421 0 -3.0 1e-06 
3.0 4.421 0 -3.0 1e-06 
0.05 4.422 0 -3.0 1e-06 
3.0 4.422 0 -3.0 1e-06 
0.05 4.423 0 -3.0 1e-06 
3.0 4.423 0 -3.0 1e-06 
0.05 4.424 0 -3.0 1e-06 
3.0 4.424 0 -3.0 1e-06 
0.05 4.425 0 -3.0 1e-06 
3.0 4.425 0 -3.0 1e-06 
0.05 4.426 0 -3.0 1e-06 
3.0 4.426 0 -3.0 1e-06 
0.05 4.427 0 -3.0 1e-06 
3.0 4.427 0 -3.0 1e-06 
0.05 4.428 0 -3.0 1e-06 
3.0 4.428 0 -3.0 1e-06 
0.05 4.429 0 -3.0 1e-06 
3.0 4.429 0 -3.0 1e-06 
0.05 4.43 0 -3.0 1e-06 
3.0 4.43 0 -3.0 1e-06 
0.05 4.431 0 -3.0 1e-06 
3.0 4.431 0 -3.0 1e-06 
0.05 4.432 0 -3.0 1e-06 
3.0 4.432 0 -3.0 1e-06 
0.05 4.433 0 -3.0 1e-06 
3.0 4.433 0 -3.0 1e-06 
0.05 4.434 0 -3.0 1e-06 
3.0 4.434 0 -3.0 1e-06 
0.05 4.435 0 -3.0 1e-06 
3.0 4.435 0 -3.0 1e-06 
0.05 4.436 0 -3.0 1e-06 
3.0 4.436 0 -3.0 1e-06 
0.05 4.437 0 -3.0 1e-06 
3.0 4.437 0 -3.0 1e-06 
0.05 4.438 0 -3.0 1e-06 
3.0 4.438 0 -3.0 1e-06 
0.05 4.439 0 -3.0 1e-06 
3.0 4.439 0 -3.0 1e-06 
0.05 4.44 0 -3.0 1e-06 
3.0 4.44 0 -3.0 1e-06 
0.05 4.441 0 -3.0 1e-06 
3.0 4.441 0 -3.0 1e-06 
0.05 4.442 0 -3.0 1e-06 
3.0 4.442 0 -3.0 1e-06 
0.05 4.443 0 -3.0 1e-06 
3.0 4.443 0 -3.0 1e-06 
0.05 4.444 0 -3.0 1e-06 
3.0 4.444 0 -3.0 1e-06 
0.05 4.445 0 -3.0 1e-06 
3.0 4.445 0 -3.0 1e-06 
0.05 4.446 0 -3.0 1e-06 
3.0 4.446 0 -3.0 1e-06 
0.05 4.447 0 -3.0 1e-06 
3.0 4.447 0 -3.0 1e-06 
0.05 4.448 0 -3.0 1e-06 
3.0 4.448 0 -3.0 1e-06 
0.05 4.449 0 -3.0 1e-06 
3.0 4.449 0 -3.0 1e-06 
0.05 4.45 0 -3.0 1e-06 
3.0 4.45 0 -3.0 1e-06 
0.05 4.451 0 -3.0 1e-06 
3.0 4.451 0 -3.0 1e-06 
0.05 4.452 0 -3.0 1e-06 
3.0 4.452 0 -3.0 1e-06 
0.05 4.453 0 -3.0 1e-06 
3.0 4.453 0 -3.0 1e-06 
0.05 4.454 0 -3.0 1e-06 
3.0 4.454 0 -3.0 1e-06 
0.05 4.455 0 -3.0 1e-06 
3.0 4.455 0 -3.0 1e-06 
0.05 4.456 0 -3.0 1e-06 
3.0 4.456 0 -3.0 1e-06 
0.05 4.457 0 -3.0 1e-06 
3.0 4.457 0 -3.0 1e-06 
0.05 4.458 0 -3.0 1e-06 
3.0 4.458 0 -3.0 1e-06 
0.05 4.459 0 -3.0 1e-06 
3.0 4.459 0 -3.0 1e-06 
0.05 4.46 0 -3.0 1e-06 
3.0 4.46 0 -3.0 1e-06 
0.05 4.461 0 -3.0 1e-06 
3.0 4.461 0 -3.0 1e-06 
0.05 4.462 0 -3.0 1e-06 
3.0 4.462 0 -3.0 1e-06 
0.05 4.463 0 -3.0 1e-06 
3.0 4.463 0 -3.0 1e-06 
0.05 4.464 0 -3.0 1e-06 
3.0 4.464 0 -3.0 1e-06 
0.05 4.465 0 -3.0 1e-06 
3.0 4.465 0 -3.0 1e-06 
0.05 4.466 0 -3.0 1e-06 
3.0 4.466 0 -3.0 1e-06 
0.05 4.467 0 -3.0 1e-06 
3.0 4.467 0 -3.0 1e-06 
0.05 4.468 0 -3.0 1e-06 
3.0 4.468 0 -3.0 1e-06 
0.05 4.469 0 -3.0 1e-06 
3.0 4.469 0 -3.0 1e-06 
0.05 4.47 0 -3.0 1e-06 
3.0 4.47 0 -3.0 1e-06 
0.05 4.471 0 -3.0 1e-06 
3.0 4.471 0 -3.0 1e-06 
0.05 4.472 0 -3.0 1e-06 
3.0 4.472 0 -3.0 1e-06 
0.05 4.473 0 -3.0 1e-06 
3.0 4.473 0 -3.0 1e-06 
0.05 4.474 0 -3.0 1e-06 
3.0 4.474 0 -3.0 1e-06 
0.05 4.475 0 -3.0 1e-06 
3.0 4.475 0 -3.0 1e-06 
0.05 4.476 0 -3.0 1e-06 
3.0 4.476 0 -3.0 1e-06 
0.05 4.477 0 -3.0 1e-06 
3.0 4.477 0 -3.0 1e-06 
0.05 4.478 0 -3.0 1e-06 
3.0 4.478 0 -3.0 1e-06 
0.05 4.479 0 -3.0 1e-06 
3.0 4.479 0 -3.0 1e-06 
0.05 4.48 0 -3.0 1e-06 
3.0 4.48 0 -3.0 1e-06 
0.05 4.481 0 -3.0 1e-06 
3.0 4.481 0 -3.0 1e-06 
0.05 4.482 0 -3.0 1e-06 
3.0 4.482 0 -3.0 1e-06 
0.05 4.483 0 -3.0 1e-06 
3.0 4.483 0 -3.0 1e-06 
0.05 4.484 0 -3.0 1e-06 
3.0 4.484 0 -3.0 1e-06 
0.05 4.485 0 -3.0 1e-06 
3.0 4.485 0 -3.0 1e-06 
0.05 4.486 0 -3.0 1e-06 
3.0 4.486 0 -3.0 1e-06 
0.05 4.487 0 -3.0 1e-06 
3.0 4.487 0 -3.0 1e-06 
0.05 4.488 0 -3.0 1e-06 
3.0 4.488 0 -3.0 1e-06 
0.05 4.489 0 -3.0 1e-06 
3.0 4.489 0 -3.0 1e-06 
0.05 4.49 0 -3.0 1e-06 
3.0 4.49 0 -3.0 1e-06 
0.05 4.491 0 -3.0 1e-06 
3.0 4.491 0 -3.0 1e-06 
0.05 4.492 0 -3.0 1e-06 
3.0 4.492 0 -3.0 1e-06 
0.05 4.493 0 -3.0 1e-06 
3.0 4.493 0 -3.0 1e-06 
0.05 4.494 0 -3.0 1e-06 
3.0 4.494 0 -3.0 1e-06 
0.05 4.495 0 -3.0 1e-06 
3.0 4.495 0 -3.0 1e-06 
0.05 4.496 0 -3.0 1e-06 
3.0 4.496 0 -3.0 1e-06 
0.05 4.497 0 -3.0 1e-06 
3.0 4.497 0 -3.0 1e-06 
0.05 4.498 0 -3.0 1e-06 
3.0 4.498 0 -3.0 1e-06 
0.05 4.499 0 -3.0 1e-06 
3.0 4.499 0 -3.0 1e-06 
0.05 4.5 0 -3.0 1e-06 
3.0 4.5 0 -3.0 1e-06 
0.05 4.501 0 -3.0 1e-06 
3.0 4.501 0 -3.0 1e-06 
0.05 4.502 0 -3.0 1e-06 
3.0 4.502 0 -3.0 1e-06 
0.05 4.503 0 -3.0 1e-06 
3.0 4.503 0 -3.0 1e-06 
0.05 4.504 0 -3.0 1e-06 
3.0 4.504 0 -3.0 1e-06 
0.05 4.505 0 -3.0 1e-06 
3.0 4.505 0 -3.0 1e-06 
0.05 4.506 0 -3.0 1e-06 
3.0 4.506 0 -3.0 1e-06 
0.05 4.507 0 -3.0 1e-06 
3.0 4.507 0 -3.0 1e-06 
0.05 4.508 0 -3.0 1e-06 
3.0 4.508 0 -3.0 1e-06 
0.05 4.509 0 -3.0 1e-06 
3.0 4.509 0 -3.0 1e-06 
0.05 4.51 0 -3.0 1e-06 
3.0 4.51 0 -3.0 1e-06 
0.05 4.511 0 -3.0 1e-06 
3.0 4.511 0 -3.0 1e-06 
0.05 4.512 0 -3.0 1e-06 
3.0 4.512 0 -3.0 1e-06 
0.05 4.513 0 -3.0 1e-06 
3.0 4.513 0 -3.0 1e-06 
0.05 4.514 0 -3.0 1e-06 
3.0 4.514 0 -3.0 1e-06 
0.05 4.515 0 -3.0 1e-06 
3.0 4.515 0 -3.0 1e-06 
0.05 4.516 0 -3.0 1e-06 
3.0 4.516 0 -3.0 1e-06 
0.05 4.517 0 -3.0 1e-06 
3.0 4.517 0 -3.0 1e-06 
0.05 4.518 0 -3.0 1e-06 
3.0 4.518 0 -3.0 1e-06 
0.05 4.519 0 -3.0 1e-06 
3.0 4.519 0 -3.0 1e-06 
0.05 4.52 0 -3.0 1e-06 
3.0 4.52 0 -3.0 1e-06 
0.05 4.521 0 -3.0 1e-06 
3.0 4.521 0 -3.0 1e-06 
0.05 4.522 0 -3.0 1e-06 
3.0 4.522 0 -3.0 1e-06 
0.05 4.523 0 -3.0 1e-06 
3.0 4.523 0 -3.0 1e-06 
0.05 4.524 0 -3.0 1e-06 
3.0 4.524 0 -3.0 1e-06 
0.05 4.525 0 -3.0 1e-06 
3.0 4.525 0 -3.0 1e-06 
0.05 4.526 0 -3.0 1e-06 
3.0 4.526 0 -3.0 1e-06 
0.05 4.527 0 -3.0 1e-06 
3.0 4.527 0 -3.0 1e-06 
0.05 4.528 0 -3.0 1e-06 
3.0 4.528 0 -3.0 1e-06 
0.05 4.529 0 -3.0 1e-06 
3.0 4.529 0 -3.0 1e-06 
0.05 4.53 0 -3.0 1e-06 
3.0 4.53 0 -3.0 1e-06 
0.05 4.531 0 -3.0 1e-06 
3.0 4.531 0 -3.0 1e-06 
0.05 4.532 0 -3.0 1e-06 
3.0 4.532 0 -3.0 1e-06 
0.05 4.533 0 -3.0 1e-06 
3.0 4.533 0 -3.0 1e-06 
0.05 4.534 0 -3.0 1e-06 
3.0 4.534 0 -3.0 1e-06 
0.05 4.535 0 -3.0 1e-06 
3.0 4.535 0 -3.0 1e-06 
0.05 4.536 0 -3.0 1e-06 
3.0 4.536 0 -3.0 1e-06 
0.05 4.537 0 -3.0 1e-06 
3.0 4.537 0 -3.0 1e-06 
0.05 4.538 0 -3.0 1e-06 
3.0 4.538 0 -3.0 1e-06 
0.05 4.539 0 -3.0 1e-06 
3.0 4.539 0 -3.0 1e-06 
0.05 4.54 0 -3.0 1e-06 
3.0 4.54 0 -3.0 1e-06 
0.05 4.541 0 -3.0 1e-06 
3.0 4.541 0 -3.0 1e-06 
0.05 4.542 0 -3.0 1e-06 
3.0 4.542 0 -3.0 1e-06 
0.05 4.543 0 -3.0 1e-06 
3.0 4.543 0 -3.0 1e-06 
0.05 4.544 0 -3.0 1e-06 
3.0 4.544 0 -3.0 1e-06 
0.05 4.545 0 -3.0 1e-06 
3.0 4.545 0 -3.0 1e-06 
0.05 4.546 0 -3.0 1e-06 
3.0 4.546 0 -3.0 1e-06 
0.05 4.547 0 -3.0 1e-06 
3.0 4.547 0 -3.0 1e-06 
0.05 4.548 0 -3.0 1e-06 
3.0 4.548 0 -3.0 1e-06 
0.05 4.549 0 -3.0 1e-06 
3.0 4.549 0 -3.0 1e-06 
0.05 4.55 0 -3.0 1e-06 
3.0 4.55 0 -3.0 1e-06 
0.05 4.551 0 -3.0 1e-06 
3.0 4.551 0 -3.0 1e-06 
0.05 4.552 0 -3.0 1e-06 
3.0 4.552 0 -3.0 1e-06 
0.05 4.553 0 -3.0 1e-06 
3.0 4.553 0 -3.0 1e-06 
0.05 4.554 0 -3.0 1e-06 
3.0 4.554 0 -3.0 1e-06 
0.05 4.555 0 -3.0 1e-06 
3.0 4.555 0 -3.0 1e-06 
0.05 4.556 0 -3.0 1e-06 
3.0 4.556 0 -3.0 1e-06 
0.05 4.557 0 -3.0 1e-06 
3.0 4.557 0 -3.0 1e-06 
0.05 4.558 0 -3.0 1e-06 
3.0 4.558 0 -3.0 1e-06 
0.05 4.559 0 -3.0 1e-06 
3.0 4.559 0 -3.0 1e-06 
0.05 4.56 0 -3.0 1e-06 
3.0 4.56 0 -3.0 1e-06 
0.05 4.561 0 -3.0 1e-06 
3.0 4.561 0 -3.0 1e-06 
0.05 4.562 0 -3.0 1e-06 
3.0 4.562 0 -3.0 1e-06 
0.05 4.563 0 -3.0 1e-06 
3.0 4.563 0 -3.0 1e-06 
0.05 4.564 0 -3.0 1e-06 
3.0 4.564 0 -3.0 1e-06 
0.05 4.565 0 -3.0 1e-06 
3.0 4.565 0 -3.0 1e-06 
0.05 4.566 0 -3.0 1e-06 
3.0 4.566 0 -3.0 1e-06 
0.05 4.567 0 -3.0 1e-06 
3.0 4.567 0 -3.0 1e-06 
0.05 4.568 0 -3.0 1e-06 
3.0 4.568 0 -3.0 1e-06 
0.05 4.569 0 -3.0 1e-06 
3.0 4.569 0 -3.0 1e-06 
0.05 4.57 0 -3.0 1e-06 
3.0 4.57 0 -3.0 1e-06 
0.05 4.571 0 -3.0 1e-06 
3.0 4.571 0 -3.0 1e-06 
0.05 4.572 0 -3.0 1e-06 
3.0 4.572 0 -3.0 1e-06 
0.05 4.573 0 -3.0 1e-06 
3.0 4.573 0 -3.0 1e-06 
0.05 4.574 0 -3.0 1e-06 
3.0 4.574 0 -3.0 1e-06 
0.05 4.575 0 -3.0 1e-06 
3.0 4.575 0 -3.0 1e-06 
0.05 4.576 0 -3.0 1e-06 
3.0 4.576 0 -3.0 1e-06 
0.05 4.577 0 -3.0 1e-06 
3.0 4.577 0 -3.0 1e-06 
0.05 4.578 0 -3.0 1e-06 
3.0 4.578 0 -3.0 1e-06 
0.05 4.579 0 -3.0 1e-06 
3.0 4.579 0 -3.0 1e-06 
0.05 4.58 0 -3.0 1e-06 
3.0 4.58 0 -3.0 1e-06 
0.05 4.581 0 -3.0 1e-06 
3.0 4.581 0 -3.0 1e-06 
0.05 4.582 0 -3.0 1e-06 
3.0 4.582 0 -3.0 1e-06 
0.05 4.583 0 -3.0 1e-06 
3.0 4.583 0 -3.0 1e-06 
0.05 4.584 0 -3.0 1e-06 
3.0 4.584 0 -3.0 1e-06 
0.05 4.585 0 -3.0 1e-06 
3.0 4.585 0 -3.0 1e-06 
0.05 4.586 0 -3.0 1e-06 
3.0 4.586 0 -3.0 1e-06 
0.05 4.587 0 -3.0 1e-06 
3.0 4.587 0 -3.0 1e-06 
0.05 4.588 0 -3.0 1e-06 
3.0 4.588 0 -3.0 1e-06 
0.05 4.589 0 -3.0 1e-06 
3.0 4.589 0 -3.0 1e-06 
0.05 4.59 0 -3.0 1e-06 
3.0 4.59 0 -3.0 1e-06 
0.05 4.591 0 -3.0 1e-06 
3.0 4.591 0 -3.0 1e-06 
0.05 4.592 0 -3.0 1e-06 
3.0 4.592 0 -3.0 1e-06 
0.05 4.593 0 -3.0 1e-06 
3.0 4.593 0 -3.0 1e-06 
0.05 4.594 0 -3.0 1e-06 
3.0 4.594 0 -3.0 1e-06 
0.05 4.595 0 -3.0 1e-06 
3.0 4.595 0 -3.0 1e-06 
0.05 4.596 0 -3.0 1e-06 
3.0 4.596 0 -3.0 1e-06 
0.05 4.597 0 -3.0 1e-06 
3.0 4.597 0 -3.0 1e-06 
0.05 4.598 0 -3.0 1e-06 
3.0 4.598 0 -3.0 1e-06 
0.05 4.599 0 -3.0 1e-06 
3.0 4.599 0 -3.0 1e-06 
0.05 4.6 0 -3.0 1e-06 
3.0 4.6 0 -3.0 1e-06 
0.05 4.601 0 -3.0 1e-06 
3.0 4.601 0 -3.0 1e-06 
0.05 4.602 0 -3.0 1e-06 
3.0 4.602 0 -3.0 1e-06 
0.05 4.603 0 -3.0 1e-06 
3.0 4.603 0 -3.0 1e-06 
0.05 4.604 0 -3.0 1e-06 
3.0 4.604 0 -3.0 1e-06 
0.05 4.605 0 -3.0 1e-06 
3.0 4.605 0 -3.0 1e-06 
0.05 4.606 0 -3.0 1e-06 
3.0 4.606 0 -3.0 1e-06 
0.05 4.607 0 -3.0 1e-06 
3.0 4.607 0 -3.0 1e-06 
0.05 4.608 0 -3.0 1e-06 
3.0 4.608 0 -3.0 1e-06 
0.05 4.609 0 -3.0 1e-06 
3.0 4.609 0 -3.0 1e-06 
0.05 4.61 0 -3.0 1e-06 
3.0 4.61 0 -3.0 1e-06 
0.05 4.611 0 -3.0 1e-06 
3.0 4.611 0 -3.0 1e-06 
0.05 4.612 0 -3.0 1e-06 
3.0 4.612 0 -3.0 1e-06 
0.05 4.613 0 -3.0 1e-06 
3.0 4.613 0 -3.0 1e-06 
0.05 4.614 0 -3.0 1e-06 
3.0 4.614 0 -3.0 1e-06 
0.05 4.615 0 -3.0 1e-06 
3.0 4.615 0 -3.0 1e-06 
0.05 4.616 0 -3.0 1e-06 
3.0 4.616 0 -3.0 1e-06 
0.05 4.617 0 -3.0 1e-06 
3.0 4.617 0 -3.0 1e-06 
0.05 4.618 0 -3.0 1e-06 
3.0 4.618 0 -3.0 1e-06 
0.05 4.619 0 -3.0 1e-06 
3.0 4.619 0 -3.0 1e-06 
0.05 4.62 0 -3.0 1e-06 
3.0 4.62 0 -3.0 1e-06 
0.05 4.621 0 -3.0 1e-06 
3.0 4.621 0 -3.0 1e-06 
0.05 4.622 0 -3.0 1e-06 
3.0 4.622 0 -3.0 1e-06 
0.05 4.623 0 -3.0 1e-06 
3.0 4.623 0 -3.0 1e-06 
0.05 4.624 0 -3.0 1e-06 
3.0 4.624 0 -3.0 1e-06 
0.05 4.625 0 -3.0 1e-06 
3.0 4.625 0 -3.0 1e-06 
0.05 4.626 0 -3.0 1e-06 
3.0 4.626 0 -3.0 1e-06 
0.05 4.627 0 -3.0 1e-06 
3.0 4.627 0 -3.0 1e-06 
0.05 4.628 0 -3.0 1e-06 
3.0 4.628 0 -3.0 1e-06 
0.05 4.629 0 -3.0 1e-06 
3.0 4.629 0 -3.0 1e-06 
0.05 4.63 0 -3.0 1e-06 
3.0 4.63 0 -3.0 1e-06 
0.05 4.631 0 -3.0 1e-06 
3.0 4.631 0 -3.0 1e-06 
0.05 4.632 0 -3.0 1e-06 
3.0 4.632 0 -3.0 1e-06 
0.05 4.633 0 -3.0 1e-06 
3.0 4.633 0 -3.0 1e-06 
0.05 4.634 0 -3.0 1e-06 
3.0 4.634 0 -3.0 1e-06 
0.05 4.635 0 -3.0 1e-06 
3.0 4.635 0 -3.0 1e-06 
0.05 4.636 0 -3.0 1e-06 
3.0 4.636 0 -3.0 1e-06 
0.05 4.637 0 -3.0 1e-06 
3.0 4.637 0 -3.0 1e-06 
0.05 4.638 0 -3.0 1e-06 
3.0 4.638 0 -3.0 1e-06 
0.05 4.639 0 -3.0 1e-06 
3.0 4.639 0 -3.0 1e-06 
0.05 4.64 0 -3.0 1e-06 
3.0 4.64 0 -3.0 1e-06 
0.05 4.641 0 -3.0 1e-06 
3.0 4.641 0 -3.0 1e-06 
0.05 4.642 0 -3.0 1e-06 
3.0 4.642 0 -3.0 1e-06 
0.05 4.643 0 -3.0 1e-06 
3.0 4.643 0 -3.0 1e-06 
0.05 4.644 0 -3.0 1e-06 
3.0 4.644 0 -3.0 1e-06 
0.05 4.645 0 -3.0 1e-06 
3.0 4.645 0 -3.0 1e-06 
0.05 4.646 0 -3.0 1e-06 
3.0 4.646 0 -3.0 1e-06 
0.05 4.647 0 -3.0 1e-06 
3.0 4.647 0 -3.0 1e-06 
0.05 4.648 0 -3.0 1e-06 
3.0 4.648 0 -3.0 1e-06 
0.05 4.649 0 -3.0 1e-06 
3.0 4.649 0 -3.0 1e-06 
0.05 4.65 0 -3.0 1e-06 
3.0 4.65 0 -3.0 1e-06 
0.05 4.651 0 -3.0 1e-06 
3.0 4.651 0 -3.0 1e-06 
0.05 4.652 0 -3.0 1e-06 
3.0 4.652 0 -3.0 1e-06 
0.05 4.653 0 -3.0 1e-06 
3.0 4.653 0 -3.0 1e-06 
0.05 4.654 0 -3.0 1e-06 
3.0 4.654 0 -3.0 1e-06 
0.05 4.655 0 -3.0 1e-06 
3.0 4.655 0 -3.0 1e-06 
0.05 4.656 0 -3.0 1e-06 
3.0 4.656 0 -3.0 1e-06 
0.05 4.657 0 -3.0 1e-06 
3.0 4.657 0 -3.0 1e-06 
0.05 4.658 0 -3.0 1e-06 
3.0 4.658 0 -3.0 1e-06 
0.05 4.659 0 -3.0 1e-06 
3.0 4.659 0 -3.0 1e-06 
0.05 4.66 0 -3.0 1e-06 
3.0 4.66 0 -3.0 1e-06 
0.05 4.661 0 -3.0 1e-06 
3.0 4.661 0 -3.0 1e-06 
0.05 4.662 0 -3.0 1e-06 
3.0 4.662 0 -3.0 1e-06 
0.05 4.663 0 -3.0 1e-06 
3.0 4.663 0 -3.0 1e-06 
0.05 4.664 0 -3.0 1e-06 
3.0 4.664 0 -3.0 1e-06 
0.05 4.665 0 -3.0 1e-06 
3.0 4.665 0 -3.0 1e-06 
0.05 4.666 0 -3.0 1e-06 
3.0 4.666 0 -3.0 1e-06 
0.05 4.667 0 -3.0 1e-06 
3.0 4.667 0 -3.0 1e-06 
0.05 4.668 0 -3.0 1e-06 
3.0 4.668 0 -3.0 1e-06 
0.05 4.669 0 -3.0 1e-06 
3.0 4.669 0 -3.0 1e-06 
0.05 4.67 0 -3.0 1e-06 
3.0 4.67 0 -3.0 1e-06 
0.05 4.671 0 -3.0 1e-06 
3.0 4.671 0 -3.0 1e-06 
0.05 4.672 0 -3.0 1e-06 
3.0 4.672 0 -3.0 1e-06 
0.05 4.673 0 -3.0 1e-06 
3.0 4.673 0 -3.0 1e-06 
0.05 4.674 0 -3.0 1e-06 
3.0 4.674 0 -3.0 1e-06 
0.05 4.675 0 -3.0 1e-06 
3.0 4.675 0 -3.0 1e-06 
0.05 4.676 0 -3.0 1e-06 
3.0 4.676 0 -3.0 1e-06 
0.05 4.677 0 -3.0 1e-06 
3.0 4.677 0 -3.0 1e-06 
0.05 4.678 0 -3.0 1e-06 
3.0 4.678 0 -3.0 1e-06 
0.05 4.679 0 -3.0 1e-06 
3.0 4.679 0 -3.0 1e-06 
0.05 4.68 0 -3.0 1e-06 
3.0 4.68 0 -3.0 1e-06 
0.05 4.681 0 -3.0 1e-06 
3.0 4.681 0 -3.0 1e-06 
0.05 4.682 0 -3.0 1e-06 
3.0 4.682 0 -3.0 1e-06 
0.05 4.683 0 -3.0 1e-06 
3.0 4.683 0 -3.0 1e-06 
0.05 4.684 0 -3.0 1e-06 
3.0 4.684 0 -3.0 1e-06 
0.05 4.685 0 -3.0 1e-06 
3.0 4.685 0 -3.0 1e-06 
0.05 4.686 0 -3.0 1e-06 
3.0 4.686 0 -3.0 1e-06 
0.05 4.687 0 -3.0 1e-06 
3.0 4.687 0 -3.0 1e-06 
0.05 4.688 0 -3.0 1e-06 
3.0 4.688 0 -3.0 1e-06 
0.05 4.689 0 -3.0 1e-06 
3.0 4.689 0 -3.0 1e-06 
0.05 4.69 0 -3.0 1e-06 
3.0 4.69 0 -3.0 1e-06 
0.05 4.691 0 -3.0 1e-06 
3.0 4.691 0 -3.0 1e-06 
0.05 4.692 0 -3.0 1e-06 
3.0 4.692 0 -3.0 1e-06 
0.05 4.693 0 -3.0 1e-06 
3.0 4.693 0 -3.0 1e-06 
0.05 4.694 0 -3.0 1e-06 
3.0 4.694 0 -3.0 1e-06 
0.05 4.695 0 -3.0 1e-06 
3.0 4.695 0 -3.0 1e-06 
0.05 4.696 0 -3.0 1e-06 
3.0 4.696 0 -3.0 1e-06 
0.05 4.697 0 -3.0 1e-06 
3.0 4.697 0 -3.0 1e-06 
0.05 4.698 0 -3.0 1e-06 
3.0 4.698 0 -3.0 1e-06 
0.05 4.699 0 -3.0 1e-06 
3.0 4.699 0 -3.0 1e-06 
0.05 4.7 0 -3.0 1e-06 
3.0 4.7 0 -3.0 1e-06 
0.05 4.701 0 -3.0 1e-06 
3.0 4.701 0 -3.0 1e-06 
0.05 4.702 0 -3.0 1e-06 
3.0 4.702 0 -3.0 1e-06 
0.05 4.703 0 -3.0 1e-06 
3.0 4.703 0 -3.0 1e-06 
0.05 4.704 0 -3.0 1e-06 
3.0 4.704 0 -3.0 1e-06 
0.05 4.705 0 -3.0 1e-06 
3.0 4.705 0 -3.0 1e-06 
0.05 4.706 0 -3.0 1e-06 
3.0 4.706 0 -3.0 1e-06 
0.05 4.707 0 -3.0 1e-06 
3.0 4.707 0 -3.0 1e-06 
0.05 4.708 0 -3.0 1e-06 
3.0 4.708 0 -3.0 1e-06 
0.05 4.709 0 -3.0 1e-06 
3.0 4.709 0 -3.0 1e-06 
0.05 4.71 0 -3.0 1e-06 
3.0 4.71 0 -3.0 1e-06 
0.05 4.711 0 -3.0 1e-06 
3.0 4.711 0 -3.0 1e-06 
0.05 4.712 0 -3.0 1e-06 
3.0 4.712 0 -3.0 1e-06 
0.05 4.713 0 -3.0 1e-06 
3.0 4.713 0 -3.0 1e-06 
0.05 4.714 0 -3.0 1e-06 
3.0 4.714 0 -3.0 1e-06 
0.05 4.715 0 -3.0 1e-06 
3.0 4.715 0 -3.0 1e-06 
0.05 4.716 0 -3.0 1e-06 
3.0 4.716 0 -3.0 1e-06 
0.05 4.717 0 -3.0 1e-06 
3.0 4.717 0 -3.0 1e-06 
0.05 4.718 0 -3.0 1e-06 
3.0 4.718 0 -3.0 1e-06 
0.05 4.719 0 -3.0 1e-06 
3.0 4.719 0 -3.0 1e-06 
0.05 4.72 0 -3.0 1e-06 
3.0 4.72 0 -3.0 1e-06 
0.05 4.721 0 -3.0 1e-06 
3.0 4.721 0 -3.0 1e-06 
0.05 4.722 0 -3.0 1e-06 
3.0 4.722 0 -3.0 1e-06 
0.05 4.723 0 -3.0 1e-06 
3.0 4.723 0 -3.0 1e-06 
0.05 4.724 0 -3.0 1e-06 
3.0 4.724 0 -3.0 1e-06 
0.05 4.725 0 -3.0 1e-06 
3.0 4.725 0 -3.0 1e-06 
0.05 4.726 0 -3.0 1e-06 
3.0 4.726 0 -3.0 1e-06 
0.05 4.727 0 -3.0 1e-06 
3.0 4.727 0 -3.0 1e-06 
0.05 4.728 0 -3.0 1e-06 
3.0 4.728 0 -3.0 1e-06 
0.05 4.729 0 -3.0 1e-06 
3.0 4.729 0 -3.0 1e-06 
0.05 4.73 0 -3.0 1e-06 
3.0 4.73 0 -3.0 1e-06 
0.05 4.731 0 -3.0 1e-06 
3.0 4.731 0 -3.0 1e-06 
0.05 4.732 0 -3.0 1e-06 
3.0 4.732 0 -3.0 1e-06 
0.05 4.733 0 -3.0 1e-06 
3.0 4.733 0 -3.0 1e-06 
0.05 4.734 0 -3.0 1e-06 
3.0 4.734 0 -3.0 1e-06 
0.05 4.735 0 -3.0 1e-06 
3.0 4.735 0 -3.0 1e-06 
0.05 4.736 0 -3.0 1e-06 
3.0 4.736 0 -3.0 1e-06 
0.05 4.737 0 -3.0 1e-06 
3.0 4.737 0 -3.0 1e-06 
0.05 4.738 0 -3.0 1e-06 
3.0 4.738 0 -3.0 1e-06 
0.05 4.739 0 -3.0 1e-06 
3.0 4.739 0 -3.0 1e-06 
0.05 4.74 0 -3.0 1e-06 
3.0 4.74 0 -3.0 1e-06 
0.05 4.741 0 -3.0 1e-06 
3.0 4.741 0 -3.0 1e-06 
0.05 4.742 0 -3.0 1e-06 
3.0 4.742 0 -3.0 1e-06 
0.05 4.743 0 -3.0 1e-06 
3.0 4.743 0 -3.0 1e-06 
0.05 4.744 0 -3.0 1e-06 
3.0 4.744 0 -3.0 1e-06 
0.05 4.745 0 -3.0 1e-06 
3.0 4.745 0 -3.0 1e-06 
0.05 4.746 0 -3.0 1e-06 
3.0 4.746 0 -3.0 1e-06 
0.05 4.747 0 -3.0 1e-06 
3.0 4.747 0 -3.0 1e-06 
0.05 4.748 0 -3.0 1e-06 
3.0 4.748 0 -3.0 1e-06 
0.05 4.749 0 -3.0 1e-06 
3.0 4.749 0 -3.0 1e-06 
0.05 4.75 0 -3.0 1e-06 
3.0 4.75 0 -3.0 1e-06 
0.05 4.751 0 -3.0 1e-06 
3.0 4.751 0 -3.0 1e-06 
0.05 4.752 0 -3.0 1e-06 
3.0 4.752 0 -3.0 1e-06 
0.05 4.753 0 -3.0 1e-06 
3.0 4.753 0 -3.0 1e-06 
0.05 4.754 0 -3.0 1e-06 
3.0 4.754 0 -3.0 1e-06 
0.05 4.755 0 -3.0 1e-06 
3.0 4.755 0 -3.0 1e-06 
0.05 4.756 0 -3.0 1e-06 
3.0 4.756 0 -3.0 1e-06 
0.05 4.757 0 -3.0 1e-06 
3.0 4.757 0 -3.0 1e-06 
0.05 4.758 0 -3.0 1e-06 
3.0 4.758 0 -3.0 1e-06 
0.05 4.759 0 -3.0 1e-06 
3.0 4.759 0 -3.0 1e-06 
0.05 4.76 0 -3.0 1e-06 
3.0 4.76 0 -3.0 1e-06 
0.05 4.761 0 -3.0 1e-06 
3.0 4.761 0 -3.0 1e-06 
0.05 4.762 0 -3.0 1e-06 
3.0 4.762 0 -3.0 1e-06 
0.05 4.763 0 -3.0 1e-06 
3.0 4.763 0 -3.0 1e-06 
0.05 4.764 0 -3.0 1e-06 
3.0 4.764 0 -3.0 1e-06 
0.05 4.765 0 -3.0 1e-06 
3.0 4.765 0 -3.0 1e-06 
0.05 4.766 0 -3.0 1e-06 
3.0 4.766 0 -3.0 1e-06 
0.05 4.767 0 -3.0 1e-06 
3.0 4.767 0 -3.0 1e-06 
0.05 4.768 0 -3.0 1e-06 
3.0 4.768 0 -3.0 1e-06 
0.05 4.769 0 -3.0 1e-06 
3.0 4.769 0 -3.0 1e-06 
0.05 4.77 0 -3.0 1e-06 
3.0 4.77 0 -3.0 1e-06 
0.05 4.771 0 -3.0 1e-06 
3.0 4.771 0 -3.0 1e-06 
0.05 4.772 0 -3.0 1e-06 
3.0 4.772 0 -3.0 1e-06 
0.05 4.773 0 -3.0 1e-06 
3.0 4.773 0 -3.0 1e-06 
0.05 4.774 0 -3.0 1e-06 
3.0 4.774 0 -3.0 1e-06 
0.05 4.775 0 -3.0 1e-06 
3.0 4.775 0 -3.0 1e-06 
0.05 4.776 0 -3.0 1e-06 
3.0 4.776 0 -3.0 1e-06 
0.05 4.777 0 -3.0 1e-06 
3.0 4.777 0 -3.0 1e-06 
0.05 4.778 0 -3.0 1e-06 
3.0 4.778 0 -3.0 1e-06 
0.05 4.779 0 -3.0 1e-06 
3.0 4.779 0 -3.0 1e-06 
0.05 4.78 0 -3.0 1e-06 
3.0 4.78 0 -3.0 1e-06 
0.05 4.781 0 -3.0 1e-06 
3.0 4.781 0 -3.0 1e-06 
0.05 4.782 0 -3.0 1e-06 
3.0 4.782 0 -3.0 1e-06 
0.05 4.783 0 -3.0 1e-06 
3.0 4.783 0 -3.0 1e-06 
0.05 4.784 0 -3.0 1e-06 
3.0 4.784 0 -3.0 1e-06 
0.05 4.785 0 -3.0 1e-06 
3.0 4.785 0 -3.0 1e-06 
0.05 4.786 0 -3.0 1e-06 
3.0 4.786 0 -3.0 1e-06 
0.05 4.787 0 -3.0 1e-06 
3.0 4.787 0 -3.0 1e-06 
0.05 4.788 0 -3.0 1e-06 
3.0 4.788 0 -3.0 1e-06 
0.05 4.789 0 -3.0 1e-06 
3.0 4.789 0 -3.0 1e-06 
0.05 4.79 0 -3.0 1e-06 
3.0 4.79 0 -3.0 1e-06 
0.05 4.791 0 -3.0 1e-06 
3.0 4.791 0 -3.0 1e-06 
0.05 4.792 0 -3.0 1e-06 
3.0 4.792 0 -3.0 1e-06 
0.05 4.793 0 -3.0 1e-06 
3.0 4.793 0 -3.0 1e-06 
0.05 4.794 0 -3.0 1e-06 
3.0 4.794 0 -3.0 1e-06 
0.05 4.795 0 -3.0 1e-06 
3.0 4.795 0 -3.0 1e-06 
0.05 4.796 0 -3.0 1e-06 
3.0 4.796 0 -3.0 1e-06 
0.05 4.797 0 -3.0 1e-06 
3.0 4.797 0 -3.0 1e-06 
0.05 4.798 0 -3.0 1e-06 
3.0 4.798 0 -3.0 1e-06 
0.05 4.799 0 -3.0 1e-06 
3.0 4.799 0 -3.0 1e-06 
0.05 4.8 0 -3.0 1e-06 
3.0 4.8 0 -3.0 1e-06 
0.05 4.801 0 -3.0 1e-06 
3.0 4.801 0 -3.0 1e-06 
0.05 4.802 0 -3.0 1e-06 
3.0 4.802 0 -3.0 1e-06 
0.05 4.803 0 -3.0 1e-06 
3.0 4.803 0 -3.0 1e-06 
0.05 4.804 0 -3.0 1e-06 
3.0 4.804 0 -3.0 1e-06 
0.05 4.805 0 -3.0 1e-06 
3.0 4.805 0 -3.0 1e-06 
0.05 4.806 0 -3.0 1e-06 
3.0 4.806 0 -3.0 1e-06 
0.05 4.807 0 -3.0 1e-06 
3.0 4.807 0 -3.0 1e-06 
0.05 4.808 0 -3.0 1e-06 
3.0 4.808 0 -3.0 1e-06 
0.05 4.809 0 -3.0 1e-06 
3.0 4.809 0 -3.0 1e-06 
0.05 4.81 0 -3.0 1e-06 
3.0 4.81 0 -3.0 1e-06 
0.05 4.811 0 -3.0 1e-06 
3.0 4.811 0 -3.0 1e-06 
0.05 4.812 0 -3.0 1e-06 
3.0 4.812 0 -3.0 1e-06 
0.05 4.813 0 -3.0 1e-06 
3.0 4.813 0 -3.0 1e-06 
0.05 4.814 0 -3.0 1e-06 
3.0 4.814 0 -3.0 1e-06 
0.05 4.815 0 -3.0 1e-06 
3.0 4.815 0 -3.0 1e-06 
0.05 4.816 0 -3.0 1e-06 
3.0 4.816 0 -3.0 1e-06 
0.05 4.817 0 -3.0 1e-06 
3.0 4.817 0 -3.0 1e-06 
0.05 4.818 0 -3.0 1e-06 
3.0 4.818 0 -3.0 1e-06 
0.05 4.819 0 -3.0 1e-06 
3.0 4.819 0 -3.0 1e-06 
0.05 4.82 0 -3.0 1e-06 
3.0 4.82 0 -3.0 1e-06 
0.05 4.821 0 -3.0 1e-06 
3.0 4.821 0 -3.0 1e-06 
0.05 4.822 0 -3.0 1e-06 
3.0 4.822 0 -3.0 1e-06 
0.05 4.823 0 -3.0 1e-06 
3.0 4.823 0 -3.0 1e-06 
0.05 4.824 0 -3.0 1e-06 
3.0 4.824 0 -3.0 1e-06 
0.05 4.825 0 -3.0 1e-06 
3.0 4.825 0 -3.0 1e-06 
0.05 4.826 0 -3.0 1e-06 
3.0 4.826 0 -3.0 1e-06 
0.05 4.827 0 -3.0 1e-06 
3.0 4.827 0 -3.0 1e-06 
0.05 4.828 0 -3.0 1e-06 
3.0 4.828 0 -3.0 1e-06 
0.05 4.829 0 -3.0 1e-06 
3.0 4.829 0 -3.0 1e-06 
0.05 4.83 0 -3.0 1e-06 
3.0 4.83 0 -3.0 1e-06 
0.05 4.831 0 -3.0 1e-06 
3.0 4.831 0 -3.0 1e-06 
0.05 4.832 0 -3.0 1e-06 
3.0 4.832 0 -3.0 1e-06 
0.05 4.833 0 -3.0 1e-06 
3.0 4.833 0 -3.0 1e-06 
0.05 4.834 0 -3.0 1e-06 
3.0 4.834 0 -3.0 1e-06 
0.05 4.835 0 -3.0 1e-06 
3.0 4.835 0 -3.0 1e-06 
0.05 4.836 0 -3.0 1e-06 
3.0 4.836 0 -3.0 1e-06 
0.05 4.837 0 -3.0 1e-06 
3.0 4.837 0 -3.0 1e-06 
0.05 4.838 0 -3.0 1e-06 
3.0 4.838 0 -3.0 1e-06 
0.05 4.839 0 -3.0 1e-06 
3.0 4.839 0 -3.0 1e-06 
0.05 4.84 0 -3.0 1e-06 
3.0 4.84 0 -3.0 1e-06 
0.05 4.841 0 -3.0 1e-06 
3.0 4.841 0 -3.0 1e-06 
0.05 4.842 0 -3.0 1e-06 
3.0 4.842 0 -3.0 1e-06 
0.05 4.843 0 -3.0 1e-06 
3.0 4.843 0 -3.0 1e-06 
0.05 4.844 0 -3.0 1e-06 
3.0 4.844 0 -3.0 1e-06 
0.05 4.845 0 -3.0 1e-06 
3.0 4.845 0 -3.0 1e-06 
0.05 4.846 0 -3.0 1e-06 
3.0 4.846 0 -3.0 1e-06 
0.05 4.847 0 -3.0 1e-06 
3.0 4.847 0 -3.0 1e-06 
0.05 4.848 0 -3.0 1e-06 
3.0 4.848 0 -3.0 1e-06 
0.05 4.849 0 -3.0 1e-06 
3.0 4.849 0 -3.0 1e-06 
0.05 4.85 0 -3.0 1e-06 
3.0 4.85 0 -3.0 1e-06 
0.05 4.851 0 -3.0 1e-06 
3.0 4.851 0 -3.0 1e-06 
0.05 4.852 0 -3.0 1e-06 
3.0 4.852 0 -3.0 1e-06 
0.05 4.853 0 -3.0 1e-06 
3.0 4.853 0 -3.0 1e-06 
0.05 4.854 0 -3.0 1e-06 
3.0 4.854 0 -3.0 1e-06 
0.05 4.855 0 -3.0 1e-06 
3.0 4.855 0 -3.0 1e-06 
0.05 4.856 0 -3.0 1e-06 
3.0 4.856 0 -3.0 1e-06 
0.05 4.857 0 -3.0 1e-06 
3.0 4.857 0 -3.0 1e-06 
0.05 4.858 0 -3.0 1e-06 
3.0 4.858 0 -3.0 1e-06 
0.05 4.859 0 -3.0 1e-06 
3.0 4.859 0 -3.0 1e-06 
0.05 4.86 0 -3.0 1e-06 
3.0 4.86 0 -3.0 1e-06 
0.05 4.861 0 -3.0 1e-06 
3.0 4.861 0 -3.0 1e-06 
0.05 4.862 0 -3.0 1e-06 
3.0 4.862 0 -3.0 1e-06 
0.05 4.863 0 -3.0 1e-06 
3.0 4.863 0 -3.0 1e-06 
0.05 4.864 0 -3.0 1e-06 
3.0 4.864 0 -3.0 1e-06 
0.05 4.865 0 -3.0 1e-06 
3.0 4.865 0 -3.0 1e-06 
0.05 4.866 0 -3.0 1e-06 
3.0 4.866 0 -3.0 1e-06 
0.05 4.867 0 -3.0 1e-06 
3.0 4.867 0 -3.0 1e-06 
0.05 4.868 0 -3.0 1e-06 
3.0 4.868 0 -3.0 1e-06 
0.05 4.869 0 -3.0 1e-06 
3.0 4.869 0 -3.0 1e-06 
0.05 4.87 0 -3.0 1e-06 
3.0 4.87 0 -3.0 1e-06 
0.05 4.871 0 -3.0 1e-06 
3.0 4.871 0 -3.0 1e-06 
0.05 4.872 0 -3.0 1e-06 
3.0 4.872 0 -3.0 1e-06 
0.05 4.873 0 -3.0 1e-06 
3.0 4.873 0 -3.0 1e-06 
0.05 4.874 0 -3.0 1e-06 
3.0 4.874 0 -3.0 1e-06 
0.05 4.875 0 -3.0 1e-06 
3.0 4.875 0 -3.0 1e-06 
0.05 4.876 0 -3.0 1e-06 
3.0 4.876 0 -3.0 1e-06 
0.05 4.877 0 -3.0 1e-06 
3.0 4.877 0 -3.0 1e-06 
0.05 4.878 0 -3.0 1e-06 
3.0 4.878 0 -3.0 1e-06 
0.05 4.879 0 -3.0 1e-06 
3.0 4.879 0 -3.0 1e-06 
0.05 4.88 0 -3.0 1e-06 
3.0 4.88 0 -3.0 1e-06 
0.05 4.881 0 -3.0 1e-06 
3.0 4.881 0 -3.0 1e-06 
0.05 4.882 0 -3.0 1e-06 
3.0 4.882 0 -3.0 1e-06 
0.05 4.883 0 -3.0 1e-06 
3.0 4.883 0 -3.0 1e-06 
0.05 4.884 0 -3.0 1e-06 
3.0 4.884 0 -3.0 1e-06 
0.05 4.885 0 -3.0 1e-06 
3.0 4.885 0 -3.0 1e-06 
0.05 4.886 0 -3.0 1e-06 
3.0 4.886 0 -3.0 1e-06 
0.05 4.887 0 -3.0 1e-06 
3.0 4.887 0 -3.0 1e-06 
0.05 4.888 0 -3.0 1e-06 
3.0 4.888 0 -3.0 1e-06 
0.05 4.889 0 -3.0 1e-06 
3.0 4.889 0 -3.0 1e-06 
0.05 4.89 0 -3.0 1e-06 
3.0 4.89 0 -3.0 1e-06 
0.05 4.891 0 -3.0 1e-06 
3.0 4.891 0 -3.0 1e-06 
0.05 4.892 0 -3.0 1e-06 
3.0 4.892 0 -3.0 1e-06 
0.05 4.893 0 -3.0 1e-06 
3.0 4.893 0 -3.0 1e-06 
0.05 4.894 0 -3.0 1e-06 
3.0 4.894 0 -3.0 1e-06 
0.05 4.895 0 -3.0 1e-06 
3.0 4.895 0 -3.0 1e-06 
0.05 4.896 0 -3.0 1e-06 
3.0 4.896 0 -3.0 1e-06 
0.05 4.897 0 -3.0 1e-06 
3.0 4.897 0 -3.0 1e-06 
0.05 4.898 0 -3.0 1e-06 
3.0 4.898 0 -3.0 1e-06 
0.05 4.899 0 -3.0 1e-06 
3.0 4.899 0 -3.0 1e-06 
0.05 4.9 0 -3.0 1e-06 
3.0 4.9 0 -3.0 1e-06 
0.05 4.901 0 -3.0 1e-06 
3.0 4.901 0 -3.0 1e-06 
0.05 4.902 0 -3.0 1e-06 
3.0 4.902 0 -3.0 1e-06 
0.05 4.903 0 -3.0 1e-06 
3.0 4.903 0 -3.0 1e-06 
0.05 4.904 0 -3.0 1e-06 
3.0 4.904 0 -3.0 1e-06 
0.05 4.905 0 -3.0 1e-06 
3.0 4.905 0 -3.0 1e-06 
0.05 4.906 0 -3.0 1e-06 
3.0 4.906 0 -3.0 1e-06 
0.05 4.907 0 -3.0 1e-06 
3.0 4.907 0 -3.0 1e-06 
0.05 4.908 0 -3.0 1e-06 
3.0 4.908 0 -3.0 1e-06 
0.05 4.909 0 -3.0 1e-06 
3.0 4.909 0 -3.0 1e-06 
0.05 4.91 0 -3.0 1e-06 
3.0 4.91 0 -3.0 1e-06 
0.05 4.911 0 -3.0 1e-06 
3.0 4.911 0 -3.0 1e-06 
0.05 4.912 0 -3.0 1e-06 
3.0 4.912 0 -3.0 1e-06 
0.05 4.913 0 -3.0 1e-06 
3.0 4.913 0 -3.0 1e-06 
0.05 4.914 0 -3.0 1e-06 
3.0 4.914 0 -3.0 1e-06 
0.05 4.915 0 -3.0 1e-06 
3.0 4.915 0 -3.0 1e-06 
0.05 4.916 0 -3.0 1e-06 
3.0 4.916 0 -3.0 1e-06 
0.05 4.917 0 -3.0 1e-06 
3.0 4.917 0 -3.0 1e-06 
0.05 4.918 0 -3.0 1e-06 
3.0 4.918 0 -3.0 1e-06 
0.05 4.919 0 -3.0 1e-06 
3.0 4.919 0 -3.0 1e-06 
0.05 4.92 0 -3.0 1e-06 
3.0 4.92 0 -3.0 1e-06 
0.05 4.921 0 -3.0 1e-06 
3.0 4.921 0 -3.0 1e-06 
0.05 4.922 0 -3.0 1e-06 
3.0 4.922 0 -3.0 1e-06 
0.05 4.923 0 -3.0 1e-06 
3.0 4.923 0 -3.0 1e-06 
0.05 4.924 0 -3.0 1e-06 
3.0 4.924 0 -3.0 1e-06 
0.05 4.925 0 -3.0 1e-06 
3.0 4.925 0 -3.0 1e-06 
0.05 4.926 0 -3.0 1e-06 
3.0 4.926 0 -3.0 1e-06 
0.05 4.927 0 -3.0 1e-06 
3.0 4.927 0 -3.0 1e-06 
0.05 4.928 0 -3.0 1e-06 
3.0 4.928 0 -3.0 1e-06 
0.05 4.929 0 -3.0 1e-06 
3.0 4.929 0 -3.0 1e-06 
0.05 4.93 0 -3.0 1e-06 
3.0 4.93 0 -3.0 1e-06 
0.05 4.931 0 -3.0 1e-06 
3.0 4.931 0 -3.0 1e-06 
0.05 4.932 0 -3.0 1e-06 
3.0 4.932 0 -3.0 1e-06 
0.05 4.933 0 -3.0 1e-06 
3.0 4.933 0 -3.0 1e-06 
0.05 4.934 0 -3.0 1e-06 
3.0 4.934 0 -3.0 1e-06 
0.05 4.935 0 -3.0 1e-06 
3.0 4.935 0 -3.0 1e-06 
0.05 4.936 0 -3.0 1e-06 
3.0 4.936 0 -3.0 1e-06 
0.05 4.937 0 -3.0 1e-06 
3.0 4.937 0 -3.0 1e-06 
0.05 4.938 0 -3.0 1e-06 
3.0 4.938 0 -3.0 1e-06 
0.05 4.939 0 -3.0 1e-06 
3.0 4.939 0 -3.0 1e-06 
0.05 4.94 0 -3.0 1e-06 
3.0 4.94 0 -3.0 1e-06 
0.05 4.941 0 -3.0 1e-06 
3.0 4.941 0 -3.0 1e-06 
0.05 4.942 0 -3.0 1e-06 
3.0 4.942 0 -3.0 1e-06 
0.05 4.943 0 -3.0 1e-06 
3.0 4.943 0 -3.0 1e-06 
0.05 4.944 0 -3.0 1e-06 
3.0 4.944 0 -3.0 1e-06 
0.05 4.945 0 -3.0 1e-06 
3.0 4.945 0 -3.0 1e-06 
0.05 4.946 0 -3.0 1e-06 
3.0 4.946 0 -3.0 1e-06 
0.05 4.947 0 -3.0 1e-06 
3.0 4.947 0 -3.0 1e-06 
0.05 4.948 0 -3.0 1e-06 
3.0 4.948 0 -3.0 1e-06 
0.05 4.949 0 -3.0 1e-06 
3.0 4.949 0 -3.0 1e-06 
0.05 4.95 0 -3.0 1e-06 
3.0 4.95 0 -3.0 1e-06 
0.05 4.951 0 -3.0 1e-06 
3.0 4.951 0 -3.0 1e-06 
0.05 4.952 0 -3.0 1e-06 
3.0 4.952 0 -3.0 1e-06 
0.05 4.953 0 -3.0 1e-06 
3.0 4.953 0 -3.0 1e-06 
0.05 4.954 0 -3.0 1e-06 
3.0 4.954 0 -3.0 1e-06 
0.05 4.955 0 -3.0 1e-06 
3.0 4.955 0 -3.0 1e-06 
0.05 4.956 0 -3.0 1e-06 
3.0 4.956 0 -3.0 1e-06 
0.05 4.957 0 -3.0 1e-06 
3.0 4.957 0 -3.0 1e-06 
0.05 4.958 0 -3.0 1e-06 
3.0 4.958 0 -3.0 1e-06 
0.05 4.959 0 -3.0 1e-06 
3.0 4.959 0 -3.0 1e-06 
0.05 4.96 0 -3.0 1e-06 
3.0 4.96 0 -3.0 1e-06 
0.05 4.961 0 -3.0 1e-06 
3.0 4.961 0 -3.0 1e-06 
0.05 4.962 0 -3.0 1e-06 
3.0 4.962 0 -3.0 1e-06 
0.05 4.963 0 -3.0 1e-06 
3.0 4.963 0 -3.0 1e-06 
0.05 4.964 0 -3.0 1e-06 
3.0 4.964 0 -3.0 1e-06 
0.05 4.965 0 -3.0 1e-06 
3.0 4.965 0 -3.0 1e-06 
0.05 4.966 0 -3.0 1e-06 
3.0 4.966 0 -3.0 1e-06 
0.05 4.967 0 -3.0 1e-06 
3.0 4.967 0 -3.0 1e-06 
0.05 4.968 0 -3.0 1e-06 
3.0 4.968 0 -3.0 1e-06 
0.05 4.969 0 -3.0 1e-06 
3.0 4.969 0 -3.0 1e-06 
0.05 4.97 0 -3.0 1e-06 
3.0 4.97 0 -3.0 1e-06 
0.05 4.971 0 -3.0 1e-06 
3.0 4.971 0 -3.0 1e-06 
0.05 4.972 0 -3.0 1e-06 
3.0 4.972 0 -3.0 1e-06 
0.05 4.973 0 -3.0 1e-06 
3.0 4.973 0 -3.0 1e-06 
0.05 4.974 0 -3.0 1e-06 
3.0 4.974 0 -3.0 1e-06 
0.05 4.975 0 -3.0 1e-06 
3.0 4.975 0 -3.0 1e-06 
0.05 4.976 0 -3.0 1e-06 
3.0 4.976 0 -3.0 1e-06 
0.05 4.977 0 -3.0 1e-06 
3.0 4.977 0 -3.0 1e-06 
0.05 4.978 0 -3.0 1e-06 
3.0 4.978 0 -3.0 1e-06 
0.05 4.979 0 -3.0 1e-06 
3.0 4.979 0 -3.0 1e-06 
0.05 4.98 0 -3.0 1e-06 
3.0 4.98 0 -3.0 1e-06 
0.05 4.981 0 -3.0 1e-06 
3.0 4.981 0 -3.0 1e-06 
0.05 4.982 0 -3.0 1e-06 
3.0 4.982 0 -3.0 1e-06 
0.05 4.983 0 -3.0 1e-06 
3.0 4.983 0 -3.0 1e-06 
0.05 4.984 0 -3.0 1e-06 
3.0 4.984 0 -3.0 1e-06 
0.05 4.985 0 -3.0 1e-06 
3.0 4.985 0 -3.0 1e-06 
0.05 4.986 0 -3.0 1e-06 
3.0 4.986 0 -3.0 1e-06 
0.05 4.987 0 -3.0 1e-06 
3.0 4.987 0 -3.0 1e-06 
0.05 4.988 0 -3.0 1e-06 
3.0 4.988 0 -3.0 1e-06 
0.05 4.989 0 -3.0 1e-06 
3.0 4.989 0 -3.0 1e-06 
0.05 4.99 0 -3.0 1e-06 
3.0 4.99 0 -3.0 1e-06 
0.05 4.991 0 -3.0 1e-06 
3.0 4.991 0 -3.0 1e-06 
0.05 4.992 0 -3.0 1e-06 
3.0 4.992 0 -3.0 1e-06 
0.05 4.993 0 -3.0 1e-06 
3.0 4.993 0 -3.0 1e-06 
0.05 4.994 0 -3.0 1e-06 
3.0 4.994 0 -3.0 1e-06 
0.05 4.995 0 -3.0 1e-06 
3.0 4.995 0 -3.0 1e-06 
0.05 4.996 0 -3.0 1e-06 
3.0 4.996 0 -3.0 1e-06 
0.05 4.997 0 -3.0 1e-06 
3.0 4.997 0 -3.0 1e-06 
0.05 4.998 0 -3.0 1e-06 
3.0 4.998 0 -3.0 1e-06 
0.05 4.999 0 -3.0 1e-06 
3.0 4.999 0 -3.0 1e-06 
0.05 0.0 0 0.0 1e-06 
3.0 0.0 0 0.0 1e-06 
0.05 0.001 0 0.0 1e-06 
3.0 0.001 0 0.0 1e-06 
0.05 0.002 0 0.0 1e-06 
3.0 0.002 0 0.0 1e-06 
0.05 0.003 0 0.0 1e-06 
3.0 0.003 0 0.0 1e-06 
0.05 0.004 0 0.0 1e-06 
3.0 0.004 0 0.0 1e-06 
0.05 0.005 0 0.0 1e-06 
3.0 0.005 0 0.0 1e-06 
0.05 0.006 0 0.0 1e-06 
3.0 0.006 0 0.0 1e-06 
0.05 0.007 0 0.0 1e-06 
3.0 0.007 0 0.0 1e-06 
0.05 0.008 0 0.0 1e-06 
3.0 0.008 0 0.0 1e-06 
0.05 0.009 0 0.0 1e-06 
3.0 0.009 0 0.0 1e-06 
0.05 0.01 0 0.0 1e-06 
3.0 0.01 0 0.0 1e-06 
0.05 0.011 0 0.0 1e-06 
3.0 0.011 0 0.0 1e-06 
0.05 0.012 0 0.0 1e-06 
3.0 0.012 0 0.0 1e-06 
0.05 0.013 0 0.0 1e-06 
3.0 0.013 0 0.0 1e-06 
0.05 0.014 0 0.0 1e-06 
3.0 0.014 0 0.0 1e-06 
0.05 0.015 0 0.0 1e-06 
3.0 0.015 0 0.0 1e-06 
0.05 0.016 0 0.0 1e-06 
3.0 0.016 0 0.0 1e-06 
0.05 0.017 0 0.0 1e-06 
3.0 0.017 0 0.0 1e-06 
0.05 0.018 0 0.0 1e-06 
3.0 0.018 0 0.0 1e-06 
0.05 0.019 0 0.0 1e-06 
3.0 0.019 0 0.0 1e-06 
0.05 0.02 0 0.0 1e-06 
3.0 0.02 0 0.0 1e-06 
0.05 0.021 0 0.0 1e-06 
3.0 0.021 0 0.0 1e-06 
0.05 0.022 0 0.0 1e-06 
3.0 0.022 0 0.0 1e-06 
0.05 0.023 0 0.0 1e-06 
3.0 0.023 0 0.0 1e-06 
0.05 0.024 0 0.0 1e-06 
3.0 0.024 0 0.0 1e-06 
0.05 0.025 0 0.0 1e-06 
3.0 0.025 0 0.0 1e-06 
0.05 0.026 0 0.0 1e-06 
3.0 0.026 0 0.0 1e-06 
0.05 0.027 0 0.0 1e-06 
3.0 0.027 0 0.0 1e-06 
0.05 0.028 0 0.0 1e-06 
3.0 0.028 0 0.0 1e-06 
0.05 0.029 0 0.0 1e-06 
3.0 0.029 0 0.0 1e-06 
0.05 0.03 0 0.0 1e-06 
3.0 0.03 0 0.0 1e-06 
0.05 0.031 0 0.0 1e-06 
3.0 0.031 0 0.0 1e-06 
0.05 0.032 0 0.0 1e-06 
3.0 0.032 0 0.0 1e-06 
0.05 0.033 0 0.0 1e-06 
3.0 0.033 0 0.0 1e-06 
0.05 0.034 0 0.0 1e-06 
3.0 0.034 0 0.0 1e-06 
0.05 0.035 0 0.0 1e-06 
3.0 0.035 0 0.0 1e-06 
0.05 0.036 0 0.0 1e-06 
3.0 0.036 0 0.0 1e-06 
0.05 0.037 0 0.0 1e-06 
3.0 0.037 0 0.0 1e-06 
0.05 0.038 0 0.0 1e-06 
3.0 0.038 0 0.0 1e-06 
0.05 0.039 0 0.0 1e-06 
3.0 0.039 0 0.0 1e-06 
0.05 0.04 0 0.0 1e-06 
3.0 0.04 0 0.0 1e-06 
0.05 0.041 0 0.0 1e-06 
3.0 0.041 0 0.0 1e-06 
0.05 0.042 0 0.0 1e-06 
3.0 0.042 0 0.0 1e-06 
0.05 0.043 0 0.0 1e-06 
3.0 0.043 0 0.0 1e-06 
0.05 0.044 0 0.0 1e-06 
3.0 0.044 0 0.0 1e-06 
0.05 0.045 0 0.0 1e-06 
3.0 0.045 0 0.0 1e-06 
0.05 0.046 0 0.0 1e-06 
3.0 0.046 0 0.0 1e-06 
0.05 0.047 0 0.0 1e-06 
3.0 0.047 0 0.0 1e-06 
0.05 0.048 0 0.0 1e-06 
3.0 0.048 0 0.0 1e-06 
0.05 0.049 0 0.0 1e-06 
3.0 0.049 0 0.0 1e-06 
0.05 0.05 0 0.0 1e-06 
3.0 0.05 0 0.0 1e-06 
0.05 0.051 0 0.0 1e-06 
3.0 0.051 0 0.0 1e-06 
0.05 0.052 0 0.0 1e-06 
3.0 0.052 0 0.0 1e-06 
0.05 0.053 0 0.0 1e-06 
3.0 0.053 0 0.0 1e-06 
0.05 0.054 0 0.0 1e-06 
3.0 0.054 0 0.0 1e-06 
0.05 0.055 0 0.0 1e-06 
3.0 0.055 0 0.0 1e-06 
0.05 0.056 0 0.0 1e-06 
3.0 0.056 0 0.0 1e-06 
0.05 0.057 0 0.0 1e-06 
3.0 0.057 0 0.0 1e-06 
0.05 0.058 0 0.0 1e-06 
3.0 0.058 0 0.0 1e-06 
0.05 0.059 0 0.0 1e-06 
3.0 0.059 0 0.0 1e-06 
0.05 0.06 0 0.0 1e-06 
3.0 0.06 0 0.0 1e-06 
0.05 0.061 0 0.0 1e-06 
3.0 0.061 0 0.0 1e-06 
0.05 0.062 0 0.0 1e-06 
3.0 0.062 0 0.0 1e-06 
0.05 0.063 0 0.0 1e-06 
3.0 0.063 0 0.0 1e-06 
0.05 0.064 0 0.0 1e-06 
3.0 0.064 0 0.0 1e-06 
0.05 0.065 0 0.0 1e-06 
3.0 0.065 0 0.0 1e-06 
0.05 0.066 0 0.0 1e-06 
3.0 0.066 0 0.0 1e-06 
0.05 0.067 0 0.0 1e-06 
3.0 0.067 0 0.0 1e-06 
0.05 0.068 0 0.0 1e-06 
3.0 0.068 0 0.0 1e-06 
0.05 0.069 0 0.0 1e-06 
3.0 0.069 0 0.0 1e-06 
0.05 0.07 0 0.0 1e-06 
3.0 0.07 0 0.0 1e-06 
0.05 0.071 0 0.0 1e-06 
3.0 0.071 0 0.0 1e-06 
0.05 0.072 0 0.0 1e-06 
3.0 0.072 0 0.0 1e-06 
0.05 0.073 0 0.0 1e-06 
3.0 0.073 0 0.0 1e-06 
0.05 0.074 0 0.0 1e-06 
3.0 0.074 0 0.0 1e-06 
0.05 0.075 0 0.0 1e-06 
3.0 0.075 0 0.0 1e-06 
0.05 0.076 0 0.0 1e-06 
3.0 0.076 0 0.0 1e-06 
0.05 0.077 0 0.0 1e-06 
3.0 0.077 0 0.0 1e-06 
0.05 0.078 0 0.0 1e-06 
3.0 0.078 0 0.0 1e-06 
0.05 0.079 0 0.0 1e-06 
3.0 0.079 0 0.0 1e-06 
0.05 0.08 0 0.0 1e-06 
3.0 0.08 0 0.0 1e-06 
0.05 0.081 0 0.0 1e-06 
3.0 0.081 0 0.0 1e-06 
0.05 0.082 0 0.0 1e-06 
3.0 0.082 0 0.0 1e-06 
0.05 0.083 0 0.0 1e-06 
3.0 0.083 0 0.0 1e-06 
0.05 0.084 0 0.0 1e-06 
3.0 0.084 0 0.0 1e-06 
0.05 0.085 0 0.0 1e-06 
3.0 0.085 0 0.0 1e-06 
0.05 0.086 0 0.0 1e-06 
3.0 0.086 0 0.0 1e-06 
0.05 0.087 0 0.0 1e-06 
3.0 0.087 0 0.0 1e-06 
0.05 0.088 0 0.0 1e-06 
3.0 0.088 0 0.0 1e-06 
0.05 0.089 0 0.0 1e-06 
3.0 0.089 0 0.0 1e-06 
0.05 0.09 0 0.0 1e-06 
3.0 0.09 0 0.0 1e-06 
0.05 0.091 0 0.0 1e-06 
3.0 0.091 0 0.0 1e-06 
0.05 0.092 0 0.0 1e-06 
3.0 0.092 0 0.0 1e-06 
0.05 0.093 0 0.0 1e-06 
3.0 0.093 0 0.0 1e-06 
0.05 0.094 0 0.0 1e-06 
3.0 0.094 0 0.0 1e-06 
0.05 0.095 0 0.0 1e-06 
3.0 0.095 0 0.0 1e-06 
0.05 0.096 0 0.0 1e-06 
3.0 0.096 0 0.0 1e-06 
0.05 0.097 0 0.0 1e-06 
3.0 0.097 0 0.0 1e-06 
0.05 0.098 0 0.0 1e-06 
3.0 0.098 0 0.0 1e-06 
0.05 0.099 0 0.0 1e-06 
3.0 0.099 0 0.0 1e-06 
0.05 0.1 0 0.0 1e-06 
3.0 0.1 0 0.0 1e-06 
0.05 0.101 0 0.0 1e-06 
3.0 0.101 0 0.0 1e-06 
0.05 0.102 0 0.0 1e-06 
3.0 0.102 0 0.0 1e-06 
0.05 0.103 0 0.0 1e-06 
3.0 0.103 0 0.0 1e-06 
0.05 0.104 0 0.0 1e-06 
3.0 0.104 0 0.0 1e-06 
0.05 0.105 0 0.0 1e-06 
3.0 0.105 0 0.0 1e-06 
0.05 0.106 0 0.0 1e-06 
3.0 0.106 0 0.0 1e-06 
0.05 0.107 0 0.0 1e-06 
3.0 0.107 0 0.0 1e-06 
0.05 0.108 0 0.0 1e-06 
3.0 0.108 0 0.0 1e-06 
0.05 0.109 0 0.0 1e-06 
3.0 0.109 0 0.0 1e-06 
0.05 0.11 0 0.0 1e-06 
3.0 0.11 0 0.0 1e-06 
0.05 0.111 0 0.0 1e-06 
3.0 0.111 0 0.0 1e-06 
0.05 0.112 0 0.0 1e-06 
3.0 0.112 0 0.0 1e-06 
0.05 0.113 0 0.0 1e-06 
3.0 0.113 0 0.0 1e-06 
0.05 0.114 0 0.0 1e-06 
3.0 0.114 0 0.0 1e-06 
0.05 0.115 0 0.0 1e-06 
3.0 0.115 0 0.0 1e-06 
0.05 0.116 0 0.0 1e-06 
3.0 0.116 0 0.0 1e-06 
0.05 0.117 0 0.0 1e-06 
3.0 0.117 0 0.0 1e-06 
0.05 0.118 0 0.0 1e-06 
3.0 0.118 0 0.0 1e-06 
0.05 0.119 0 0.0 1e-06 
3.0 0.119 0 0.0 1e-06 
0.05 0.12 0 0.0 1e-06 
3.0 0.12 0 0.0 1e-06 
0.05 0.121 0 0.0 1e-06 
3.0 0.121 0 0.0 1e-06 
0.05 0.122 0 0.0 1e-06 
3.0 0.122 0 0.0 1e-06 
0.05 0.123 0 0.0 1e-06 
3.0 0.123 0 0.0 1e-06 
0.05 0.124 0 0.0 1e-06 
3.0 0.124 0 0.0 1e-06 
0.05 0.125 0 0.0 1e-06 
3.0 0.125 0 0.0 1e-06 
0.05 0.126 0 0.0 1e-06 
3.0 0.126 0 0.0 1e-06 
0.05 0.127 0 0.0 1e-06 
3.0 0.127 0 0.0 1e-06 
0.05 0.128 0 0.0 1e-06 
3.0 0.128 0 0.0 1e-06 
0.05 0.129 0 0.0 1e-06 
3.0 0.129 0 0.0 1e-06 
0.05 0.13 0 0.0 1e-06 
3.0 0.13 0 0.0 1e-06 
0.05 0.131 0 0.0 1e-06 
3.0 0.131 0 0.0 1e-06 
0.05 0.132 0 0.0 1e-06 
3.0 0.132 0 0.0 1e-06 
0.05 0.133 0 0.0 1e-06 
3.0 0.133 0 0.0 1e-06 
0.05 0.134 0 0.0 1e-06 
3.0 0.134 0 0.0 1e-06 
0.05 0.135 0 0.0 1e-06 
3.0 0.135 0 0.0 1e-06 
0.05 0.136 0 0.0 1e-06 
3.0 0.136 0 0.0 1e-06 
0.05 0.137 0 0.0 1e-06 
3.0 0.137 0 0.0 1e-06 
0.05 0.138 0 0.0 1e-06 
3.0 0.138 0 0.0 1e-06 
0.05 0.139 0 0.0 1e-06 
3.0 0.139 0 0.0 1e-06 
0.05 0.14 0 0.0 1e-06 
3.0 0.14 0 0.0 1e-06 
0.05 0.141 0 0.0 1e-06 
3.0 0.141 0 0.0 1e-06 
0.05 0.142 0 0.0 1e-06 
3.0 0.142 0 0.0 1e-06 
0.05 0.143 0 0.0 1e-06 
3.0 0.143 0 0.0 1e-06 
0.05 0.144 0 0.0 1e-06 
3.0 0.144 0 0.0 1e-06 
0.05 0.145 0 0.0 1e-06 
3.0 0.145 0 0.0 1e-06 
0.05 0.146 0 0.0 1e-06 
3.0 0.146 0 0.0 1e-06 
0.05 0.147 0 0.0 1e-06 
3.0 0.147 0 0.0 1e-06 
0.05 0.148 0 0.0 1e-06 
3.0 0.148 0 0.0 1e-06 
0.05 0.149 0 0.0 1e-06 
3.0 0.149 0 0.0 1e-06 
0.05 0.15 0 0.0 1e-06 
3.0 0.15 0 0.0 1e-06 
0.05 0.151 0 0.0 1e-06 
3.0 0.151 0 0.0 1e-06 
0.05 0.152 0 0.0 1e-06 
3.0 0.152 0 0.0 1e-06 
0.05 0.153 0 0.0 1e-06 
3.0 0.153 0 0.0 1e-06 
0.05 0.154 0 0.0 1e-06 
3.0 0.154 0 0.0 1e-06 
0.05 0.155 0 0.0 1e-06 
3.0 0.155 0 0.0 1e-06 
0.05 0.156 0 0.0 1e-06 
3.0 0.156 0 0.0 1e-06 
0.05 0.157 0 0.0 1e-06 
3.0 0.157 0 0.0 1e-06 
0.05 0.158 0 0.0 1e-06 
3.0 0.158 0 0.0 1e-06 
0.05 0.159 0 0.0 1e-06 
3.0 0.159 0 0.0 1e-06 
0.05 0.16 0 0.0 1e-06 
3.0 0.16 0 0.0 1e-06 
0.05 0.161 0 0.0 1e-06 
3.0 0.161 0 0.0 1e-06 
0.05 0.162 0 0.0 1e-06 
3.0 0.162 0 0.0 1e-06 
0.05 0.163 0 0.0 1e-06 
3.0 0.163 0 0.0 1e-06 
0.05 0.164 0 0.0 1e-06 
3.0 0.164 0 0.0 1e-06 
0.05 0.165 0 0.0 1e-06 
3.0 0.165 0 0.0 1e-06 
0.05 0.166 0 0.0 1e-06 
3.0 0.166 0 0.0 1e-06 
0.05 0.167 0 0.0 1e-06 
3.0 0.167 0 0.0 1e-06 
0.05 0.168 0 0.0 1e-06 
3.0 0.168 0 0.0 1e-06 
0.05 0.169 0 0.0 1e-06 
3.0 0.169 0 0.0 1e-06 
0.05 0.17 0 0.0 1e-06 
3.0 0.17 0 0.0 1e-06 
0.05 0.171 0 0.0 1e-06 
3.0 0.171 0 0.0 1e-06 
0.05 0.172 0 0.0 1e-06 
3.0 0.172 0 0.0 1e-06 
0.05 0.173 0 0.0 1e-06 
3.0 0.173 0 0.0 1e-06 
0.05 0.174 0 0.0 1e-06 
3.0 0.174 0 0.0 1e-06 
0.05 0.175 0 0.0 1e-06 
3.0 0.175 0 0.0 1e-06 
0.05 0.176 0 0.0 1e-06 
3.0 0.176 0 0.0 1e-06 
0.05 0.177 0 0.0 1e-06 
3.0 0.177 0 0.0 1e-06 
0.05 0.178 0 0.0 1e-06 
3.0 0.178 0 0.0 1e-06 
0.05 0.179 0 0.0 1e-06 
3.0 0.179 0 0.0 1e-06 
0.05 0.18 0 0.0 1e-06 
3.0 0.18 0 0.0 1e-06 
0.05 0.181 0 0.0 1e-06 
3.0 0.181 0 0.0 1e-06 
0.05 0.182 0 0.0 1e-06 
3.0 0.182 0 0.0 1e-06 
0.05 0.183 0 0.0 1e-06 
3.0 0.183 0 0.0 1e-06 
0.05 0.184 0 0.0 1e-06 
3.0 0.184 0 0.0 1e-06 
0.05 0.185 0 0.0 1e-06 
3.0 0.185 0 0.0 1e-06 
0.05 0.186 0 0.0 1e-06 
3.0 0.186 0 0.0 1e-06 
0.05 0.187 0 0.0 1e-06 
3.0 0.187 0 0.0 1e-06 
0.05 0.188 0 0.0 1e-06 
3.0 0.188 0 0.0 1e-06 
0.05 0.189 0 0.0 1e-06 
3.0 0.189 0 0.0 1e-06 
0.05 0.19 0 0.0 1e-06 
3.0 0.19 0 0.0 1e-06 
0.05 0.191 0 0.0 1e-06 
3.0 0.191 0 0.0 1e-06 
0.05 0.192 0 0.0 1e-06 
3.0 0.192 0 0.0 1e-06 
0.05 0.193 0 0.0 1e-06 
3.0 0.193 0 0.0 1e-06 
0.05 0.194 0 0.0 1e-06 
3.0 0.194 0 0.0 1e-06 
0.05 0.195 0 0.0 1e-06 
3.0 0.195 0 0.0 1e-06 
0.05 0.196 0 0.0 1e-06 
3.0 0.196 0 0.0 1e-06 
0.05 0.197 0 0.0 1e-06 
3.0 0.197 0 0.0 1e-06 
0.05 0.198 0 0.0 1e-06 
3.0 0.198 0 0.0 1e-06 
0.05 0.199 0 0.0 1e-06 
3.0 0.199 0 0.0 1e-06 
0.05 0.2 0 0.0 1e-06 
3.0 0.2 0 0.0 1e-06 
0.05 0.201 0 0.0 1e-06 
3.0 0.201 0 0.0 1e-06 
0.05 0.202 0 0.0 1e-06 
3.0 0.202 0 0.0 1e-06 
0.05 0.203 0 0.0 1e-06 
3.0 0.203 0 0.0 1e-06 
0.05 0.204 0 0.0 1e-06 
3.0 0.204 0 0.0 1e-06 
0.05 0.205 0 0.0 1e-06 
3.0 0.205 0 0.0 1e-06 
0.05 0.206 0 0.0 1e-06 
3.0 0.206 0 0.0 1e-06 
0.05 0.207 0 0.0 1e-06 
3.0 0.207 0 0.0 1e-06 
0.05 0.208 0 0.0 1e-06 
3.0 0.208 0 0.0 1e-06 
0.05 0.209 0 0.0 1e-06 
3.0 0.209 0 0.0 1e-06 
0.05 0.21 0 0.0 1e-06 
3.0 0.21 0 0.0 1e-06 
0.05 0.211 0 0.0 1e-06 
3.0 0.211 0 0.0 1e-06 
0.05 0.212 0 0.0 1e-06 
3.0 0.212 0 0.0 1e-06 
0.05 0.213 0 0.0 1e-06 
3.0 0.213 0 0.0 1e-06 
0.05 0.214 0 0.0 1e-06 
3.0 0.214 0 0.0 1e-06 
0.05 0.215 0 0.0 1e-06 
3.0 0.215 0 0.0 1e-06 
0.05 0.216 0 0.0 1e-06 
3.0 0.216 0 0.0 1e-06 
0.05 0.217 0 0.0 1e-06 
3.0 0.217 0 0.0 1e-06 
0.05 0.218 0 0.0 1e-06 
3.0 0.218 0 0.0 1e-06 
0.05 0.219 0 0.0 1e-06 
3.0 0.219 0 0.0 1e-06 
0.05 0.22 0 0.0 1e-06 
3.0 0.22 0 0.0 1e-06 
0.05 0.221 0 0.0 1e-06 
3.0 0.221 0 0.0 1e-06 
0.05 0.222 0 0.0 1e-06 
3.0 0.222 0 0.0 1e-06 
0.05 0.223 0 0.0 1e-06 
3.0 0.223 0 0.0 1e-06 
0.05 0.224 0 0.0 1e-06 
3.0 0.224 0 0.0 1e-06 
0.05 0.225 0 0.0 1e-06 
3.0 0.225 0 0.0 1e-06 
0.05 0.226 0 0.0 1e-06 
3.0 0.226 0 0.0 1e-06 
0.05 0.227 0 0.0 1e-06 
3.0 0.227 0 0.0 1e-06 
0.05 0.228 0 0.0 1e-06 
3.0 0.228 0 0.0 1e-06 
0.05 0.229 0 0.0 1e-06 
3.0 0.229 0 0.0 1e-06 
0.05 0.23 0 0.0 1e-06 
3.0 0.23 0 0.0 1e-06 
0.05 0.231 0 0.0 1e-06 
3.0 0.231 0 0.0 1e-06 
0.05 0.232 0 0.0 1e-06 
3.0 0.232 0 0.0 1e-06 
0.05 0.233 0 0.0 1e-06 
3.0 0.233 0 0.0 1e-06 
0.05 0.234 0 0.0 1e-06 
3.0 0.234 0 0.0 1e-06 
0.05 0.235 0 0.0 1e-06 
3.0 0.235 0 0.0 1e-06 
0.05 0.236 0 0.0 1e-06 
3.0 0.236 0 0.0 1e-06 
0.05 0.237 0 0.0 1e-06 
3.0 0.237 0 0.0 1e-06 
0.05 0.238 0 0.0 1e-06 
3.0 0.238 0 0.0 1e-06 
0.05 0.239 0 0.0 1e-06 
3.0 0.239 0 0.0 1e-06 
0.05 0.24 0 0.0 1e-06 
3.0 0.24 0 0.0 1e-06 
0.05 0.241 0 0.0 1e-06 
3.0 0.241 0 0.0 1e-06 
0.05 0.242 0 0.0 1e-06 
3.0 0.242 0 0.0 1e-06 
0.05 0.243 0 0.0 1e-06 
3.0 0.243 0 0.0 1e-06 
0.05 0.244 0 0.0 1e-06 
3.0 0.244 0 0.0 1e-06 
0.05 0.245 0 0.0 1e-06 
3.0 0.245 0 0.0 1e-06 
0.05 0.246 0 0.0 1e-06 
3.0 0.246 0 0.0 1e-06 
0.05 0.247 0 0.0 1e-06 
3.0 0.247 0 0.0 1e-06 
0.05 0.248 0 0.0 1e-06 
3.0 0.248 0 0.0 1e-06 
0.05 0.249 0 0.0 1e-06 
3.0 0.249 0 0.0 1e-06 
0.05 0.25 0 0.0 1e-06 
3.0 0.25 0 0.0 1e-06 
0.05 0.251 0 0.0 1e-06 
3.0 0.251 0 0.0 1e-06 
0.05 0.252 0 0.0 1e-06 
3.0 0.252 0 0.0 1e-06 
0.05 0.253 0 0.0 1e-06 
3.0 0.253 0 0.0 1e-06 
0.05 0.254 0 0.0 1e-06 
3.0 0.254 0 0.0 1e-06 
0.05 0.255 0 0.0 1e-06 
3.0 0.255 0 0.0 1e-06 
0.05 0.256 0 0.0 1e-06 
3.0 0.256 0 0.0 1e-06 
0.05 0.257 0 0.0 1e-06 
3.0 0.257 0 0.0 1e-06 
0.05 0.258 0 0.0 1e-06 
3.0 0.258 0 0.0 1e-06 
0.05 0.259 0 0.0 1e-06 
3.0 0.259 0 0.0 1e-06 
0.05 0.26 0 0.0 1e-06 
3.0 0.26 0 0.0 1e-06 
0.05 0.261 0 0.0 1e-06 
3.0 0.261 0 0.0 1e-06 
0.05 0.262 0 0.0 1e-06 
3.0 0.262 0 0.0 1e-06 
0.05 0.263 0 0.0 1e-06 
3.0 0.263 0 0.0 1e-06 
0.05 0.264 0 0.0 1e-06 
3.0 0.264 0 0.0 1e-06 
0.05 0.265 0 0.0 1e-06 
3.0 0.265 0 0.0 1e-06 
0.05 0.266 0 0.0 1e-06 
3.0 0.266 0 0.0 1e-06 
0.05 0.267 0 0.0 1e-06 
3.0 0.267 0 0.0 1e-06 
0.05 0.268 0 0.0 1e-06 
3.0 0.268 0 0.0 1e-06 
0.05 0.269 0 0.0 1e-06 
3.0 0.269 0 0.0 1e-06 
0.05 0.27 0 0.0 1e-06 
3.0 0.27 0 0.0 1e-06 
0.05 0.271 0 0.0 1e-06 
3.0 0.271 0 0.0 1e-06 
0.05 0.272 0 0.0 1e-06 
3.0 0.272 0 0.0 1e-06 
0.05 0.273 0 0.0 1e-06 
3.0 0.273 0 0.0 1e-06 
0.05 0.274 0 0.0 1e-06 
3.0 0.274 0 0.0 1e-06 
0.05 0.275 0 0.0 1e-06 
3.0 0.275 0 0.0 1e-06 
0.05 0.276 0 0.0 1e-06 
3.0 0.276 0 0.0 1e-06 
0.05 0.277 0 0.0 1e-06 
3.0 0.277 0 0.0 1e-06 
0.05 0.278 0 0.0 1e-06 
3.0 0.278 0 0.0 1e-06 
0.05 0.279 0 0.0 1e-06 
3.0 0.279 0 0.0 1e-06 
0.05 0.28 0 0.0 1e-06 
3.0 0.28 0 0.0 1e-06 
0.05 0.281 0 0.0 1e-06 
3.0 0.281 0 0.0 1e-06 
0.05 0.282 0 0.0 1e-06 
3.0 0.282 0 0.0 1e-06 
0.05 0.283 0 0.0 1e-06 
3.0 0.283 0 0.0 1e-06 
0.05 0.284 0 0.0 1e-06 
3.0 0.284 0 0.0 1e-06 
0.05 0.285 0 0.0 1e-06 
3.0 0.285 0 0.0 1e-06 
0.05 0.286 0 0.0 1e-06 
3.0 0.286 0 0.0 1e-06 
0.05 0.287 0 0.0 1e-06 
3.0 0.287 0 0.0 1e-06 
0.05 0.288 0 0.0 1e-06 
3.0 0.288 0 0.0 1e-06 
0.05 0.289 0 0.0 1e-06 
3.0 0.289 0 0.0 1e-06 
0.05 0.29 0 0.0 1e-06 
3.0 0.29 0 0.0 1e-06 
0.05 0.291 0 0.0 1e-06 
3.0 0.291 0 0.0 1e-06 
0.05 0.292 0 0.0 1e-06 
3.0 0.292 0 0.0 1e-06 
0.05 0.293 0 0.0 1e-06 
3.0 0.293 0 0.0 1e-06 
0.05 0.294 0 0.0 1e-06 
3.0 0.294 0 0.0 1e-06 
0.05 0.295 0 0.0 1e-06 
3.0 0.295 0 0.0 1e-06 
0.05 0.296 0 0.0 1e-06 
3.0 0.296 0 0.0 1e-06 
0.05 0.297 0 0.0 1e-06 
3.0 0.297 0 0.0 1e-06 
0.05 0.298 0 0.0 1e-06 
3.0 0.298 0 0.0 1e-06 
0.05 0.299 0 0.0 1e-06 
3.0 0.299 0 0.0 1e-06 
0.05 0.3 0 0.0 1e-06 
3.0 0.3 0 0.0 1e-06 
0.05 0.301 0 0.0 1e-06 
3.0 0.301 0 0.0 1e-06 
0.05 0.302 0 0.0 1e-06 
3.0 0.302 0 0.0 1e-06 
0.05 0.303 0 0.0 1e-06 
3.0 0.303 0 0.0 1e-06 
0.05 0.304 0 0.0 1e-06 
3.0 0.304 0 0.0 1e-06 
0.05 0.305 0 0.0 1e-06 
3.0 0.305 0 0.0 1e-06 
0.05 0.306 0 0.0 1e-06 
3.0 0.306 0 0.0 1e-06 
0.05 0.307 0 0.0 1e-06 
3.0 0.307 0 0.0 1e-06 
0.05 0.308 0 0.0 1e-06 
3.0 0.308 0 0.0 1e-06 
0.05 0.309 0 0.0 1e-06 
3.0 0.309 0 0.0 1e-06 
0.05 0.31 0 0.0 1e-06 
3.0 0.31 0 0.0 1e-06 
0.05 0.311 0 0.0 1e-06 
3.0 0.311 0 0.0 1e-06 
0.05 0.312 0 0.0 1e-06 
3.0 0.312 0 0.0 1e-06 
0.05 0.313 0 0.0 1e-06 
3.0 0.313 0 0.0 1e-06 
0.05 0.314 0 0.0 1e-06 
3.0 0.314 0 0.0 1e-06 
0.05 0.315 0 0.0 1e-06 
3.0 0.315 0 0.0 1e-06 
0.05 0.316 0 0.0 1e-06 
3.0 0.316 0 0.0 1e-06 
0.05 0.317 0 0.0 1e-06 
3.0 0.317 0 0.0 1e-06 
0.05 0.318 0 0.0 1e-06 
3.0 0.318 0 0.0 1e-06 
0.05 0.319 0 0.0 1e-06 
3.0 0.319 0 0.0 1e-06 
0.05 0.32 0 0.0 1e-06 
3.0 0.32 0 0.0 1e-06 
0.05 0.321 0 0.0 1e-06 
3.0 0.321 0 0.0 1e-06 
0.05 0.322 0 0.0 1e-06 
3.0 0.322 0 0.0 1e-06 
0.05 0.323 0 0.0 1e-06 
3.0 0.323 0 0.0 1e-06 
0.05 0.324 0 0.0 1e-06 
3.0 0.324 0 0.0 1e-06 
0.05 0.325 0 0.0 1e-06 
3.0 0.325 0 0.0 1e-06 
0.05 0.326 0 0.0 1e-06 
3.0 0.326 0 0.0 1e-06 
0.05 0.327 0 0.0 1e-06 
3.0 0.327 0 0.0 1e-06 
0.05 0.328 0 0.0 1e-06 
3.0 0.328 0 0.0 1e-06 
0.05 0.329 0 0.0 1e-06 
3.0 0.329 0 0.0 1e-06 
0.05 0.33 0 0.0 1e-06 
3.0 0.33 0 0.0 1e-06 
0.05 0.331 0 0.0 1e-06 
3.0 0.331 0 0.0 1e-06 
0.05 0.332 0 0.0 1e-06 
3.0 0.332 0 0.0 1e-06 
0.05 0.333 0 0.0 1e-06 
3.0 0.333 0 0.0 1e-06 
0.05 0.334 0 0.0 1e-06 
3.0 0.334 0 0.0 1e-06 
0.05 0.335 0 0.0 1e-06 
3.0 0.335 0 0.0 1e-06 
0.05 0.336 0 0.0 1e-06 
3.0 0.336 0 0.0 1e-06 
0.05 0.337 0 0.0 1e-06 
3.0 0.337 0 0.0 1e-06 
0.05 0.338 0 0.0 1e-06 
3.0 0.338 0 0.0 1e-06 
0.05 0.339 0 0.0 1e-06 
3.0 0.339 0 0.0 1e-06 
0.05 0.34 0 0.0 1e-06 
3.0 0.34 0 0.0 1e-06 
0.05 0.341 0 0.0 1e-06 
3.0 0.341 0 0.0 1e-06 
0.05 0.342 0 0.0 1e-06 
3.0 0.342 0 0.0 1e-06 
0.05 0.343 0 0.0 1e-06 
3.0 0.343 0 0.0 1e-06 
0.05 0.344 0 0.0 1e-06 
3.0 0.344 0 0.0 1e-06 
0.05 0.345 0 0.0 1e-06 
3.0 0.345 0 0.0 1e-06 
0.05 0.346 0 0.0 1e-06 
3.0 0.346 0 0.0 1e-06 
0.05 0.347 0 0.0 1e-06 
3.0 0.347 0 0.0 1e-06 
0.05 0.348 0 0.0 1e-06 
3.0 0.348 0 0.0 1e-06 
0.05 0.349 0 0.0 1e-06 
3.0 0.349 0 0.0 1e-06 
0.05 0.35 0 0.0 1e-06 
3.0 0.35 0 0.0 1e-06 
0.05 0.351 0 0.0 1e-06 
3.0 0.351 0 0.0 1e-06 
0.05 0.352 0 0.0 1e-06 
3.0 0.352 0 0.0 1e-06 
0.05 0.353 0 0.0 1e-06 
3.0 0.353 0 0.0 1e-06 
0.05 0.354 0 0.0 1e-06 
3.0 0.354 0 0.0 1e-06 
0.05 0.355 0 0.0 1e-06 
3.0 0.355 0 0.0 1e-06 
0.05 0.356 0 0.0 1e-06 
3.0 0.356 0 0.0 1e-06 
0.05 0.357 0 0.0 1e-06 
3.0 0.357 0 0.0 1e-06 
0.05 0.358 0 0.0 1e-06 
3.0 0.358 0 0.0 1e-06 
0.05 0.359 0 0.0 1e-06 
3.0 0.359 0 0.0 1e-06 
0.05 0.36 0 0.0 1e-06 
3.0 0.36 0 0.0 1e-06 
0.05 0.361 0 0.0 1e-06 
3.0 0.361 0 0.0 1e-06 
0.05 0.362 0 0.0 1e-06 
3.0 0.362 0 0.0 1e-06 
0.05 0.363 0 0.0 1e-06 
3.0 0.363 0 0.0 1e-06 
0.05 0.364 0 0.0 1e-06 
3.0 0.364 0 0.0 1e-06 
0.05 0.365 0 0.0 1e-06 
3.0 0.365 0 0.0 1e-06 
0.05 0.366 0 0.0 1e-06 
3.0 0.366 0 0.0 1e-06 
0.05 0.367 0 0.0 1e-06 
3.0 0.367 0 0.0 1e-06 
0.05 0.368 0 0.0 1e-06 
3.0 0.368 0 0.0 1e-06 
0.05 0.369 0 0.0 1e-06 
3.0 0.369 0 0.0 1e-06 
0.05 0.37 0 0.0 1e-06 
3.0 0.37 0 0.0 1e-06 
0.05 0.371 0 0.0 1e-06 
3.0 0.371 0 0.0 1e-06 
0.05 0.372 0 0.0 1e-06 
3.0 0.372 0 0.0 1e-06 
0.05 0.373 0 0.0 1e-06 
3.0 0.373 0 0.0 1e-06 
0.05 0.374 0 0.0 1e-06 
3.0 0.374 0 0.0 1e-06 
0.05 0.375 0 0.0 1e-06 
3.0 0.375 0 0.0 1e-06 
0.05 0.376 0 0.0 1e-06 
3.0 0.376 0 0.0 1e-06 
0.05 0.377 0 0.0 1e-06 
3.0 0.377 0 0.0 1e-06 
0.05 0.378 0 0.0 1e-06 
3.0 0.378 0 0.0 1e-06 
0.05 0.379 0 0.0 1e-06 
3.0 0.379 0 0.0 1e-06 
0.05 0.38 0 0.0 1e-06 
3.0 0.38 0 0.0 1e-06 
0.05 0.381 0 0.0 1e-06 
3.0 0.381 0 0.0 1e-06 
0.05 0.382 0 0.0 1e-06 
3.0 0.382 0 0.0 1e-06 
0.05 0.383 0 0.0 1e-06 
3.0 0.383 0 0.0 1e-06 
0.05 0.384 0 0.0 1e-06 
3.0 0.384 0 0.0 1e-06 
0.05 0.385 0 0.0 1e-06 
3.0 0.385 0 0.0 1e-06 
0.05 0.386 0 0.0 1e-06 
3.0 0.386 0 0.0 1e-06 
0.05 0.387 0 0.0 1e-06 
3.0 0.387 0 0.0 1e-06 
0.05 0.388 0 0.0 1e-06 
3.0 0.388 0 0.0 1e-06 
0.05 0.389 0 0.0 1e-06 
3.0 0.389 0 0.0 1e-06 
0.05 0.39 0 0.0 1e-06 
3.0 0.39 0 0.0 1e-06 
0.05 0.391 0 0.0 1e-06 
3.0 0.391 0 0.0 1e-06 
0.05 0.392 0 0.0 1e-06 
3.0 0.392 0 0.0 1e-06 
0.05 0.393 0 0.0 1e-06 
3.0 0.393 0 0.0 1e-06 
0.05 0.394 0 0.0 1e-06 
3.0 0.394 0 0.0 1e-06 
0.05 0.395 0 0.0 1e-06 
3.0 0.395 0 0.0 1e-06 
0.05 0.396 0 0.0 1e-06 
3.0 0.396 0 0.0 1e-06 
0.05 0.397 0 0.0 1e-06 
3.0 0.397 0 0.0 1e-06 
0.05 0.398 0 0.0 1e-06 
3.0 0.398 0 0.0 1e-06 
0.05 0.399 0 0.0 1e-06 
3.0 0.399 0 0.0 1e-06 
0.05 0.4 0 0.0 1e-06 
3.0 0.4 0 0.0 1e-06 
0.05 0.401 0 0.0 1e-06 
3.0 0.401 0 0.0 1e-06 
0.05 0.402 0 0.0 1e-06 
3.0 0.402 0 0.0 1e-06 
0.05 0.403 0 0.0 1e-06 
3.0 0.403 0 0.0 1e-06 
0.05 0.404 0 0.0 1e-06 
3.0 0.404 0 0.0 1e-06 
0.05 0.405 0 0.0 1e-06 
3.0 0.405 0 0.0 1e-06 
0.05 0.406 0 0.0 1e-06 
3.0 0.406 0 0.0 1e-06 
0.05 0.407 0 0.0 1e-06 
3.0 0.407 0 0.0 1e-06 
0.05 0.408 0 0.0 1e-06 
3.0 0.408 0 0.0 1e-06 
0.05 0.409 0 0.0 1e-06 
3.0 0.409 0 0.0 1e-06 
0.05 0.41 0 0.0 1e-06 
3.0 0.41 0 0.0 1e-06 
0.05 0.411 0 0.0 1e-06 
3.0 0.411 0 0.0 1e-06 
0.05 0.412 0 0.0 1e-06 
3.0 0.412 0 0.0 1e-06 
0.05 0.413 0 0.0 1e-06 
3.0 0.413 0 0.0 1e-06 
0.05 0.414 0 0.0 1e-06 
3.0 0.414 0 0.0 1e-06 
0.05 0.415 0 0.0 1e-06 
3.0 0.415 0 0.0 1e-06 
0.05 0.416 0 0.0 1e-06 
3.0 0.416 0 0.0 1e-06 
0.05 0.417 0 0.0 1e-06 
3.0 0.417 0 0.0 1e-06 
0.05 0.418 0 0.0 1e-06 
3.0 0.418 0 0.0 1e-06 
0.05 0.419 0 0.0 1e-06 
3.0 0.419 0 0.0 1e-06 
0.05 0.42 0 0.0 1e-06 
3.0 0.42 0 0.0 1e-06 
0.05 0.421 0 0.0 1e-06 
3.0 0.421 0 0.0 1e-06 
0.05 0.422 0 0.0 1e-06 
3.0 0.422 0 0.0 1e-06 
0.05 0.423 0 0.0 1e-06 
3.0 0.423 0 0.0 1e-06 
0.05 0.424 0 0.0 1e-06 
3.0 0.424 0 0.0 1e-06 
0.05 0.425 0 0.0 1e-06 
3.0 0.425 0 0.0 1e-06 
0.05 0.426 0 0.0 1e-06 
3.0 0.426 0 0.0 1e-06 
0.05 0.427 0 0.0 1e-06 
3.0 0.427 0 0.0 1e-06 
0.05 0.428 0 0.0 1e-06 
3.0 0.428 0 0.0 1e-06 
0.05 0.429 0 0.0 1e-06 
3.0 0.429 0 0.0 1e-06 
0.05 0.43 0 0.0 1e-06 
3.0 0.43 0 0.0 1e-06 
0.05 0.431 0 0.0 1e-06 
3.0 0.431 0 0.0 1e-06 
0.05 0.432 0 0.0 1e-06 
3.0 0.432 0 0.0 1e-06 
0.05 0.433 0 0.0 1e-06 
3.0 0.433 0 0.0 1e-06 
0.05 0.434 0 0.0 1e-06 
3.0 0.434 0 0.0 1e-06 
0.05 0.435 0 0.0 1e-06 
3.0 0.435 0 0.0 1e-06 
0.05 0.436 0 0.0 1e-06 
3.0 0.436 0 0.0 1e-06 
0.05 0.437 0 0.0 1e-06 
3.0 0.437 0 0.0 1e-06 
0.05 0.438 0 0.0 1e-06 
3.0 0.438 0 0.0 1e-06 
0.05 0.439 0 0.0 1e-06 
3.0 0.439 0 0.0 1e-06 
0.05 0.44 0 0.0 1e-06 
3.0 0.44 0 0.0 1e-06 
0.05 0.441 0 0.0 1e-06 
3.0 0.441 0 0.0 1e-06 
0.05 0.442 0 0.0 1e-06 
3.0 0.442 0 0.0 1e-06 
0.05 0.443 0 0.0 1e-06 
3.0 0.443 0 0.0 1e-06 
0.05 0.444 0 0.0 1e-06 
3.0 0.444 0 0.0 1e-06 
0.05 0.445 0 0.0 1e-06 
3.0 0.445 0 0.0 1e-06 
0.05 0.446 0 0.0 1e-06 
3.0 0.446 0 0.0 1e-06 
0.05 0.447 0 0.0 1e-06 
3.0 0.447 0 0.0 1e-06 
0.05 0.448 0 0.0 1e-06 
3.0 0.448 0 0.0 1e-06 
0.05 0.449 0 0.0 1e-06 
3.0 0.449 0 0.0 1e-06 
0.05 0.45 0 0.0 1e-06 
3.0 0.45 0 0.0 1e-06 
0.05 0.451 0 0.0 1e-06 
3.0 0.451 0 0.0 1e-06 
0.05 0.452 0 0.0 1e-06 
3.0 0.452 0 0.0 1e-06 
0.05 0.453 0 0.0 1e-06 
3.0 0.453 0 0.0 1e-06 
0.05 0.454 0 0.0 1e-06 
3.0 0.454 0 0.0 1e-06 
0.05 0.455 0 0.0 1e-06 
3.0 0.455 0 0.0 1e-06 
0.05 0.456 0 0.0 1e-06 
3.0 0.456 0 0.0 1e-06 
0.05 0.457 0 0.0 1e-06 
3.0 0.457 0 0.0 1e-06 
0.05 0.458 0 0.0 1e-06 
3.0 0.458 0 0.0 1e-06 
0.05 0.459 0 0.0 1e-06 
3.0 0.459 0 0.0 1e-06 
0.05 0.46 0 0.0 1e-06 
3.0 0.46 0 0.0 1e-06 
0.05 0.461 0 0.0 1e-06 
3.0 0.461 0 0.0 1e-06 
0.05 0.462 0 0.0 1e-06 
3.0 0.462 0 0.0 1e-06 
0.05 0.463 0 0.0 1e-06 
3.0 0.463 0 0.0 1e-06 
0.05 0.464 0 0.0 1e-06 
3.0 0.464 0 0.0 1e-06 
0.05 0.465 0 0.0 1e-06 
3.0 0.465 0 0.0 1e-06 
0.05 0.466 0 0.0 1e-06 
3.0 0.466 0 0.0 1e-06 
0.05 0.467 0 0.0 1e-06 
3.0 0.467 0 0.0 1e-06 
0.05 0.468 0 0.0 1e-06 
3.0 0.468 0 0.0 1e-06 
0.05 0.469 0 0.0 1e-06 
3.0 0.469 0 0.0 1e-06 
0.05 0.47 0 0.0 1e-06 
3.0 0.47 0 0.0 1e-06 
0.05 0.471 0 0.0 1e-06 
3.0 0.471 0 0.0 1e-06 
0.05 0.472 0 0.0 1e-06 
3.0 0.472 0 0.0 1e-06 
0.05 0.473 0 0.0 1e-06 
3.0 0.473 0 0.0 1e-06 
0.05 0.474 0 0.0 1e-06 
3.0 0.474 0 0.0 1e-06 
0.05 0.475 0 0.0 1e-06 
3.0 0.475 0 0.0 1e-06 
0.05 0.476 0 0.0 1e-06 
3.0 0.476 0 0.0 1e-06 
0.05 0.477 0 0.0 1e-06 
3.0 0.477 0 0.0 1e-06 
0.05 0.478 0 0.0 1e-06 
3.0 0.478 0 0.0 1e-06 
0.05 0.479 0 0.0 1e-06 
3.0 0.479 0 0.0 1e-06 
0.05 0.48 0 0.0 1e-06 
3.0 0.48 0 0.0 1e-06 
0.05 0.481 0 0.0 1e-06 
3.0 0.481 0 0.0 1e-06 
0.05 0.482 0 0.0 1e-06 
3.0 0.482 0 0.0 1e-06 
0.05 0.483 0 0.0 1e-06 
3.0 0.483 0 0.0 1e-06 
0.05 0.484 0 0.0 1e-06 
3.0 0.484 0 0.0 1e-06 
0.05 0.485 0 0.0 1e-06 
3.0 0.485 0 0.0 1e-06 
0.05 0.486 0 0.0 1e-06 
3.0 0.486 0 0.0 1e-06 
0.05 0.487 0 0.0 1e-06 
3.0 0.487 0 0.0 1e-06 
0.05 0.488 0 0.0 1e-06 
3.0 0.488 0 0.0 1e-06 
0.05 0.489 0 0.0 1e-06 
3.0 0.489 0 0.0 1e-06 
0.05 0.49 0 0.0 1e-06 
3.0 0.49 0 0.0 1e-06 
0.05 0.491 0 0.0 1e-06 
3.0 0.491 0 0.0 1e-06 
0.05 0.492 0 0.0 1e-06 
3.0 0.492 0 0.0 1e-06 
0.05 0.493 0 0.0 1e-06 
3.0 0.493 0 0.0 1e-06 
0.05 0.494 0 0.0 1e-06 
3.0 0.494 0 0.0 1e-06 
0.05 0.495 0 0.0 1e-06 
3.0 0.495 0 0.0 1e-06 
0.05 0.496 0 0.0 1e-06 
3.0 0.496 0 0.0 1e-06 
0.05 0.497 0 0.0 1e-06 
3.0 0.497 0 0.0 1e-06 
0.05 0.498 0 0.0 1e-06 
3.0 0.498 0 0.0 1e-06 
0.05 0.499 0 0.0 1e-06 
3.0 0.499 0 0.0 1e-06 
0.05 0.5 0 0.0 1e-06 
3.0 0.5 0 0.0 1e-06 
0.05 0.501 0 0.0 1e-06 
3.0 0.501 0 0.0 1e-06 
0.05 0.502 0 0.0 1e-06 
3.0 0.502 0 0.0 1e-06 
0.05 0.503 0 0.0 1e-06 
3.0 0.503 0 0.0 1e-06 
0.05 0.504 0 0.0 1e-06 
3.0 0.504 0 0.0 1e-06 
0.05 0.505 0 0.0 1e-06 
3.0 0.505 0 0.0 1e-06 
0.05 0.506 0 0.0 1e-06 
3.0 0.506 0 0.0 1e-06 
0.05 0.507 0 0.0 1e-06 
3.0 0.507 0 0.0 1e-06 
0.05 0.508 0 0.0 1e-06 
3.0 0.508 0 0.0 1e-06 
0.05 0.509 0 0.0 1e-06 
3.0 0.509 0 0.0 1e-06 
0.05 0.51 0 0.0 1e-06 
3.0 0.51 0 0.0 1e-06 
0.05 0.511 0 0.0 1e-06 
3.0 0.511 0 0.0 1e-06 
0.05 0.512 0 0.0 1e-06 
3.0 0.512 0 0.0 1e-06 
0.05 0.513 0 0.0 1e-06 
3.0 0.513 0 0.0 1e-06 
0.05 0.514 0 0.0 1e-06 
3.0 0.514 0 0.0 1e-06 
0.05 0.515 0 0.0 1e-06 
3.0 0.515 0 0.0 1e-06 
0.05 0.516 0 0.0 1e-06 
3.0 0.516 0 0.0 1e-06 
0.05 0.517 0 0.0 1e-06 
3.0 0.517 0 0.0 1e-06 
0.05 0.518 0 0.0 1e-06 
3.0 0.518 0 0.0 1e-06 
0.05 0.519 0 0.0 1e-06 
3.0 0.519 0 0.0 1e-06 
0.05 0.52 0 0.0 1e-06 
3.0 0.52 0 0.0 1e-06 
0.05 0.521 0 0.0 1e-06 
3.0 0.521 0 0.0 1e-06 
0.05 0.522 0 0.0 1e-06 
3.0 0.522 0 0.0 1e-06 
0.05 0.523 0 0.0 1e-06 
3.0 0.523 0 0.0 1e-06 
0.05 0.524 0 0.0 1e-06 
3.0 0.524 0 0.0 1e-06 
0.05 0.525 0 0.0 1e-06 
3.0 0.525 0 0.0 1e-06 
0.05 0.526 0 0.0 1e-06 
3.0 0.526 0 0.0 1e-06 
0.05 0.527 0 0.0 1e-06 
3.0 0.527 0 0.0 1e-06 
0.05 0.528 0 0.0 1e-06 
3.0 0.528 0 0.0 1e-06 
0.05 0.529 0 0.0 1e-06 
3.0 0.529 0 0.0 1e-06 
0.05 0.53 0 0.0 1e-06 
3.0 0.53 0 0.0 1e-06 
0.05 0.531 0 0.0 1e-06 
3.0 0.531 0 0.0 1e-06 
0.05 0.532 0 0.0 1e-06 
3.0 0.532 0 0.0 1e-06 
0.05 0.533 0 0.0 1e-06 
3.0 0.533 0 0.0 1e-06 
0.05 0.534 0 0.0 1e-06 
3.0 0.534 0 0.0 1e-06 
0.05 0.535 0 0.0 1e-06 
3.0 0.535 0 0.0 1e-06 
0.05 0.536 0 0.0 1e-06 
3.0 0.536 0 0.0 1e-06 
0.05 0.537 0 0.0 1e-06 
3.0 0.537 0 0.0 1e-06 
0.05 0.538 0 0.0 1e-06 
3.0 0.538 0 0.0 1e-06 
0.05 0.539 0 0.0 1e-06 
3.0 0.539 0 0.0 1e-06 
0.05 0.54 0 0.0 1e-06 
3.0 0.54 0 0.0 1e-06 
0.05 0.541 0 0.0 1e-06 
3.0 0.541 0 0.0 1e-06 
0.05 0.542 0 0.0 1e-06 
3.0 0.542 0 0.0 1e-06 
0.05 0.543 0 0.0 1e-06 
3.0 0.543 0 0.0 1e-06 
0.05 0.544 0 0.0 1e-06 
3.0 0.544 0 0.0 1e-06 
0.05 0.545 0 0.0 1e-06 
3.0 0.545 0 0.0 1e-06 
0.05 0.546 0 0.0 1e-06 
3.0 0.546 0 0.0 1e-06 
0.05 0.547 0 0.0 1e-06 
3.0 0.547 0 0.0 1e-06 
0.05 0.548 0 0.0 1e-06 
3.0 0.548 0 0.0 1e-06 
0.05 0.549 0 0.0 1e-06 
3.0 0.549 0 0.0 1e-06 
0.05 0.55 0 0.0 1e-06 
3.0 0.55 0 0.0 1e-06 
0.05 0.551 0 0.0 1e-06 
3.0 0.551 0 0.0 1e-06 
0.05 0.552 0 0.0 1e-06 
3.0 0.552 0 0.0 1e-06 
0.05 0.553 0 0.0 1e-06 
3.0 0.553 0 0.0 1e-06 
0.05 0.554 0 0.0 1e-06 
3.0 0.554 0 0.0 1e-06 
0.05 0.555 0 0.0 1e-06 
3.0 0.555 0 0.0 1e-06 
0.05 0.556 0 0.0 1e-06 
3.0 0.556 0 0.0 1e-06 
0.05 0.557 0 0.0 1e-06 
3.0 0.557 0 0.0 1e-06 
0.05 0.558 0 0.0 1e-06 
3.0 0.558 0 0.0 1e-06 
0.05 0.559 0 0.0 1e-06 
3.0 0.559 0 0.0 1e-06 
0.05 0.56 0 0.0 1e-06 
3.0 0.56 0 0.0 1e-06 
0.05 0.561 0 0.0 1e-06 
3.0 0.561 0 0.0 1e-06 
0.05 0.562 0 0.0 1e-06 
3.0 0.562 0 0.0 1e-06 
0.05 0.563 0 0.0 1e-06 
3.0 0.563 0 0.0 1e-06 
0.05 0.564 0 0.0 1e-06 
3.0 0.564 0 0.0 1e-06 
0.05 0.565 0 0.0 1e-06 
3.0 0.565 0 0.0 1e-06 
0.05 0.566 0 0.0 1e-06 
3.0 0.566 0 0.0 1e-06 
0.05 0.567 0 0.0 1e-06 
3.0 0.567 0 0.0 1e-06 
0.05 0.568 0 0.0 1e-06 
3.0 0.568 0 0.0 1e-06 
0.05 0.569 0 0.0 1e-06 
3.0 0.569 0 0.0 1e-06 
0.05 0.57 0 0.0 1e-06 
3.0 0.57 0 0.0 1e-06 
0.05 0.571 0 0.0 1e-06 
3.0 0.571 0 0.0 1e-06 
0.05 0.572 0 0.0 1e-06 
3.0 0.572 0 0.0 1e-06 
0.05 0.573 0 0.0 1e-06 
3.0 0.573 0 0.0 1e-06 
0.05 0.574 0 0.0 1e-06 
3.0 0.574 0 0.0 1e-06 
0.05 0.575 0 0.0 1e-06 
3.0 0.575 0 0.0 1e-06 
0.05 0.576 0 0.0 1e-06 
3.0 0.576 0 0.0 1e-06 
0.05 0.577 0 0.0 1e-06 
3.0 0.577 0 0.0 1e-06 
0.05 0.578 0 0.0 1e-06 
3.0 0.578 0 0.0 1e-06 
0.05 0.579 0 0.0 1e-06 
3.0 0.579 0 0.0 1e-06 
0.05 0.58 0 0.0 1e-06 
3.0 0.58 0 0.0 1e-06 
0.05 0.581 0 0.0 1e-06 
3.0 0.581 0 0.0 1e-06 
0.05 0.582 0 0.0 1e-06 
3.0 0.582 0 0.0 1e-06 
0.05 0.583 0 0.0 1e-06 
3.0 0.583 0 0.0 1e-06 
0.05 0.584 0 0.0 1e-06 
3.0 0.584 0 0.0 1e-06 
0.05 0.585 0 0.0 1e-06 
3.0 0.585 0 0.0 1e-06 
0.05 0.586 0 0.0 1e-06 
3.0 0.586 0 0.0 1e-06 
0.05 0.587 0 0.0 1e-06 
3.0 0.587 0 0.0 1e-06 
0.05 0.588 0 0.0 1e-06 
3.0 0.588 0 0.0 1e-06 
0.05 0.589 0 0.0 1e-06 
3.0 0.589 0 0.0 1e-06 
0.05 0.59 0 0.0 1e-06 
3.0 0.59 0 0.0 1e-06 
0.05 0.591 0 0.0 1e-06 
3.0 0.591 0 0.0 1e-06 
0.05 0.592 0 0.0 1e-06 
3.0 0.592 0 0.0 1e-06 
0.05 0.593 0 0.0 1e-06 
3.0 0.593 0 0.0 1e-06 
0.05 0.594 0 0.0 1e-06 
3.0 0.594 0 0.0 1e-06 
0.05 0.595 0 0.0 1e-06 
3.0 0.595 0 0.0 1e-06 
0.05 0.596 0 0.0 1e-06 
3.0 0.596 0 0.0 1e-06 
0.05 0.597 0 0.0 1e-06 
3.0 0.597 0 0.0 1e-06 
0.05 0.598 0 0.0 1e-06 
3.0 0.598 0 0.0 1e-06 
0.05 0.599 0 0.0 1e-06 
3.0 0.599 0 0.0 1e-06 
0.05 0.6 0 0.0 1e-06 
3.0 0.6 0 0.0 1e-06 
0.05 0.601 0 0.0 1e-06 
3.0 0.601 0 0.0 1e-06 
0.05 0.602 0 0.0 1e-06 
3.0 0.602 0 0.0 1e-06 
0.05 0.603 0 0.0 1e-06 
3.0 0.603 0 0.0 1e-06 
0.05 0.604 0 0.0 1e-06 
3.0 0.604 0 0.0 1e-06 
0.05 0.605 0 0.0 1e-06 
3.0 0.605 0 0.0 1e-06 
0.05 0.606 0 0.0 1e-06 
3.0 0.606 0 0.0 1e-06 
0.05 0.607 0 0.0 1e-06 
3.0 0.607 0 0.0 1e-06 
0.05 0.608 0 0.0 1e-06 
3.0 0.608 0 0.0 1e-06 
0.05 0.609 0 0.0 1e-06 
3.0 0.609 0 0.0 1e-06 
0.05 0.61 0 0.0 1e-06 
3.0 0.61 0 0.0 1e-06 
0.05 0.611 0 0.0 1e-06 
3.0 0.611 0 0.0 1e-06 
0.05 0.612 0 0.0 1e-06 
3.0 0.612 0 0.0 1e-06 
0.05 0.613 0 0.0 1e-06 
3.0 0.613 0 0.0 1e-06 
0.05 0.614 0 0.0 1e-06 
3.0 0.614 0 0.0 1e-06 
0.05 0.615 0 0.0 1e-06 
3.0 0.615 0 0.0 1e-06 
0.05 0.616 0 0.0 1e-06 
3.0 0.616 0 0.0 1e-06 
0.05 0.617 0 0.0 1e-06 
3.0 0.617 0 0.0 1e-06 
0.05 0.618 0 0.0 1e-06 
3.0 0.618 0 0.0 1e-06 
0.05 0.619 0 0.0 1e-06 
3.0 0.619 0 0.0 1e-06 
0.05 0.62 0 0.0 1e-06 
3.0 0.62 0 0.0 1e-06 
0.05 0.621 0 0.0 1e-06 
3.0 0.621 0 0.0 1e-06 
0.05 0.622 0 0.0 1e-06 
3.0 0.622 0 0.0 1e-06 
0.05 0.623 0 0.0 1e-06 
3.0 0.623 0 0.0 1e-06 
0.05 0.624 0 0.0 1e-06 
3.0 0.624 0 0.0 1e-06 
0.05 0.625 0 0.0 1e-06 
3.0 0.625 0 0.0 1e-06 
0.05 0.626 0 0.0 1e-06 
3.0 0.626 0 0.0 1e-06 
0.05 0.627 0 0.0 1e-06 
3.0 0.627 0 0.0 1e-06 
0.05 0.628 0 0.0 1e-06 
3.0 0.628 0 0.0 1e-06 
0.05 0.629 0 0.0 1e-06 
3.0 0.629 0 0.0 1e-06 
0.05 0.63 0 0.0 1e-06 
3.0 0.63 0 0.0 1e-06 
0.05 0.631 0 0.0 1e-06 
3.0 0.631 0 0.0 1e-06 
0.05 0.632 0 0.0 1e-06 
3.0 0.632 0 0.0 1e-06 
0.05 0.633 0 0.0 1e-06 
3.0 0.633 0 0.0 1e-06 
0.05 0.634 0 0.0 1e-06 
3.0 0.634 0 0.0 1e-06 
0.05 0.635 0 0.0 1e-06 
3.0 0.635 0 0.0 1e-06 
0.05 0.636 0 0.0 1e-06 
3.0 0.636 0 0.0 1e-06 
0.05 0.637 0 0.0 1e-06 
3.0 0.637 0 0.0 1e-06 
0.05 0.638 0 0.0 1e-06 
3.0 0.638 0 0.0 1e-06 
0.05 0.639 0 0.0 1e-06 
3.0 0.639 0 0.0 1e-06 
0.05 0.64 0 0.0 1e-06 
3.0 0.64 0 0.0 1e-06 
0.05 0.641 0 0.0 1e-06 
3.0 0.641 0 0.0 1e-06 
0.05 0.642 0 0.0 1e-06 
3.0 0.642 0 0.0 1e-06 
0.05 0.643 0 0.0 1e-06 
3.0 0.643 0 0.0 1e-06 
0.05 0.644 0 0.0 1e-06 
3.0 0.644 0 0.0 1e-06 
0.05 0.645 0 0.0 1e-06 
3.0 0.645 0 0.0 1e-06 
0.05 0.646 0 0.0 1e-06 
3.0 0.646 0 0.0 1e-06 
0.05 0.647 0 0.0 1e-06 
3.0 0.647 0 0.0 1e-06 
0.05 0.648 0 0.0 1e-06 
3.0 0.648 0 0.0 1e-06 
0.05 0.649 0 0.0 1e-06 
3.0 0.649 0 0.0 1e-06 
0.05 0.65 0 0.0 1e-06 
3.0 0.65 0 0.0 1e-06 
0.05 0.651 0 0.0 1e-06 
3.0 0.651 0 0.0 1e-06 
0.05 0.652 0 0.0 1e-06 
3.0 0.652 0 0.0 1e-06 
0.05 0.653 0 0.0 1e-06 
3.0 0.653 0 0.0 1e-06 
0.05 0.654 0 0.0 1e-06 
3.0 0.654 0 0.0 1e-06 
0.05 0.655 0 0.0 1e-06 
3.0 0.655 0 0.0 1e-06 
0.05 0.656 0 0.0 1e-06 
3.0 0.656 0 0.0 1e-06 
0.05 0.657 0 0.0 1e-06 
3.0 0.657 0 0.0 1e-06 
0.05 0.658 0 0.0 1e-06 
3.0 0.658 0 0.0 1e-06 
0.05 0.659 0 0.0 1e-06 
3.0 0.659 0 0.0 1e-06 
0.05 0.66 0 0.0 1e-06 
3.0 0.66 0 0.0 1e-06 
0.05 0.661 0 0.0 1e-06 
3.0 0.661 0 0.0 1e-06 
0.05 0.662 0 0.0 1e-06 
3.0 0.662 0 0.0 1e-06 
0.05 0.663 0 0.0 1e-06 
3.0 0.663 0 0.0 1e-06 
0.05 0.664 0 0.0 1e-06 
3.0 0.664 0 0.0 1e-06 
0.05 0.665 0 0.0 1e-06 
3.0 0.665 0 0.0 1e-06 
0.05 0.666 0 0.0 1e-06 
3.0 0.666 0 0.0 1e-06 
0.05 0.667 0 0.0 1e-06 
3.0 0.667 0 0.0 1e-06 
0.05 0.668 0 0.0 1e-06 
3.0 0.668 0 0.0 1e-06 
0.05 0.669 0 0.0 1e-06 
3.0 0.669 0 0.0 1e-06 
0.05 0.67 0 0.0 1e-06 
3.0 0.67 0 0.0 1e-06 
0.05 0.671 0 0.0 1e-06 
3.0 0.671 0 0.0 1e-06 
0.05 0.672 0 0.0 1e-06 
3.0 0.672 0 0.0 1e-06 
0.05 0.673 0 0.0 1e-06 
3.0 0.673 0 0.0 1e-06 
0.05 0.674 0 0.0 1e-06 
3.0 0.674 0 0.0 1e-06 
0.05 0.675 0 0.0 1e-06 
3.0 0.675 0 0.0 1e-06 
0.05 0.676 0 0.0 1e-06 
3.0 0.676 0 0.0 1e-06 
0.05 0.677 0 0.0 1e-06 
3.0 0.677 0 0.0 1e-06 
0.05 0.678 0 0.0 1e-06 
3.0 0.678 0 0.0 1e-06 
0.05 0.679 0 0.0 1e-06 
3.0 0.679 0 0.0 1e-06 
0.05 0.68 0 0.0 1e-06 
3.0 0.68 0 0.0 1e-06 
0.05 0.681 0 0.0 1e-06 
3.0 0.681 0 0.0 1e-06 
0.05 0.682 0 0.0 1e-06 
3.0 0.682 0 0.0 1e-06 
0.05 0.683 0 0.0 1e-06 
3.0 0.683 0 0.0 1e-06 
0.05 0.684 0 0.0 1e-06 
3.0 0.684 0 0.0 1e-06 
0.05 0.685 0 0.0 1e-06 
3.0 0.685 0 0.0 1e-06 
0.05 0.686 0 0.0 1e-06 
3.0 0.686 0 0.0 1e-06 
0.05 0.687 0 0.0 1e-06 
3.0 0.687 0 0.0 1e-06 
0.05 0.688 0 0.0 1e-06 
3.0 0.688 0 0.0 1e-06 
0.05 0.689 0 0.0 1e-06 
3.0 0.689 0 0.0 1e-06 
0.05 0.69 0 0.0 1e-06 
3.0 0.69 0 0.0 1e-06 
0.05 0.691 0 0.0 1e-06 
3.0 0.691 0 0.0 1e-06 
0.05 0.692 0 0.0 1e-06 
3.0 0.692 0 0.0 1e-06 
0.05 0.693 0 0.0 1e-06 
3.0 0.693 0 0.0 1e-06 
0.05 0.694 0 0.0 1e-06 
3.0 0.694 0 0.0 1e-06 
0.05 0.695 0 0.0 1e-06 
3.0 0.695 0 0.0 1e-06 
0.05 0.696 0 0.0 1e-06 
3.0 0.696 0 0.0 1e-06 
0.05 0.697 0 0.0 1e-06 
3.0 0.697 0 0.0 1e-06 
0.05 0.698 0 0.0 1e-06 
3.0 0.698 0 0.0 1e-06 
0.05 0.699 0 0.0 1e-06 
3.0 0.699 0 0.0 1e-06 
0.05 0.7 0 0.0 1e-06 
3.0 0.7 0 0.0 1e-06 
0.05 0.701 0 0.0 1e-06 
3.0 0.701 0 0.0 1e-06 
0.05 0.702 0 0.0 1e-06 
3.0 0.702 0 0.0 1e-06 
0.05 0.703 0 0.0 1e-06 
3.0 0.703 0 0.0 1e-06 
0.05 0.704 0 0.0 1e-06 
3.0 0.704 0 0.0 1e-06 
0.05 0.705 0 0.0 1e-06 
3.0 0.705 0 0.0 1e-06 
0.05 0.706 0 0.0 1e-06 
3.0 0.706 0 0.0 1e-06 
0.05 0.707 0 0.0 1e-06 
3.0 0.707 0 0.0 1e-06 
0.05 0.708 0 0.0 1e-06 
3.0 0.708 0 0.0 1e-06 
0.05 0.709 0 0.0 1e-06 
3.0 0.709 0 0.0 1e-06 
0.05 0.71 0 0.0 1e-06 
3.0 0.71 0 0.0 1e-06 
0.05 0.711 0 0.0 1e-06 
3.0 0.711 0 0.0 1e-06 
0.05 0.712 0 0.0 1e-06 
3.0 0.712 0 0.0 1e-06 
0.05 0.713 0 0.0 1e-06 
3.0 0.713 0 0.0 1e-06 
0.05 0.714 0 0.0 1e-06 
3.0 0.714 0 0.0 1e-06 
0.05 0.715 0 0.0 1e-06 
3.0 0.715 0 0.0 1e-06 
0.05 0.716 0 0.0 1e-06 
3.0 0.716 0 0.0 1e-06 
0.05 0.717 0 0.0 1e-06 
3.0 0.717 0 0.0 1e-06 
0.05 0.718 0 0.0 1e-06 
3.0 0.718 0 0.0 1e-06 
0.05 0.719 0 0.0 1e-06 
3.0 0.719 0 0.0 1e-06 
0.05 0.72 0 0.0 1e-06 
3.0 0.72 0 0.0 1e-06 
0.05 0.721 0 0.0 1e-06 
3.0 0.721 0 0.0 1e-06 
0.05 0.722 0 0.0 1e-06 
3.0 0.722 0 0.0 1e-06 
0.05 0.723 0 0.0 1e-06 
3.0 0.723 0 0.0 1e-06 
0.05 0.724 0 0.0 1e-06 
3.0 0.724 0 0.0 1e-06 
0.05 0.725 0 0.0 1e-06 
3.0 0.725 0 0.0 1e-06 
0.05 0.726 0 0.0 1e-06 
3.0 0.726 0 0.0 1e-06 
0.05 0.727 0 0.0 1e-06 
3.0 0.727 0 0.0 1e-06 
0.05 0.728 0 0.0 1e-06 
3.0 0.728 0 0.0 1e-06 
0.05 0.729 0 0.0 1e-06 
3.0 0.729 0 0.0 1e-06 
0.05 0.73 0 0.0 1e-06 
3.0 0.73 0 0.0 1e-06 
0.05 0.731 0 0.0 1e-06 
3.0 0.731 0 0.0 1e-06 
0.05 0.732 0 0.0 1e-06 
3.0 0.732 0 0.0 1e-06 
0.05 0.733 0 0.0 1e-06 
3.0 0.733 0 0.0 1e-06 
0.05 0.734 0 0.0 1e-06 
3.0 0.734 0 0.0 1e-06 
0.05 0.735 0 0.0 1e-06 
3.0 0.735 0 0.0 1e-06 
0.05 0.736 0 0.0 1e-06 
3.0 0.736 0 0.0 1e-06 
0.05 0.737 0 0.0 1e-06 
3.0 0.737 0 0.0 1e-06 
0.05 0.738 0 0.0 1e-06 
3.0 0.738 0 0.0 1e-06 
0.05 0.739 0 0.0 1e-06 
3.0 0.739 0 0.0 1e-06 
0.05 0.74 0 0.0 1e-06 
3.0 0.74 0 0.0 1e-06 
0.05 0.741 0 0.0 1e-06 
3.0 0.741 0 0.0 1e-06 
0.05 0.742 0 0.0 1e-06 
3.0 0.742 0 0.0 1e-06 
0.05 0.743 0 0.0 1e-06 
3.0 0.743 0 0.0 1e-06 
0.05 0.744 0 0.0 1e-06 
3.0 0.744 0 0.0 1e-06 
0.05 0.745 0 0.0 1e-06 
3.0 0.745 0 0.0 1e-06 
0.05 0.746 0 0.0 1e-06 
3.0 0.746 0 0.0 1e-06 
0.05 0.747 0 0.0 1e-06 
3.0 0.747 0 0.0 1e-06 
0.05 0.748 0 0.0 1e-06 
3.0 0.748 0 0.0 1e-06 
0.05 0.749 0 0.0 1e-06 
3.0 0.749 0 0.0 1e-06 
0.05 0.75 0 0.0 1e-06 
3.0 0.75 0 0.0 1e-06 
0.05 0.751 0 0.0 1e-06 
3.0 0.751 0 0.0 1e-06 
0.05 0.752 0 0.0 1e-06 
3.0 0.752 0 0.0 1e-06 
0.05 0.753 0 0.0 1e-06 
3.0 0.753 0 0.0 1e-06 
0.05 0.754 0 0.0 1e-06 
3.0 0.754 0 0.0 1e-06 
0.05 0.755 0 0.0 1e-06 
3.0 0.755 0 0.0 1e-06 
0.05 0.756 0 0.0 1e-06 
3.0 0.756 0 0.0 1e-06 
0.05 0.757 0 0.0 1e-06 
3.0 0.757 0 0.0 1e-06 
0.05 0.758 0 0.0 1e-06 
3.0 0.758 0 0.0 1e-06 
0.05 0.759 0 0.0 1e-06 
3.0 0.759 0 0.0 1e-06 
0.05 0.76 0 0.0 1e-06 
3.0 0.76 0 0.0 1e-06 
0.05 0.761 0 0.0 1e-06 
3.0 0.761 0 0.0 1e-06 
0.05 0.762 0 0.0 1e-06 
3.0 0.762 0 0.0 1e-06 
0.05 0.763 0 0.0 1e-06 
3.0 0.763 0 0.0 1e-06 
0.05 0.764 0 0.0 1e-06 
3.0 0.764 0 0.0 1e-06 
0.05 0.765 0 0.0 1e-06 
3.0 0.765 0 0.0 1e-06 
0.05 0.766 0 0.0 1e-06 
3.0 0.766 0 0.0 1e-06 
0.05 0.767 0 0.0 1e-06 
3.0 0.767 0 0.0 1e-06 
0.05 0.768 0 0.0 1e-06 
3.0 0.768 0 0.0 1e-06 
0.05 0.769 0 0.0 1e-06 
3.0 0.769 0 0.0 1e-06 
0.05 0.77 0 0.0 1e-06 
3.0 0.77 0 0.0 1e-06 
0.05 0.771 0 0.0 1e-06 
3.0 0.771 0 0.0 1e-06 
0.05 0.772 0 0.0 1e-06 
3.0 0.772 0 0.0 1e-06 
0.05 0.773 0 0.0 1e-06 
3.0 0.773 0 0.0 1e-06 
0.05 0.774 0 0.0 1e-06 
3.0 0.774 0 0.0 1e-06 
0.05 0.775 0 0.0 1e-06 
3.0 0.775 0 0.0 1e-06 
0.05 0.776 0 0.0 1e-06 
3.0 0.776 0 0.0 1e-06 
0.05 0.777 0 0.0 1e-06 
3.0 0.777 0 0.0 1e-06 
0.05 0.778 0 0.0 1e-06 
3.0 0.778 0 0.0 1e-06 
0.05 0.779 0 0.0 1e-06 
3.0 0.779 0 0.0 1e-06 
0.05 0.78 0 0.0 1e-06 
3.0 0.78 0 0.0 1e-06 
0.05 0.781 0 0.0 1e-06 
3.0 0.781 0 0.0 1e-06 
0.05 0.782 0 0.0 1e-06 
3.0 0.782 0 0.0 1e-06 
0.05 0.783 0 0.0 1e-06 
3.0 0.783 0 0.0 1e-06 
0.05 0.784 0 0.0 1e-06 
3.0 0.784 0 0.0 1e-06 
0.05 0.785 0 0.0 1e-06 
3.0 0.785 0 0.0 1e-06 
0.05 0.786 0 0.0 1e-06 
3.0 0.786 0 0.0 1e-06 
0.05 0.787 0 0.0 1e-06 
3.0 0.787 0 0.0 1e-06 
0.05 0.788 0 0.0 1e-06 
3.0 0.788 0 0.0 1e-06 
0.05 0.789 0 0.0 1e-06 
3.0 0.789 0 0.0 1e-06 
0.05 0.79 0 0.0 1e-06 
3.0 0.79 0 0.0 1e-06 
0.05 0.791 0 0.0 1e-06 
3.0 0.791 0 0.0 1e-06 
0.05 0.792 0 0.0 1e-06 
3.0 0.792 0 0.0 1e-06 
0.05 0.793 0 0.0 1e-06 
3.0 0.793 0 0.0 1e-06 
0.05 0.794 0 0.0 1e-06 
3.0 0.794 0 0.0 1e-06 
0.05 0.795 0 0.0 1e-06 
3.0 0.795 0 0.0 1e-06 
0.05 0.796 0 0.0 1e-06 
3.0 0.796 0 0.0 1e-06 
0.05 0.797 0 0.0 1e-06 
3.0 0.797 0 0.0 1e-06 
0.05 0.798 0 0.0 1e-06 
3.0 0.798 0 0.0 1e-06 
0.05 0.799 0 0.0 1e-06 
3.0 0.799 0 0.0 1e-06 
0.05 0.8 0 0.0 1e-06 
3.0 0.8 0 0.0 1e-06 
0.05 0.801 0 0.0 1e-06 
3.0 0.801 0 0.0 1e-06 
0.05 0.802 0 0.0 1e-06 
3.0 0.802 0 0.0 1e-06 
0.05 0.803 0 0.0 1e-06 
3.0 0.803 0 0.0 1e-06 
0.05 0.804 0 0.0 1e-06 
3.0 0.804 0 0.0 1e-06 
0.05 0.805 0 0.0 1e-06 
3.0 0.805 0 0.0 1e-06 
0.05 0.806 0 0.0 1e-06 
3.0 0.806 0 0.0 1e-06 
0.05 0.807 0 0.0 1e-06 
3.0 0.807 0 0.0 1e-06 
0.05 0.808 0 0.0 1e-06 
3.0 0.808 0 0.0 1e-06 
0.05 0.809 0 0.0 1e-06 
3.0 0.809 0 0.0 1e-06 
0.05 0.81 0 0.0 1e-06 
3.0 0.81 0 0.0 1e-06 
0.05 0.811 0 0.0 1e-06 
3.0 0.811 0 0.0 1e-06 
0.05 0.812 0 0.0 1e-06 
3.0 0.812 0 0.0 1e-06 
0.05 0.813 0 0.0 1e-06 
3.0 0.813 0 0.0 1e-06 
0.05 0.814 0 0.0 1e-06 
3.0 0.814 0 0.0 1e-06 
0.05 0.815 0 0.0 1e-06 
3.0 0.815 0 0.0 1e-06 
0.05 0.816 0 0.0 1e-06 
3.0 0.816 0 0.0 1e-06 
0.05 0.817 0 0.0 1e-06 
3.0 0.817 0 0.0 1e-06 
0.05 0.818 0 0.0 1e-06 
3.0 0.818 0 0.0 1e-06 
0.05 0.819 0 0.0 1e-06 
3.0 0.819 0 0.0 1e-06 
0.05 0.82 0 0.0 1e-06 
3.0 0.82 0 0.0 1e-06 
0.05 0.821 0 0.0 1e-06 
3.0 0.821 0 0.0 1e-06 
0.05 0.822 0 0.0 1e-06 
3.0 0.822 0 0.0 1e-06 
0.05 0.823 0 0.0 1e-06 
3.0 0.823 0 0.0 1e-06 
0.05 0.824 0 0.0 1e-06 
3.0 0.824 0 0.0 1e-06 
0.05 0.825 0 0.0 1e-06 
3.0 0.825 0 0.0 1e-06 
0.05 0.826 0 0.0 1e-06 
3.0 0.826 0 0.0 1e-06 
0.05 0.827 0 0.0 1e-06 
3.0 0.827 0 0.0 1e-06 
0.05 0.828 0 0.0 1e-06 
3.0 0.828 0 0.0 1e-06 
0.05 0.829 0 0.0 1e-06 
3.0 0.829 0 0.0 1e-06 
0.05 0.83 0 0.0 1e-06 
3.0 0.83 0 0.0 1e-06 
0.05 0.831 0 0.0 1e-06 
3.0 0.831 0 0.0 1e-06 
0.05 0.832 0 0.0 1e-06 
3.0 0.832 0 0.0 1e-06 
0.05 0.833 0 0.0 1e-06 
3.0 0.833 0 0.0 1e-06 
0.05 0.834 0 0.0 1e-06 
3.0 0.834 0 0.0 1e-06 
0.05 0.835 0 0.0 1e-06 
3.0 0.835 0 0.0 1e-06 
0.05 0.836 0 0.0 1e-06 
3.0 0.836 0 0.0 1e-06 
0.05 0.837 0 0.0 1e-06 
3.0 0.837 0 0.0 1e-06 
0.05 0.838 0 0.0 1e-06 
3.0 0.838 0 0.0 1e-06 
0.05 0.839 0 0.0 1e-06 
3.0 0.839 0 0.0 1e-06 
0.05 0.84 0 0.0 1e-06 
3.0 0.84 0 0.0 1e-06 
0.05 0.841 0 0.0 1e-06 
3.0 0.841 0 0.0 1e-06 
0.05 0.842 0 0.0 1e-06 
3.0 0.842 0 0.0 1e-06 
0.05 0.843 0 0.0 1e-06 
3.0 0.843 0 0.0 1e-06 
0.05 0.844 0 0.0 1e-06 
3.0 0.844 0 0.0 1e-06 
0.05 0.845 0 0.0 1e-06 
3.0 0.845 0 0.0 1e-06 
0.05 0.846 0 0.0 1e-06 
3.0 0.846 0 0.0 1e-06 
0.05 0.847 0 0.0 1e-06 
3.0 0.847 0 0.0 1e-06 
0.05 0.848 0 0.0 1e-06 
3.0 0.848 0 0.0 1e-06 
0.05 0.849 0 0.0 1e-06 
3.0 0.849 0 0.0 1e-06 
0.05 0.85 0 0.0 1e-06 
3.0 0.85 0 0.0 1e-06 
0.05 0.851 0 0.0 1e-06 
3.0 0.851 0 0.0 1e-06 
0.05 0.852 0 0.0 1e-06 
3.0 0.852 0 0.0 1e-06 
0.05 0.853 0 0.0 1e-06 
3.0 0.853 0 0.0 1e-06 
0.05 0.854 0 0.0 1e-06 
3.0 0.854 0 0.0 1e-06 
0.05 0.855 0 0.0 1e-06 
3.0 0.855 0 0.0 1e-06 
0.05 0.856 0 0.0 1e-06 
3.0 0.856 0 0.0 1e-06 
0.05 0.857 0 0.0 1e-06 
3.0 0.857 0 0.0 1e-06 
0.05 0.858 0 0.0 1e-06 
3.0 0.858 0 0.0 1e-06 
0.05 0.859 0 0.0 1e-06 
3.0 0.859 0 0.0 1e-06 
0.05 0.86 0 0.0 1e-06 
3.0 0.86 0 0.0 1e-06 
0.05 0.861 0 0.0 1e-06 
3.0 0.861 0 0.0 1e-06 
0.05 0.862 0 0.0 1e-06 
3.0 0.862 0 0.0 1e-06 
0.05 0.863 0 0.0 1e-06 
3.0 0.863 0 0.0 1e-06 
0.05 0.864 0 0.0 1e-06 
3.0 0.864 0 0.0 1e-06 
0.05 0.865 0 0.0 1e-06 
3.0 0.865 0 0.0 1e-06 
0.05 0.866 0 0.0 1e-06 
3.0 0.866 0 0.0 1e-06 
0.05 0.867 0 0.0 1e-06 
3.0 0.867 0 0.0 1e-06 
0.05 0.868 0 0.0 1e-06 
3.0 0.868 0 0.0 1e-06 
0.05 0.869 0 0.0 1e-06 
3.0 0.869 0 0.0 1e-06 
0.05 0.87 0 0.0 1e-06 
3.0 0.87 0 0.0 1e-06 
0.05 0.871 0 0.0 1e-06 
3.0 0.871 0 0.0 1e-06 
0.05 0.872 0 0.0 1e-06 
3.0 0.872 0 0.0 1e-06 
0.05 0.873 0 0.0 1e-06 
3.0 0.873 0 0.0 1e-06 
0.05 0.874 0 0.0 1e-06 
3.0 0.874 0 0.0 1e-06 
0.05 0.875 0 0.0 1e-06 
3.0 0.875 0 0.0 1e-06 
0.05 0.876 0 0.0 1e-06 
3.0 0.876 0 0.0 1e-06 
0.05 0.877 0 0.0 1e-06 
3.0 0.877 0 0.0 1e-06 
0.05 0.878 0 0.0 1e-06 
3.0 0.878 0 0.0 1e-06 
0.05 0.879 0 0.0 1e-06 
3.0 0.879 0 0.0 1e-06 
0.05 0.88 0 0.0 1e-06 
3.0 0.88 0 0.0 1e-06 
0.05 0.881 0 0.0 1e-06 
3.0 0.881 0 0.0 1e-06 
0.05 0.882 0 0.0 1e-06 
3.0 0.882 0 0.0 1e-06 
0.05 0.883 0 0.0 1e-06 
3.0 0.883 0 0.0 1e-06 
0.05 0.884 0 0.0 1e-06 
3.0 0.884 0 0.0 1e-06 
0.05 0.885 0 0.0 1e-06 
3.0 0.885 0 0.0 1e-06 
0.05 0.886 0 0.0 1e-06 
3.0 0.886 0 0.0 1e-06 
0.05 0.887 0 0.0 1e-06 
3.0 0.887 0 0.0 1e-06 
0.05 0.888 0 0.0 1e-06 
3.0 0.888 0 0.0 1e-06 
0.05 0.889 0 0.0 1e-06 
3.0 0.889 0 0.0 1e-06 
0.05 0.89 0 0.0 1e-06 
3.0 0.89 0 0.0 1e-06 
0.05 0.891 0 0.0 1e-06 
3.0 0.891 0 0.0 1e-06 
0.05 0.892 0 0.0 1e-06 
3.0 0.892 0 0.0 1e-06 
0.05 0.893 0 0.0 1e-06 
3.0 0.893 0 0.0 1e-06 
0.05 0.894 0 0.0 1e-06 
3.0 0.894 0 0.0 1e-06 
0.05 0.895 0 0.0 1e-06 
3.0 0.895 0 0.0 1e-06 
0.05 0.896 0 0.0 1e-06 
3.0 0.896 0 0.0 1e-06 
0.05 0.897 0 0.0 1e-06 
3.0 0.897 0 0.0 1e-06 
0.05 0.898 0 0.0 1e-06 
3.0 0.898 0 0.0 1e-06 
0.05 0.899 0 0.0 1e-06 
3.0 0.899 0 0.0 1e-06 
0.05 0.9 0 0.0 1e-06 
3.0 0.9 0 0.0 1e-06 
0.05 0.901 0 0.0 1e-06 
3.0 0.901 0 0.0 1e-06 
0.05 0.902 0 0.0 1e-06 
3.0 0.902 0 0.0 1e-06 
0.05 0.903 0 0.0 1e-06 
3.0 0.903 0 0.0 1e-06 
0.05 0.904 0 0.0 1e-06 
3.0 0.904 0 0.0 1e-06 
0.05 0.905 0 0.0 1e-06 
3.0 0.905 0 0.0 1e-06 
0.05 0.906 0 0.0 1e-06 
3.0 0.906 0 0.0 1e-06 
0.05 0.907 0 0.0 1e-06 
3.0 0.907 0 0.0 1e-06 
0.05 0.908 0 0.0 1e-06 
3.0 0.908 0 0.0 1e-06 
0.05 0.909 0 0.0 1e-06 
3.0 0.909 0 0.0 1e-06 
0.05 0.91 0 0.0 1e-06 
3.0 0.91 0 0.0 1e-06 
0.05 0.911 0 0.0 1e-06 
3.0 0.911 0 0.0 1e-06 
0.05 0.912 0 0.0 1e-06 
3.0 0.912 0 0.0 1e-06 
0.05 0.913 0 0.0 1e-06 
3.0 0.913 0 0.0 1e-06 
0.05 0.914 0 0.0 1e-06 
3.0 0.914 0 0.0 1e-06 
0.05 0.915 0 0.0 1e-06 
3.0 0.915 0 0.0 1e-06 
0.05 0.916 0 0.0 1e-06 
3.0 0.916 0 0.0 1e-06 
0.05 0.917 0 0.0 1e-06 
3.0 0.917 0 0.0 1e-06 
0.05 0.918 0 0.0 1e-06 
3.0 0.918 0 0.0 1e-06 
0.05 0.919 0 0.0 1e-06 
3.0 0.919 0 0.0 1e-06 
0.05 0.92 0 0.0 1e-06 
3.0 0.92 0 0.0 1e-06 
0.05 0.921 0 0.0 1e-06 
3.0 0.921 0 0.0 1e-06 
0.05 0.922 0 0.0 1e-06 
3.0 0.922 0 0.0 1e-06 
0.05 0.923 0 0.0 1e-06 
3.0 0.923 0 0.0 1e-06 
0.05 0.924 0 0.0 1e-06 
3.0 0.924 0 0.0 1e-06 
0.05 0.925 0 0.0 1e-06 
3.0 0.925 0 0.0 1e-06 
0.05 0.926 0 0.0 1e-06 
3.0 0.926 0 0.0 1e-06 
0.05 0.927 0 0.0 1e-06 
3.0 0.927 0 0.0 1e-06 
0.05 0.928 0 0.0 1e-06 
3.0 0.928 0 0.0 1e-06 
0.05 0.929 0 0.0 1e-06 
3.0 0.929 0 0.0 1e-06 
0.05 0.93 0 0.0 1e-06 
3.0 0.93 0 0.0 1e-06 
0.05 0.931 0 0.0 1e-06 
3.0 0.931 0 0.0 1e-06 
0.05 0.932 0 0.0 1e-06 
3.0 0.932 0 0.0 1e-06 
0.05 0.933 0 0.0 1e-06 
3.0 0.933 0 0.0 1e-06 
0.05 0.934 0 0.0 1e-06 
3.0 0.934 0 0.0 1e-06 
0.05 0.935 0 0.0 1e-06 
3.0 0.935 0 0.0 1e-06 
0.05 0.936 0 0.0 1e-06 
3.0 0.936 0 0.0 1e-06 
0.05 0.937 0 0.0 1e-06 
3.0 0.937 0 0.0 1e-06 
0.05 0.938 0 0.0 1e-06 
3.0 0.938 0 0.0 1e-06 
0.05 0.939 0 0.0 1e-06 
3.0 0.939 0 0.0 1e-06 
0.05 0.94 0 0.0 1e-06 
3.0 0.94 0 0.0 1e-06 
0.05 0.941 0 0.0 1e-06 
3.0 0.941 0 0.0 1e-06 
0.05 0.942 0 0.0 1e-06 
3.0 0.942 0 0.0 1e-06 
0.05 0.943 0 0.0 1e-06 
3.0 0.943 0 0.0 1e-06 
0.05 0.944 0 0.0 1e-06 
3.0 0.944 0 0.0 1e-06 
0.05 0.945 0 0.0 1e-06 
3.0 0.945 0 0.0 1e-06 
0.05 0.946 0 0.0 1e-06 
3.0 0.946 0 0.0 1e-06 
0.05 0.947 0 0.0 1e-06 
3.0 0.947 0 0.0 1e-06 
0.05 0.948 0 0.0 1e-06 
3.0 0.948 0 0.0 1e-06 
0.05 0.949 0 0.0 1e-06 
3.0 0.949 0 0.0 1e-06 
0.05 0.95 0 0.0 1e-06 
3.0 0.95 0 0.0 1e-06 
0.05 0.951 0 0.0 1e-06 
3.0 0.951 0 0.0 1e-06 
0.05 0.952 0 0.0 1e-06 
3.0 0.952 0 0.0 1e-06 
0.05 0.953 0 0.0 1e-06 
3.0 0.953 0 0.0 1e-06 
0.05 0.954 0 0.0 1e-06 
3.0 0.954 0 0.0 1e-06 
0.05 0.955 0 0.0 1e-06 
3.0 0.955 0 0.0 1e-06 
0.05 0.956 0 0.0 1e-06 
3.0 0.956 0 0.0 1e-06 
0.05 0.957 0 0.0 1e-06 
3.0 0.957 0 0.0 1e-06 
0.05 0.958 0 0.0 1e-06 
3.0 0.958 0 0.0 1e-06 
0.05 0.959 0 0.0 1e-06 
3.0 0.959 0 0.0 1e-06 
0.05 0.96 0 0.0 1e-06 
3.0 0.96 0 0.0 1e-06 
0.05 0.961 0 0.0 1e-06 
3.0 0.961 0 0.0 1e-06 
0.05 0.962 0 0.0 1e-06 
3.0 0.962 0 0.0 1e-06 
0.05 0.963 0 0.0 1e-06 
3.0 0.963 0 0.0 1e-06 
0.05 0.964 0 0.0 1e-06 
3.0 0.964 0 0.0 1e-06 
0.05 0.965 0 0.0 1e-06 
3.0 0.965 0 0.0 1e-06 
0.05 0.966 0 0.0 1e-06 
3.0 0.966 0 0.0 1e-06 
0.05 0.967 0 0.0 1e-06 
3.0 0.967 0 0.0 1e-06 
0.05 0.968 0 0.0 1e-06 
3.0 0.968 0 0.0 1e-06 
0.05 0.969 0 0.0 1e-06 
3.0 0.969 0 0.0 1e-06 
0.05 0.97 0 0.0 1e-06 
3.0 0.97 0 0.0 1e-06 
0.05 0.971 0 0.0 1e-06 
3.0 0.971 0 0.0 1e-06 
0.05 0.972 0 0.0 1e-06 
3.0 0.972 0 0.0 1e-06 
0.05 0.973 0 0.0 1e-06 
3.0 0.973 0 0.0 1e-06 
0.05 0.974 0 0.0 1e-06 
3.0 0.974 0 0.0 1e-06 
0.05 0.975 0 0.0 1e-06 
3.0 0.975 0 0.0 1e-06 
0.05 0.976 0 0.0 1e-06 
3.0 0.976 0 0.0 1e-06 
0.05 0.977 0 0.0 1e-06 
3.0 0.977 0 0.0 1e-06 
0.05 0.978 0 0.0 1e-06 
3.0 0.978 0 0.0 1e-06 
0.05 0.979 0 0.0 1e-06 
3.0 0.979 0 0.0 1e-06 
0.05 0.98 0 0.0 1e-06 
3.0 0.98 0 0.0 1e-06 
0.05 0.981 0 0.0 1e-06 
3.0 0.981 0 0.0 1e-06 
0.05 0.982 0 0.0 1e-06 
3.0 0.982 0 0.0 1e-06 
0.05 0.983 0 0.0 1e-06 
3.0 0.983 0 0.0 1e-06 
0.05 0.984 0 0.0 1e-06 
3.0 0.984 0 0.0 1e-06 
0.05 0.985 0 0.0 1e-06 
3.0 0.985 0 0.0 1e-06 
0.05 0.986 0 0.0 1e-06 
3.0 0.986 0 0.0 1e-06 
0.05 0.987 0 0.0 1e-06 
3.0 0.987 0 0.0 1e-06 
0.05 0.988 0 0.0 1e-06 
3.0 0.988 0 0.0 1e-06 
0.05 0.989 0 0.0 1e-06 
3.0 0.989 0 0.0 1e-06 
0.05 0.99 0 0.0 1e-06 
3.0 0.99 0 0.0 1e-06 
0.05 0.991 0 0.0 1e-06 
3.0 0.991 0 0.0 1e-06 
0.05 0.992 0 0.0 1e-06 
3.0 0.992 0 0.0 1e-06 
0.05 0.993 0 0.0 1e-06 
3.0 0.993 0 0.0 1e-06 
0.05 0.994 0 0.0 1e-06 
3.0 0.994 0 0.0 1e-06 
0.05 0.995 0 0.0 1e-06 
3.0 0.995 0 0.0 1e-06 
0.05 0.996 0 0.0 1e-06 
3.0 0.996 0 0.0 1e-06 
0.05 0.997 0 0.0 1e-06 
3.0 0.997 0 0.0 1e-06 
0.05 0.998 0 0.0 1e-06 
3.0 0.998 0 0.0 1e-06 
0.05 0.999 0 0.0 1e-06 
3.0 0.999 0 0.0 1e-06 
0.05 1.0 0 0.0 1e-06 
3.0 1.0 0 0.0 1e-06 
0.05 1.001 0 0.0 1e-06 
3.0 1.001 0 0.0 1e-06 
0.05 1.002 0 0.0 1e-06 
3.0 1.002 0 0.0 1e-06 
0.05 1.003 0 0.0 1e-06 
3.0 1.003 0 0.0 1e-06 
0.05 1.004 0 0.0 1e-06 
3.0 1.004 0 0.0 1e-06 
0.05 1.005 0 0.0 1e-06 
3.0 1.005 0 0.0 1e-06 
0.05 1.006 0 0.0 1e-06 
3.0 1.006 0 0.0 1e-06 
0.05 1.007 0 0.0 1e-06 
3.0 1.007 0 0.0 1e-06 
0.05 1.008 0 0.0 1e-06 
3.0 1.008 0 0.0 1e-06 
0.05 1.009 0 0.0 1e-06 
3.0 1.009 0 0.0 1e-06 
0.05 1.01 0 0.0 1e-06 
3.0 1.01 0 0.0 1e-06 
0.05 1.011 0 0.0 1e-06 
3.0 1.011 0 0.0 1e-06 
0.05 1.012 0 0.0 1e-06 
3.0 1.012 0 0.0 1e-06 
0.05 1.013 0 0.0 1e-06 
3.0 1.013 0 0.0 1e-06 
0.05 1.014 0 0.0 1e-06 
3.0 1.014 0 0.0 1e-06 
0.05 1.015 0 0.0 1e-06 
3.0 1.015 0 0.0 1e-06 
0.05 1.016 0 0.0 1e-06 
3.0 1.016 0 0.0 1e-06 
0.05 1.017 0 0.0 1e-06 
3.0 1.017 0 0.0 1e-06 
0.05 1.018 0 0.0 1e-06 
3.0 1.018 0 0.0 1e-06 
0.05 1.019 0 0.0 1e-06 
3.0 1.019 0 0.0 1e-06 
0.05 1.02 0 0.0 1e-06 
3.0 1.02 0 0.0 1e-06 
0.05 1.021 0 0.0 1e-06 
3.0 1.021 0 0.0 1e-06 
0.05 1.022 0 0.0 1e-06 
3.0 1.022 0 0.0 1e-06 
0.05 1.023 0 0.0 1e-06 
3.0 1.023 0 0.0 1e-06 
0.05 1.024 0 0.0 1e-06 
3.0 1.024 0 0.0 1e-06 
0.05 1.025 0 0.0 1e-06 
3.0 1.025 0 0.0 1e-06 
0.05 1.026 0 0.0 1e-06 
3.0 1.026 0 0.0 1e-06 
0.05 1.027 0 0.0 1e-06 
3.0 1.027 0 0.0 1e-06 
0.05 1.028 0 0.0 1e-06 
3.0 1.028 0 0.0 1e-06 
0.05 1.029 0 0.0 1e-06 
3.0 1.029 0 0.0 1e-06 
0.05 1.03 0 0.0 1e-06 
3.0 1.03 0 0.0 1e-06 
0.05 1.031 0 0.0 1e-06 
3.0 1.031 0 0.0 1e-06 
0.05 1.032 0 0.0 1e-06 
3.0 1.032 0 0.0 1e-06 
0.05 1.033 0 0.0 1e-06 
3.0 1.033 0 0.0 1e-06 
0.05 1.034 0 0.0 1e-06 
3.0 1.034 0 0.0 1e-06 
0.05 1.035 0 0.0 1e-06 
3.0 1.035 0 0.0 1e-06 
0.05 1.036 0 0.0 1e-06 
3.0 1.036 0 0.0 1e-06 
0.05 1.037 0 0.0 1e-06 
3.0 1.037 0 0.0 1e-06 
0.05 1.038 0 0.0 1e-06 
3.0 1.038 0 0.0 1e-06 
0.05 1.039 0 0.0 1e-06 
3.0 1.039 0 0.0 1e-06 
0.05 1.04 0 0.0 1e-06 
3.0 1.04 0 0.0 1e-06 
0.05 1.041 0 0.0 1e-06 
3.0 1.041 0 0.0 1e-06 
0.05 1.042 0 0.0 1e-06 
3.0 1.042 0 0.0 1e-06 
0.05 1.043 0 0.0 1e-06 
3.0 1.043 0 0.0 1e-06 
0.05 1.044 0 0.0 1e-06 
3.0 1.044 0 0.0 1e-06 
0.05 1.045 0 0.0 1e-06 
3.0 1.045 0 0.0 1e-06 
0.05 1.046 0 0.0 1e-06 
3.0 1.046 0 0.0 1e-06 
0.05 1.047 0 0.0 1e-06 
3.0 1.047 0 0.0 1e-06 
0.05 1.048 0 0.0 1e-06 
3.0 1.048 0 0.0 1e-06 
0.05 1.049 0 0.0 1e-06 
3.0 1.049 0 0.0 1e-06 
0.05 1.05 0 0.0 1e-06 
3.0 1.05 0 0.0 1e-06 
0.05 1.051 0 0.0 1e-06 
3.0 1.051 0 0.0 1e-06 
0.05 1.052 0 0.0 1e-06 
3.0 1.052 0 0.0 1e-06 
0.05 1.053 0 0.0 1e-06 
3.0 1.053 0 0.0 1e-06 
0.05 1.054 0 0.0 1e-06 
3.0 1.054 0 0.0 1e-06 
0.05 1.055 0 0.0 1e-06 
3.0 1.055 0 0.0 1e-06 
0.05 1.056 0 0.0 1e-06 
3.0 1.056 0 0.0 1e-06 
0.05 1.057 0 0.0 1e-06 
3.0 1.057 0 0.0 1e-06 
0.05 1.058 0 0.0 1e-06 
3.0 1.058 0 0.0 1e-06 
0.05 1.059 0 0.0 1e-06 
3.0 1.059 0 0.0 1e-06 
0.05 1.06 0 0.0 1e-06 
3.0 1.06 0 0.0 1e-06 
0.05 1.061 0 0.0 1e-06 
3.0 1.061 0 0.0 1e-06 
0.05 1.062 0 0.0 1e-06 
3.0 1.062 0 0.0 1e-06 
0.05 1.063 0 0.0 1e-06 
3.0 1.063 0 0.0 1e-06 
0.05 1.064 0 0.0 1e-06 
3.0 1.064 0 0.0 1e-06 
0.05 1.065 0 0.0 1e-06 
3.0 1.065 0 0.0 1e-06 
0.05 1.066 0 0.0 1e-06 
3.0 1.066 0 0.0 1e-06 
0.05 1.067 0 0.0 1e-06 
3.0 1.067 0 0.0 1e-06 
0.05 1.068 0 0.0 1e-06 
3.0 1.068 0 0.0 1e-06 
0.05 1.069 0 0.0 1e-06 
3.0 1.069 0 0.0 1e-06 
0.05 1.07 0 0.0 1e-06 
3.0 1.07 0 0.0 1e-06 
0.05 1.071 0 0.0 1e-06 
3.0 1.071 0 0.0 1e-06 
0.05 1.072 0 0.0 1e-06 
3.0 1.072 0 0.0 1e-06 
0.05 1.073 0 0.0 1e-06 
3.0 1.073 0 0.0 1e-06 
0.05 1.074 0 0.0 1e-06 
3.0 1.074 0 0.0 1e-06 
0.05 1.075 0 0.0 1e-06 
3.0 1.075 0 0.0 1e-06 
0.05 1.076 0 0.0 1e-06 
3.0 1.076 0 0.0 1e-06 
0.05 1.077 0 0.0 1e-06 
3.0 1.077 0 0.0 1e-06 
0.05 1.078 0 0.0 1e-06 
3.0 1.078 0 0.0 1e-06 
0.05 1.079 0 0.0 1e-06 
3.0 1.079 0 0.0 1e-06 
0.05 1.08 0 0.0 1e-06 
3.0 1.08 0 0.0 1e-06 
0.05 1.081 0 0.0 1e-06 
3.0 1.081 0 0.0 1e-06 
0.05 1.082 0 0.0 1e-06 
3.0 1.082 0 0.0 1e-06 
0.05 1.083 0 0.0 1e-06 
3.0 1.083 0 0.0 1e-06 
0.05 1.084 0 0.0 1e-06 
3.0 1.084 0 0.0 1e-06 
0.05 1.085 0 0.0 1e-06 
3.0 1.085 0 0.0 1e-06 
0.05 1.086 0 0.0 1e-06 
3.0 1.086 0 0.0 1e-06 
0.05 1.087 0 0.0 1e-06 
3.0 1.087 0 0.0 1e-06 
0.05 1.088 0 0.0 1e-06 
3.0 1.088 0 0.0 1e-06 
0.05 1.089 0 0.0 1e-06 
3.0 1.089 0 0.0 1e-06 
0.05 1.09 0 0.0 1e-06 
3.0 1.09 0 0.0 1e-06 
0.05 1.091 0 0.0 1e-06 
3.0 1.091 0 0.0 1e-06 
0.05 1.092 0 0.0 1e-06 
3.0 1.092 0 0.0 1e-06 
0.05 1.093 0 0.0 1e-06 
3.0 1.093 0 0.0 1e-06 
0.05 1.094 0 0.0 1e-06 
3.0 1.094 0 0.0 1e-06 
0.05 1.095 0 0.0 1e-06 
3.0 1.095 0 0.0 1e-06 
0.05 1.096 0 0.0 1e-06 
3.0 1.096 0 0.0 1e-06 
0.05 1.097 0 0.0 1e-06 
3.0 1.097 0 0.0 1e-06 
0.05 1.098 0 0.0 1e-06 
3.0 1.098 0 0.0 1e-06 
0.05 1.099 0 0.0 1e-06 
3.0 1.099 0 0.0 1e-06 
0.05 1.1 0 0.0 1e-06 
3.0 1.1 0 0.0 1e-06 
0.05 1.101 0 0.0 1e-06 
3.0 1.101 0 0.0 1e-06 
0.05 1.102 0 0.0 1e-06 
3.0 1.102 0 0.0 1e-06 
0.05 1.103 0 0.0 1e-06 
3.0 1.103 0 0.0 1e-06 
0.05 1.104 0 0.0 1e-06 
3.0 1.104 0 0.0 1e-06 
0.05 1.105 0 0.0 1e-06 
3.0 1.105 0 0.0 1e-06 
0.05 1.106 0 0.0 1e-06 
3.0 1.106 0 0.0 1e-06 
0.05 1.107 0 0.0 1e-06 
3.0 1.107 0 0.0 1e-06 
0.05 1.108 0 0.0 1e-06 
3.0 1.108 0 0.0 1e-06 
0.05 1.109 0 0.0 1e-06 
3.0 1.109 0 0.0 1e-06 
0.05 1.11 0 0.0 1e-06 
3.0 1.11 0 0.0 1e-06 
0.05 1.111 0 0.0 1e-06 
3.0 1.111 0 0.0 1e-06 
0.05 1.112 0 0.0 1e-06 
3.0 1.112 0 0.0 1e-06 
0.05 1.113 0 0.0 1e-06 
3.0 1.113 0 0.0 1e-06 
0.05 1.114 0 0.0 1e-06 
3.0 1.114 0 0.0 1e-06 
0.05 1.115 0 0.0 1e-06 
3.0 1.115 0 0.0 1e-06 
0.05 1.116 0 0.0 1e-06 
3.0 1.116 0 0.0 1e-06 
0.05 1.117 0 0.0 1e-06 
3.0 1.117 0 0.0 1e-06 
0.05 1.118 0 0.0 1e-06 
3.0 1.118 0 0.0 1e-06 
0.05 1.119 0 0.0 1e-06 
3.0 1.119 0 0.0 1e-06 
0.05 1.12 0 0.0 1e-06 
3.0 1.12 0 0.0 1e-06 
0.05 1.121 0 0.0 1e-06 
3.0 1.121 0 0.0 1e-06 
0.05 1.122 0 0.0 1e-06 
3.0 1.122 0 0.0 1e-06 
0.05 1.123 0 0.0 1e-06 
3.0 1.123 0 0.0 1e-06 
0.05 1.124 0 0.0 1e-06 
3.0 1.124 0 0.0 1e-06 
0.05 1.125 0 0.0 1e-06 
3.0 1.125 0 0.0 1e-06 
0.05 1.126 0 0.0 1e-06 
3.0 1.126 0 0.0 1e-06 
0.05 1.127 0 0.0 1e-06 
3.0 1.127 0 0.0 1e-06 
0.05 1.128 0 0.0 1e-06 
3.0 1.128 0 0.0 1e-06 
0.05 1.129 0 0.0 1e-06 
3.0 1.129 0 0.0 1e-06 
0.05 1.13 0 0.0 1e-06 
3.0 1.13 0 0.0 1e-06 
0.05 1.131 0 0.0 1e-06 
3.0 1.131 0 0.0 1e-06 
0.05 1.132 0 0.0 1e-06 
3.0 1.132 0 0.0 1e-06 
0.05 1.133 0 0.0 1e-06 
3.0 1.133 0 0.0 1e-06 
0.05 1.134 0 0.0 1e-06 
3.0 1.134 0 0.0 1e-06 
0.05 1.135 0 0.0 1e-06 
3.0 1.135 0 0.0 1e-06 
0.05 1.136 0 0.0 1e-06 
3.0 1.136 0 0.0 1e-06 
0.05 1.137 0 0.0 1e-06 
3.0 1.137 0 0.0 1e-06 
0.05 1.138 0 0.0 1e-06 
3.0 1.138 0 0.0 1e-06 
0.05 1.139 0 0.0 1e-06 
3.0 1.139 0 0.0 1e-06 
0.05 1.14 0 0.0 1e-06 
3.0 1.14 0 0.0 1e-06 
0.05 1.141 0 0.0 1e-06 
3.0 1.141 0 0.0 1e-06 
0.05 1.142 0 0.0 1e-06 
3.0 1.142 0 0.0 1e-06 
0.05 1.143 0 0.0 1e-06 
3.0 1.143 0 0.0 1e-06 
0.05 1.144 0 0.0 1e-06 
3.0 1.144 0 0.0 1e-06 
0.05 1.145 0 0.0 1e-06 
3.0 1.145 0 0.0 1e-06 
0.05 1.146 0 0.0 1e-06 
3.0 1.146 0 0.0 1e-06 
0.05 1.147 0 0.0 1e-06 
3.0 1.147 0 0.0 1e-06 
0.05 1.148 0 0.0 1e-06 
3.0 1.148 0 0.0 1e-06 
0.05 1.149 0 0.0 1e-06 
3.0 1.149 0 0.0 1e-06 
0.05 1.15 0 0.0 1e-06 
3.0 1.15 0 0.0 1e-06 
0.05 1.151 0 0.0 1e-06 
3.0 1.151 0 0.0 1e-06 
0.05 1.152 0 0.0 1e-06 
3.0 1.152 0 0.0 1e-06 
0.05 1.153 0 0.0 1e-06 
3.0 1.153 0 0.0 1e-06 
0.05 1.154 0 0.0 1e-06 
3.0 1.154 0 0.0 1e-06 
0.05 1.155 0 0.0 1e-06 
3.0 1.155 0 0.0 1e-06 
0.05 1.156 0 0.0 1e-06 
3.0 1.156 0 0.0 1e-06 
0.05 1.157 0 0.0 1e-06 
3.0 1.157 0 0.0 1e-06 
0.05 1.158 0 0.0 1e-06 
3.0 1.158 0 0.0 1e-06 
0.05 1.159 0 0.0 1e-06 
3.0 1.159 0 0.0 1e-06 
0.05 1.16 0 0.0 1e-06 
3.0 1.16 0 0.0 1e-06 
0.05 1.161 0 0.0 1e-06 
3.0 1.161 0 0.0 1e-06 
0.05 1.162 0 0.0 1e-06 
3.0 1.162 0 0.0 1e-06 
0.05 1.163 0 0.0 1e-06 
3.0 1.163 0 0.0 1e-06 
0.05 1.164 0 0.0 1e-06 
3.0 1.164 0 0.0 1e-06 
0.05 1.165 0 0.0 1e-06 
3.0 1.165 0 0.0 1e-06 
0.05 1.166 0 0.0 1e-06 
3.0 1.166 0 0.0 1e-06 
0.05 1.167 0 0.0 1e-06 
3.0 1.167 0 0.0 1e-06 
0.05 1.168 0 0.0 1e-06 
3.0 1.168 0 0.0 1e-06 
0.05 1.169 0 0.0 1e-06 
3.0 1.169 0 0.0 1e-06 
0.05 1.17 0 0.0 1e-06 
3.0 1.17 0 0.0 1e-06 
0.05 1.171 0 0.0 1e-06 
3.0 1.171 0 0.0 1e-06 
0.05 1.172 0 0.0 1e-06 
3.0 1.172 0 0.0 1e-06 
0.05 1.173 0 0.0 1e-06 
3.0 1.173 0 0.0 1e-06 
0.05 1.174 0 0.0 1e-06 
3.0 1.174 0 0.0 1e-06 
0.05 1.175 0 0.0 1e-06 
3.0 1.175 0 0.0 1e-06 
0.05 1.176 0 0.0 1e-06 
3.0 1.176 0 0.0 1e-06 
0.05 1.177 0 0.0 1e-06 
3.0 1.177 0 0.0 1e-06 
0.05 1.178 0 0.0 1e-06 
3.0 1.178 0 0.0 1e-06 
0.05 1.179 0 0.0 1e-06 
3.0 1.179 0 0.0 1e-06 
0.05 1.18 0 0.0 1e-06 
3.0 1.18 0 0.0 1e-06 
0.05 1.181 0 0.0 1e-06 
3.0 1.181 0 0.0 1e-06 
0.05 1.182 0 0.0 1e-06 
3.0 1.182 0 0.0 1e-06 
0.05 1.183 0 0.0 1e-06 
3.0 1.183 0 0.0 1e-06 
0.05 1.184 0 0.0 1e-06 
3.0 1.184 0 0.0 1e-06 
0.05 1.185 0 0.0 1e-06 
3.0 1.185 0 0.0 1e-06 
0.05 1.186 0 0.0 1e-06 
3.0 1.186 0 0.0 1e-06 
0.05 1.187 0 0.0 1e-06 
3.0 1.187 0 0.0 1e-06 
0.05 1.188 0 0.0 1e-06 
3.0 1.188 0 0.0 1e-06 
0.05 1.189 0 0.0 1e-06 
3.0 1.189 0 0.0 1e-06 
0.05 1.19 0 0.0 1e-06 
3.0 1.19 0 0.0 1e-06 
0.05 1.191 0 0.0 1e-06 
3.0 1.191 0 0.0 1e-06 
0.05 1.192 0 0.0 1e-06 
3.0 1.192 0 0.0 1e-06 
0.05 1.193 0 0.0 1e-06 
3.0 1.193 0 0.0 1e-06 
0.05 1.194 0 0.0 1e-06 
3.0 1.194 0 0.0 1e-06 
0.05 1.195 0 0.0 1e-06 
3.0 1.195 0 0.0 1e-06 
0.05 1.196 0 0.0 1e-06 
3.0 1.196 0 0.0 1e-06 
0.05 1.197 0 0.0 1e-06 
3.0 1.197 0 0.0 1e-06 
0.05 1.198 0 0.0 1e-06 
3.0 1.198 0 0.0 1e-06 
0.05 1.199 0 0.0 1e-06 
3.0 1.199 0 0.0 1e-06 
0.05 1.2 0 0.0 1e-06 
3.0 1.2 0 0.0 1e-06 
0.05 1.201 0 0.0 1e-06 
3.0 1.201 0 0.0 1e-06 
0.05 1.202 0 0.0 1e-06 
3.0 1.202 0 0.0 1e-06 
0.05 1.203 0 0.0 1e-06 
3.0 1.203 0 0.0 1e-06 
0.05 1.204 0 0.0 1e-06 
3.0 1.204 0 0.0 1e-06 
0.05 1.205 0 0.0 1e-06 
3.0 1.205 0 0.0 1e-06 
0.05 1.206 0 0.0 1e-06 
3.0 1.206 0 0.0 1e-06 
0.05 1.207 0 0.0 1e-06 
3.0 1.207 0 0.0 1e-06 
0.05 1.208 0 0.0 1e-06 
3.0 1.208 0 0.0 1e-06 
0.05 1.209 0 0.0 1e-06 
3.0 1.209 0 0.0 1e-06 
0.05 1.21 0 0.0 1e-06 
3.0 1.21 0 0.0 1e-06 
0.05 1.211 0 0.0 1e-06 
3.0 1.211 0 0.0 1e-06 
0.05 1.212 0 0.0 1e-06 
3.0 1.212 0 0.0 1e-06 
0.05 1.213 0 0.0 1e-06 
3.0 1.213 0 0.0 1e-06 
0.05 1.214 0 0.0 1e-06 
3.0 1.214 0 0.0 1e-06 
0.05 1.215 0 0.0 1e-06 
3.0 1.215 0 0.0 1e-06 
0.05 1.216 0 0.0 1e-06 
3.0 1.216 0 0.0 1e-06 
0.05 1.217 0 0.0 1e-06 
3.0 1.217 0 0.0 1e-06 
0.05 1.218 0 0.0 1e-06 
3.0 1.218 0 0.0 1e-06 
0.05 1.219 0 0.0 1e-06 
3.0 1.219 0 0.0 1e-06 
0.05 1.22 0 0.0 1e-06 
3.0 1.22 0 0.0 1e-06 
0.05 1.221 0 0.0 1e-06 
3.0 1.221 0 0.0 1e-06 
0.05 1.222 0 0.0 1e-06 
3.0 1.222 0 0.0 1e-06 
0.05 1.223 0 0.0 1e-06 
3.0 1.223 0 0.0 1e-06 
0.05 1.224 0 0.0 1e-06 
3.0 1.224 0 0.0 1e-06 
0.05 1.225 0 0.0 1e-06 
3.0 1.225 0 0.0 1e-06 
0.05 1.226 0 0.0 1e-06 
3.0 1.226 0 0.0 1e-06 
0.05 1.227 0 0.0 1e-06 
3.0 1.227 0 0.0 1e-06 
0.05 1.228 0 0.0 1e-06 
3.0 1.228 0 0.0 1e-06 
0.05 1.229 0 0.0 1e-06 
3.0 1.229 0 0.0 1e-06 
0.05 1.23 0 0.0 1e-06 
3.0 1.23 0 0.0 1e-06 
0.05 1.231 0 0.0 1e-06 
3.0 1.231 0 0.0 1e-06 
0.05 1.232 0 0.0 1e-06 
3.0 1.232 0 0.0 1e-06 
0.05 1.233 0 0.0 1e-06 
3.0 1.233 0 0.0 1e-06 
0.05 1.234 0 0.0 1e-06 
3.0 1.234 0 0.0 1e-06 
0.05 1.235 0 0.0 1e-06 
3.0 1.235 0 0.0 1e-06 
0.05 1.236 0 0.0 1e-06 
3.0 1.236 0 0.0 1e-06 
0.05 1.237 0 0.0 1e-06 
3.0 1.237 0 0.0 1e-06 
0.05 1.238 0 0.0 1e-06 
3.0 1.238 0 0.0 1e-06 
0.05 1.239 0 0.0 1e-06 
3.0 1.239 0 0.0 1e-06 
0.05 1.24 0 0.0 1e-06 
3.0 1.24 0 0.0 1e-06 
0.05 1.241 0 0.0 1e-06 
3.0 1.241 0 0.0 1e-06 
0.05 1.242 0 0.0 1e-06 
3.0 1.242 0 0.0 1e-06 
0.05 1.243 0 0.0 1e-06 
3.0 1.243 0 0.0 1e-06 
0.05 1.244 0 0.0 1e-06 
3.0 1.244 0 0.0 1e-06 
0.05 1.245 0 0.0 1e-06 
3.0 1.245 0 0.0 1e-06 
0.05 1.246 0 0.0 1e-06 
3.0 1.246 0 0.0 1e-06 
0.05 1.247 0 0.0 1e-06 
3.0 1.247 0 0.0 1e-06 
0.05 1.248 0 0.0 1e-06 
3.0 1.248 0 0.0 1e-06 
0.05 1.249 0 0.0 1e-06 
3.0 1.249 0 0.0 1e-06 
0.05 1.25 0 0.0 1e-06 
3.0 1.25 0 0.0 1e-06 
0.05 1.251 0 0.0 1e-06 
3.0 1.251 0 0.0 1e-06 
0.05 1.252 0 0.0 1e-06 
3.0 1.252 0 0.0 1e-06 
0.05 1.253 0 0.0 1e-06 
3.0 1.253 0 0.0 1e-06 
0.05 1.254 0 0.0 1e-06 
3.0 1.254 0 0.0 1e-06 
0.05 1.255 0 0.0 1e-06 
3.0 1.255 0 0.0 1e-06 
0.05 1.256 0 0.0 1e-06 
3.0 1.256 0 0.0 1e-06 
0.05 1.257 0 0.0 1e-06 
3.0 1.257 0 0.0 1e-06 
0.05 1.258 0 0.0 1e-06 
3.0 1.258 0 0.0 1e-06 
0.05 1.259 0 0.0 1e-06 
3.0 1.259 0 0.0 1e-06 
0.05 1.26 0 0.0 1e-06 
3.0 1.26 0 0.0 1e-06 
0.05 1.261 0 0.0 1e-06 
3.0 1.261 0 0.0 1e-06 
0.05 1.262 0 0.0 1e-06 
3.0 1.262 0 0.0 1e-06 
0.05 1.263 0 0.0 1e-06 
3.0 1.263 0 0.0 1e-06 
0.05 1.264 0 0.0 1e-06 
3.0 1.264 0 0.0 1e-06 
0.05 1.265 0 0.0 1e-06 
3.0 1.265 0 0.0 1e-06 
0.05 1.266 0 0.0 1e-06 
3.0 1.266 0 0.0 1e-06 
0.05 1.267 0 0.0 1e-06 
3.0 1.267 0 0.0 1e-06 
0.05 1.268 0 0.0 1e-06 
3.0 1.268 0 0.0 1e-06 
0.05 1.269 0 0.0 1e-06 
3.0 1.269 0 0.0 1e-06 
0.05 1.27 0 0.0 1e-06 
3.0 1.27 0 0.0 1e-06 
0.05 1.271 0 0.0 1e-06 
3.0 1.271 0 0.0 1e-06 
0.05 1.272 0 0.0 1e-06 
3.0 1.272 0 0.0 1e-06 
0.05 1.273 0 0.0 1e-06 
3.0 1.273 0 0.0 1e-06 
0.05 1.274 0 0.0 1e-06 
3.0 1.274 0 0.0 1e-06 
0.05 1.275 0 0.0 1e-06 
3.0 1.275 0 0.0 1e-06 
0.05 1.276 0 0.0 1e-06 
3.0 1.276 0 0.0 1e-06 
0.05 1.277 0 0.0 1e-06 
3.0 1.277 0 0.0 1e-06 
0.05 1.278 0 0.0 1e-06 
3.0 1.278 0 0.0 1e-06 
0.05 1.279 0 0.0 1e-06 
3.0 1.279 0 0.0 1e-06 
0.05 1.28 0 0.0 1e-06 
3.0 1.28 0 0.0 1e-06 
0.05 1.281 0 0.0 1e-06 
3.0 1.281 0 0.0 1e-06 
0.05 1.282 0 0.0 1e-06 
3.0 1.282 0 0.0 1e-06 
0.05 1.283 0 0.0 1e-06 
3.0 1.283 0 0.0 1e-06 
0.05 1.284 0 0.0 1e-06 
3.0 1.284 0 0.0 1e-06 
0.05 1.285 0 0.0 1e-06 
3.0 1.285 0 0.0 1e-06 
0.05 1.286 0 0.0 1e-06 
3.0 1.286 0 0.0 1e-06 
0.05 1.287 0 0.0 1e-06 
3.0 1.287 0 0.0 1e-06 
0.05 1.288 0 0.0 1e-06 
3.0 1.288 0 0.0 1e-06 
0.05 1.289 0 0.0 1e-06 
3.0 1.289 0 0.0 1e-06 
0.05 1.29 0 0.0 1e-06 
3.0 1.29 0 0.0 1e-06 
0.05 1.291 0 0.0 1e-06 
3.0 1.291 0 0.0 1e-06 
0.05 1.292 0 0.0 1e-06 
3.0 1.292 0 0.0 1e-06 
0.05 1.293 0 0.0 1e-06 
3.0 1.293 0 0.0 1e-06 
0.05 1.294 0 0.0 1e-06 
3.0 1.294 0 0.0 1e-06 
0.05 1.295 0 0.0 1e-06 
3.0 1.295 0 0.0 1e-06 
0.05 1.296 0 0.0 1e-06 
3.0 1.296 0 0.0 1e-06 
0.05 1.297 0 0.0 1e-06 
3.0 1.297 0 0.0 1e-06 
0.05 1.298 0 0.0 1e-06 
3.0 1.298 0 0.0 1e-06 
0.05 1.299 0 0.0 1e-06 
3.0 1.299 0 0.0 1e-06 
0.05 1.3 0 0.0 1e-06 
3.0 1.3 0 0.0 1e-06 
0.05 1.301 0 0.0 1e-06 
3.0 1.301 0 0.0 1e-06 
0.05 1.302 0 0.0 1e-06 
3.0 1.302 0 0.0 1e-06 
0.05 1.303 0 0.0 1e-06 
3.0 1.303 0 0.0 1e-06 
0.05 1.304 0 0.0 1e-06 
3.0 1.304 0 0.0 1e-06 
0.05 1.305 0 0.0 1e-06 
3.0 1.305 0 0.0 1e-06 
0.05 1.306 0 0.0 1e-06 
3.0 1.306 0 0.0 1e-06 
0.05 1.307 0 0.0 1e-06 
3.0 1.307 0 0.0 1e-06 
0.05 1.308 0 0.0 1e-06 
3.0 1.308 0 0.0 1e-06 
0.05 1.309 0 0.0 1e-06 
3.0 1.309 0 0.0 1e-06 
0.05 1.31 0 0.0 1e-06 
3.0 1.31 0 0.0 1e-06 
0.05 1.311 0 0.0 1e-06 
3.0 1.311 0 0.0 1e-06 
0.05 1.312 0 0.0 1e-06 
3.0 1.312 0 0.0 1e-06 
0.05 1.313 0 0.0 1e-06 
3.0 1.313 0 0.0 1e-06 
0.05 1.314 0 0.0 1e-06 
3.0 1.314 0 0.0 1e-06 
0.05 1.315 0 0.0 1e-06 
3.0 1.315 0 0.0 1e-06 
0.05 1.316 0 0.0 1e-06 
3.0 1.316 0 0.0 1e-06 
0.05 1.317 0 0.0 1e-06 
3.0 1.317 0 0.0 1e-06 
0.05 1.318 0 0.0 1e-06 
3.0 1.318 0 0.0 1e-06 
0.05 1.319 0 0.0 1e-06 
3.0 1.319 0 0.0 1e-06 
0.05 1.32 0 0.0 1e-06 
3.0 1.32 0 0.0 1e-06 
0.05 1.321 0 0.0 1e-06 
3.0 1.321 0 0.0 1e-06 
0.05 1.322 0 0.0 1e-06 
3.0 1.322 0 0.0 1e-06 
0.05 1.323 0 0.0 1e-06 
3.0 1.323 0 0.0 1e-06 
0.05 1.324 0 0.0 1e-06 
3.0 1.324 0 0.0 1e-06 
0.05 1.325 0 0.0 1e-06 
3.0 1.325 0 0.0 1e-06 
0.05 1.326 0 0.0 1e-06 
3.0 1.326 0 0.0 1e-06 
0.05 1.327 0 0.0 1e-06 
3.0 1.327 0 0.0 1e-06 
0.05 1.328 0 0.0 1e-06 
3.0 1.328 0 0.0 1e-06 
0.05 1.329 0 0.0 1e-06 
3.0 1.329 0 0.0 1e-06 
0.05 1.33 0 0.0 1e-06 
3.0 1.33 0 0.0 1e-06 
0.05 1.331 0 0.0 1e-06 
3.0 1.331 0 0.0 1e-06 
0.05 1.332 0 0.0 1e-06 
3.0 1.332 0 0.0 1e-06 
0.05 1.333 0 0.0 1e-06 
3.0 1.333 0 0.0 1e-06 
0.05 1.334 0 0.0 1e-06 
3.0 1.334 0 0.0 1e-06 
0.05 1.335 0 0.0 1e-06 
3.0 1.335 0 0.0 1e-06 
0.05 1.336 0 0.0 1e-06 
3.0 1.336 0 0.0 1e-06 
0.05 1.337 0 0.0 1e-06 
3.0 1.337 0 0.0 1e-06 
0.05 1.338 0 0.0 1e-06 
3.0 1.338 0 0.0 1e-06 
0.05 1.339 0 0.0 1e-06 
3.0 1.339 0 0.0 1e-06 
0.05 1.34 0 0.0 1e-06 
3.0 1.34 0 0.0 1e-06 
0.05 1.341 0 0.0 1e-06 
3.0 1.341 0 0.0 1e-06 
0.05 1.342 0 0.0 1e-06 
3.0 1.342 0 0.0 1e-06 
0.05 1.343 0 0.0 1e-06 
3.0 1.343 0 0.0 1e-06 
0.05 1.344 0 0.0 1e-06 
3.0 1.344 0 0.0 1e-06 
0.05 1.345 0 0.0 1e-06 
3.0 1.345 0 0.0 1e-06 
0.05 1.346 0 0.0 1e-06 
3.0 1.346 0 0.0 1e-06 
0.05 1.347 0 0.0 1e-06 
3.0 1.347 0 0.0 1e-06 
0.05 1.348 0 0.0 1e-06 
3.0 1.348 0 0.0 1e-06 
0.05 1.349 0 0.0 1e-06 
3.0 1.349 0 0.0 1e-06 
0.05 1.35 0 0.0 1e-06 
3.0 1.35 0 0.0 1e-06 
0.05 1.351 0 0.0 1e-06 
3.0 1.351 0 0.0 1e-06 
0.05 1.352 0 0.0 1e-06 
3.0 1.352 0 0.0 1e-06 
0.05 1.353 0 0.0 1e-06 
3.0 1.353 0 0.0 1e-06 
0.05 1.354 0 0.0 1e-06 
3.0 1.354 0 0.0 1e-06 
0.05 1.355 0 0.0 1e-06 
3.0 1.355 0 0.0 1e-06 
0.05 1.356 0 0.0 1e-06 
3.0 1.356 0 0.0 1e-06 
0.05 1.357 0 0.0 1e-06 
3.0 1.357 0 0.0 1e-06 
0.05 1.358 0 0.0 1e-06 
3.0 1.358 0 0.0 1e-06 
0.05 1.359 0 0.0 1e-06 
3.0 1.359 0 0.0 1e-06 
0.05 1.36 0 0.0 1e-06 
3.0 1.36 0 0.0 1e-06 
0.05 1.361 0 0.0 1e-06 
3.0 1.361 0 0.0 1e-06 
0.05 1.362 0 0.0 1e-06 
3.0 1.362 0 0.0 1e-06 
0.05 1.363 0 0.0 1e-06 
3.0 1.363 0 0.0 1e-06 
0.05 1.364 0 0.0 1e-06 
3.0 1.364 0 0.0 1e-06 
0.05 1.365 0 0.0 1e-06 
3.0 1.365 0 0.0 1e-06 
0.05 1.366 0 0.0 1e-06 
3.0 1.366 0 0.0 1e-06 
0.05 1.367 0 0.0 1e-06 
3.0 1.367 0 0.0 1e-06 
0.05 1.368 0 0.0 1e-06 
3.0 1.368 0 0.0 1e-06 
0.05 1.369 0 0.0 1e-06 
3.0 1.369 0 0.0 1e-06 
0.05 1.37 0 0.0 1e-06 
3.0 1.37 0 0.0 1e-06 
0.05 1.371 0 0.0 1e-06 
3.0 1.371 0 0.0 1e-06 
0.05 1.372 0 0.0 1e-06 
3.0 1.372 0 0.0 1e-06 
0.05 1.373 0 0.0 1e-06 
3.0 1.373 0 0.0 1e-06 
0.05 1.374 0 0.0 1e-06 
3.0 1.374 0 0.0 1e-06 
0.05 1.375 0 0.0 1e-06 
3.0 1.375 0 0.0 1e-06 
0.05 1.376 0 0.0 1e-06 
3.0 1.376 0 0.0 1e-06 
0.05 1.377 0 0.0 1e-06 
3.0 1.377 0 0.0 1e-06 
0.05 1.378 0 0.0 1e-06 
3.0 1.378 0 0.0 1e-06 
0.05 1.379 0 0.0 1e-06 
3.0 1.379 0 0.0 1e-06 
0.05 1.38 0 0.0 1e-06 
3.0 1.38 0 0.0 1e-06 
0.05 1.381 0 0.0 1e-06 
3.0 1.381 0 0.0 1e-06 
0.05 1.382 0 0.0 1e-06 
3.0 1.382 0 0.0 1e-06 
0.05 1.383 0 0.0 1e-06 
3.0 1.383 0 0.0 1e-06 
0.05 1.384 0 0.0 1e-06 
3.0 1.384 0 0.0 1e-06 
0.05 1.385 0 0.0 1e-06 
3.0 1.385 0 0.0 1e-06 
0.05 1.386 0 0.0 1e-06 
3.0 1.386 0 0.0 1e-06 
0.05 1.387 0 0.0 1e-06 
3.0 1.387 0 0.0 1e-06 
0.05 1.388 0 0.0 1e-06 
3.0 1.388 0 0.0 1e-06 
0.05 1.389 0 0.0 1e-06 
3.0 1.389 0 0.0 1e-06 
0.05 1.39 0 0.0 1e-06 
3.0 1.39 0 0.0 1e-06 
0.05 1.391 0 0.0 1e-06 
3.0 1.391 0 0.0 1e-06 
0.05 1.392 0 0.0 1e-06 
3.0 1.392 0 0.0 1e-06 
0.05 1.393 0 0.0 1e-06 
3.0 1.393 0 0.0 1e-06 
0.05 1.394 0 0.0 1e-06 
3.0 1.394 0 0.0 1e-06 
0.05 1.395 0 0.0 1e-06 
3.0 1.395 0 0.0 1e-06 
0.05 1.396 0 0.0 1e-06 
3.0 1.396 0 0.0 1e-06 
0.05 1.397 0 0.0 1e-06 
3.0 1.397 0 0.0 1e-06 
0.05 1.398 0 0.0 1e-06 
3.0 1.398 0 0.0 1e-06 
0.05 1.399 0 0.0 1e-06 
3.0 1.399 0 0.0 1e-06 
0.05 1.4 0 0.0 1e-06 
3.0 1.4 0 0.0 1e-06 
0.05 1.401 0 0.0 1e-06 
3.0 1.401 0 0.0 1e-06 
0.05 1.402 0 0.0 1e-06 
3.0 1.402 0 0.0 1e-06 
0.05 1.403 0 0.0 1e-06 
3.0 1.403 0 0.0 1e-06 
0.05 1.404 0 0.0 1e-06 
3.0 1.404 0 0.0 1e-06 
0.05 1.405 0 0.0 1e-06 
3.0 1.405 0 0.0 1e-06 
0.05 1.406 0 0.0 1e-06 
3.0 1.406 0 0.0 1e-06 
0.05 1.407 0 0.0 1e-06 
3.0 1.407 0 0.0 1e-06 
0.05 1.408 0 0.0 1e-06 
3.0 1.408 0 0.0 1e-06 
0.05 1.409 0 0.0 1e-06 
3.0 1.409 0 0.0 1e-06 
0.05 1.41 0 0.0 1e-06 
3.0 1.41 0 0.0 1e-06 
0.05 1.411 0 0.0 1e-06 
3.0 1.411 0 0.0 1e-06 
0.05 1.412 0 0.0 1e-06 
3.0 1.412 0 0.0 1e-06 
0.05 1.413 0 0.0 1e-06 
3.0 1.413 0 0.0 1e-06 
0.05 1.414 0 0.0 1e-06 
3.0 1.414 0 0.0 1e-06 
0.05 1.415 0 0.0 1e-06 
3.0 1.415 0 0.0 1e-06 
0.05 1.416 0 0.0 1e-06 
3.0 1.416 0 0.0 1e-06 
0.05 1.417 0 0.0 1e-06 
3.0 1.417 0 0.0 1e-06 
0.05 1.418 0 0.0 1e-06 
3.0 1.418 0 0.0 1e-06 
0.05 1.419 0 0.0 1e-06 
3.0 1.419 0 0.0 1e-06 
0.05 1.42 0 0.0 1e-06 
3.0 1.42 0 0.0 1e-06 
0.05 1.421 0 0.0 1e-06 
3.0 1.421 0 0.0 1e-06 
0.05 1.422 0 0.0 1e-06 
3.0 1.422 0 0.0 1e-06 
0.05 1.423 0 0.0 1e-06 
3.0 1.423 0 0.0 1e-06 
0.05 1.424 0 0.0 1e-06 
3.0 1.424 0 0.0 1e-06 
0.05 1.425 0 0.0 1e-06 
3.0 1.425 0 0.0 1e-06 
0.05 1.426 0 0.0 1e-06 
3.0 1.426 0 0.0 1e-06 
0.05 1.427 0 0.0 1e-06 
3.0 1.427 0 0.0 1e-06 
0.05 1.428 0 0.0 1e-06 
3.0 1.428 0 0.0 1e-06 
0.05 1.429 0 0.0 1e-06 
3.0 1.429 0 0.0 1e-06 
0.05 1.43 0 0.0 1e-06 
3.0 1.43 0 0.0 1e-06 
0.05 1.431 0 0.0 1e-06 
3.0 1.431 0 0.0 1e-06 
0.05 1.432 0 0.0 1e-06 
3.0 1.432 0 0.0 1e-06 
0.05 1.433 0 0.0 1e-06 
3.0 1.433 0 0.0 1e-06 
0.05 1.434 0 0.0 1e-06 
3.0 1.434 0 0.0 1e-06 
0.05 1.435 0 0.0 1e-06 
3.0 1.435 0 0.0 1e-06 
0.05 1.436 0 0.0 1e-06 
3.0 1.436 0 0.0 1e-06 
0.05 1.437 0 0.0 1e-06 
3.0 1.437 0 0.0 1e-06 
0.05 1.438 0 0.0 1e-06 
3.0 1.438 0 0.0 1e-06 
0.05 1.439 0 0.0 1e-06 
3.0 1.439 0 0.0 1e-06 
0.05 1.44 0 0.0 1e-06 
3.0 1.44 0 0.0 1e-06 
0.05 1.441 0 0.0 1e-06 
3.0 1.441 0 0.0 1e-06 
0.05 1.442 0 0.0 1e-06 
3.0 1.442 0 0.0 1e-06 
0.05 1.443 0 0.0 1e-06 
3.0 1.443 0 0.0 1e-06 
0.05 1.444 0 0.0 1e-06 
3.0 1.444 0 0.0 1e-06 
0.05 1.445 0 0.0 1e-06 
3.0 1.445 0 0.0 1e-06 
0.05 1.446 0 0.0 1e-06 
3.0 1.446 0 0.0 1e-06 
0.05 1.447 0 0.0 1e-06 
3.0 1.447 0 0.0 1e-06 
0.05 1.448 0 0.0 1e-06 
3.0 1.448 0 0.0 1e-06 
0.05 1.449 0 0.0 1e-06 
3.0 1.449 0 0.0 1e-06 
0.05 1.45 0 0.0 1e-06 
3.0 1.45 0 0.0 1e-06 
0.05 1.451 0 0.0 1e-06 
3.0 1.451 0 0.0 1e-06 
0.05 1.452 0 0.0 1e-06 
3.0 1.452 0 0.0 1e-06 
0.05 1.453 0 0.0 1e-06 
3.0 1.453 0 0.0 1e-06 
0.05 1.454 0 0.0 1e-06 
3.0 1.454 0 0.0 1e-06 
0.05 1.455 0 0.0 1e-06 
3.0 1.455 0 0.0 1e-06 
0.05 1.456 0 0.0 1e-06 
3.0 1.456 0 0.0 1e-06 
0.05 1.457 0 0.0 1e-06 
3.0 1.457 0 0.0 1e-06 
0.05 1.458 0 0.0 1e-06 
3.0 1.458 0 0.0 1e-06 
0.05 1.459 0 0.0 1e-06 
3.0 1.459 0 0.0 1e-06 
0.05 1.46 0 0.0 1e-06 
3.0 1.46 0 0.0 1e-06 
0.05 1.461 0 0.0 1e-06 
3.0 1.461 0 0.0 1e-06 
0.05 1.462 0 0.0 1e-06 
3.0 1.462 0 0.0 1e-06 
0.05 1.463 0 0.0 1e-06 
3.0 1.463 0 0.0 1e-06 
0.05 1.464 0 0.0 1e-06 
3.0 1.464 0 0.0 1e-06 
0.05 1.465 0 0.0 1e-06 
3.0 1.465 0 0.0 1e-06 
0.05 1.466 0 0.0 1e-06 
3.0 1.466 0 0.0 1e-06 
0.05 1.467 0 0.0 1e-06 
3.0 1.467 0 0.0 1e-06 
0.05 1.468 0 0.0 1e-06 
3.0 1.468 0 0.0 1e-06 
0.05 1.469 0 0.0 1e-06 
3.0 1.469 0 0.0 1e-06 
0.05 1.47 0 0.0 1e-06 
3.0 1.47 0 0.0 1e-06 
0.05 1.471 0 0.0 1e-06 
3.0 1.471 0 0.0 1e-06 
0.05 1.472 0 0.0 1e-06 
3.0 1.472 0 0.0 1e-06 
0.05 1.473 0 0.0 1e-06 
3.0 1.473 0 0.0 1e-06 
0.05 1.474 0 0.0 1e-06 
3.0 1.474 0 0.0 1e-06 
0.05 1.475 0 0.0 1e-06 
3.0 1.475 0 0.0 1e-06 
0.05 1.476 0 0.0 1e-06 
3.0 1.476 0 0.0 1e-06 
0.05 1.477 0 0.0 1e-06 
3.0 1.477 0 0.0 1e-06 
0.05 1.478 0 0.0 1e-06 
3.0 1.478 0 0.0 1e-06 
0.05 1.479 0 0.0 1e-06 
3.0 1.479 0 0.0 1e-06 
0.05 1.48 0 0.0 1e-06 
3.0 1.48 0 0.0 1e-06 
0.05 1.481 0 0.0 1e-06 
3.0 1.481 0 0.0 1e-06 
0.05 1.482 0 0.0 1e-06 
3.0 1.482 0 0.0 1e-06 
0.05 1.483 0 0.0 1e-06 
3.0 1.483 0 0.0 1e-06 
0.05 1.484 0 0.0 1e-06 
3.0 1.484 0 0.0 1e-06 
0.05 1.485 0 0.0 1e-06 
3.0 1.485 0 0.0 1e-06 
0.05 1.486 0 0.0 1e-06 
3.0 1.486 0 0.0 1e-06 
0.05 1.487 0 0.0 1e-06 
3.0 1.487 0 0.0 1e-06 
0.05 1.488 0 0.0 1e-06 
3.0 1.488 0 0.0 1e-06 
0.05 1.489 0 0.0 1e-06 
3.0 1.489 0 0.0 1e-06 
0.05 1.49 0 0.0 1e-06 
3.0 1.49 0 0.0 1e-06 
0.05 1.491 0 0.0 1e-06 
3.0 1.491 0 0.0 1e-06 
0.05 1.492 0 0.0 1e-06 
3.0 1.492 0 0.0 1e-06 
0.05 1.493 0 0.0 1e-06 
3.0 1.493 0 0.0 1e-06 
0.05 1.494 0 0.0 1e-06 
3.0 1.494 0 0.0 1e-06 
0.05 1.495 0 0.0 1e-06 
3.0 1.495 0 0.0 1e-06 
0.05 1.496 0 0.0 1e-06 
3.0 1.496 0 0.0 1e-06 
0.05 1.497 0 0.0 1e-06 
3.0 1.497 0 0.0 1e-06 
0.05 1.498 0 0.0 1e-06 
3.0 1.498 0 0.0 1e-06 
0.05 1.499 0 0.0 1e-06 
3.0 1.499 0 0.0 1e-06 
0.05 1.5 0 0.0 1e-06 
3.0 1.5 0 0.0 1e-06 
0.05 1.501 0 0.0 1e-06 
3.0 1.501 0 0.0 1e-06 
0.05 1.502 0 0.0 1e-06 
3.0 1.502 0 0.0 1e-06 
0.05 1.503 0 0.0 1e-06 
3.0 1.503 0 0.0 1e-06 
0.05 1.504 0 0.0 1e-06 
3.0 1.504 0 0.0 1e-06 
0.05 1.505 0 0.0 1e-06 
3.0 1.505 0 0.0 1e-06 
0.05 1.506 0 0.0 1e-06 
3.0 1.506 0 0.0 1e-06 
0.05 1.507 0 0.0 1e-06 
3.0 1.507 0 0.0 1e-06 
0.05 1.508 0 0.0 1e-06 
3.0 1.508 0 0.0 1e-06 
0.05 1.509 0 0.0 1e-06 
3.0 1.509 0 0.0 1e-06 
0.05 1.51 0 0.0 1e-06 
3.0 1.51 0 0.0 1e-06 
0.05 1.511 0 0.0 1e-06 
3.0 1.511 0 0.0 1e-06 
0.05 1.512 0 0.0 1e-06 
3.0 1.512 0 0.0 1e-06 
0.05 1.513 0 0.0 1e-06 
3.0 1.513 0 0.0 1e-06 
0.05 1.514 0 0.0 1e-06 
3.0 1.514 0 0.0 1e-06 
0.05 1.515 0 0.0 1e-06 
3.0 1.515 0 0.0 1e-06 
0.05 1.516 0 0.0 1e-06 
3.0 1.516 0 0.0 1e-06 
0.05 1.517 0 0.0 1e-06 
3.0 1.517 0 0.0 1e-06 
0.05 1.518 0 0.0 1e-06 
3.0 1.518 0 0.0 1e-06 
0.05 1.519 0 0.0 1e-06 
3.0 1.519 0 0.0 1e-06 
0.05 1.52 0 0.0 1e-06 
3.0 1.52 0 0.0 1e-06 
0.05 1.521 0 0.0 1e-06 
3.0 1.521 0 0.0 1e-06 
0.05 1.522 0 0.0 1e-06 
3.0 1.522 0 0.0 1e-06 
0.05 1.523 0 0.0 1e-06 
3.0 1.523 0 0.0 1e-06 
0.05 1.524 0 0.0 1e-06 
3.0 1.524 0 0.0 1e-06 
0.05 1.525 0 0.0 1e-06 
3.0 1.525 0 0.0 1e-06 
0.05 1.526 0 0.0 1e-06 
3.0 1.526 0 0.0 1e-06 
0.05 1.527 0 0.0 1e-06 
3.0 1.527 0 0.0 1e-06 
0.05 1.528 0 0.0 1e-06 
3.0 1.528 0 0.0 1e-06 
0.05 1.529 0 0.0 1e-06 
3.0 1.529 0 0.0 1e-06 
0.05 1.53 0 0.0 1e-06 
3.0 1.53 0 0.0 1e-06 
0.05 1.531 0 0.0 1e-06 
3.0 1.531 0 0.0 1e-06 
0.05 1.532 0 0.0 1e-06 
3.0 1.532 0 0.0 1e-06 
0.05 1.533 0 0.0 1e-06 
3.0 1.533 0 0.0 1e-06 
0.05 1.534 0 0.0 1e-06 
3.0 1.534 0 0.0 1e-06 
0.05 1.535 0 0.0 1e-06 
3.0 1.535 0 0.0 1e-06 
0.05 1.536 0 0.0 1e-06 
3.0 1.536 0 0.0 1e-06 
0.05 1.537 0 0.0 1e-06 
3.0 1.537 0 0.0 1e-06 
0.05 1.538 0 0.0 1e-06 
3.0 1.538 0 0.0 1e-06 
0.05 1.539 0 0.0 1e-06 
3.0 1.539 0 0.0 1e-06 
0.05 1.54 0 0.0 1e-06 
3.0 1.54 0 0.0 1e-06 
0.05 1.541 0 0.0 1e-06 
3.0 1.541 0 0.0 1e-06 
0.05 1.542 0 0.0 1e-06 
3.0 1.542 0 0.0 1e-06 
0.05 1.543 0 0.0 1e-06 
3.0 1.543 0 0.0 1e-06 
0.05 1.544 0 0.0 1e-06 
3.0 1.544 0 0.0 1e-06 
0.05 1.545 0 0.0 1e-06 
3.0 1.545 0 0.0 1e-06 
0.05 1.546 0 0.0 1e-06 
3.0 1.546 0 0.0 1e-06 
0.05 1.547 0 0.0 1e-06 
3.0 1.547 0 0.0 1e-06 
0.05 1.548 0 0.0 1e-06 
3.0 1.548 0 0.0 1e-06 
0.05 1.549 0 0.0 1e-06 
3.0 1.549 0 0.0 1e-06 
0.05 1.55 0 0.0 1e-06 
3.0 1.55 0 0.0 1e-06 
0.05 1.551 0 0.0 1e-06 
3.0 1.551 0 0.0 1e-06 
0.05 1.552 0 0.0 1e-06 
3.0 1.552 0 0.0 1e-06 
0.05 1.553 0 0.0 1e-06 
3.0 1.553 0 0.0 1e-06 
0.05 1.554 0 0.0 1e-06 
3.0 1.554 0 0.0 1e-06 
0.05 1.555 0 0.0 1e-06 
3.0 1.555 0 0.0 1e-06 
0.05 1.556 0 0.0 1e-06 
3.0 1.556 0 0.0 1e-06 
0.05 1.557 0 0.0 1e-06 
3.0 1.557 0 0.0 1e-06 
0.05 1.558 0 0.0 1e-06 
3.0 1.558 0 0.0 1e-06 
0.05 1.559 0 0.0 1e-06 
3.0 1.559 0 0.0 1e-06 
0.05 1.56 0 0.0 1e-06 
3.0 1.56 0 0.0 1e-06 
0.05 1.561 0 0.0 1e-06 
3.0 1.561 0 0.0 1e-06 
0.05 1.562 0 0.0 1e-06 
3.0 1.562 0 0.0 1e-06 
0.05 1.563 0 0.0 1e-06 
3.0 1.563 0 0.0 1e-06 
0.05 1.564 0 0.0 1e-06 
3.0 1.564 0 0.0 1e-06 
0.05 1.565 0 0.0 1e-06 
3.0 1.565 0 0.0 1e-06 
0.05 1.566 0 0.0 1e-06 
3.0 1.566 0 0.0 1e-06 
0.05 1.567 0 0.0 1e-06 
3.0 1.567 0 0.0 1e-06 
0.05 1.568 0 0.0 1e-06 
3.0 1.568 0 0.0 1e-06 
0.05 1.569 0 0.0 1e-06 
3.0 1.569 0 0.0 1e-06 
0.05 1.57 0 0.0 1e-06 
3.0 1.57 0 0.0 1e-06 
0.05 1.571 0 0.0 1e-06 
3.0 1.571 0 0.0 1e-06 
0.05 1.572 0 0.0 1e-06 
3.0 1.572 0 0.0 1e-06 
0.05 1.573 0 0.0 1e-06 
3.0 1.573 0 0.0 1e-06 
0.05 1.574 0 0.0 1e-06 
3.0 1.574 0 0.0 1e-06 
0.05 1.575 0 0.0 1e-06 
3.0 1.575 0 0.0 1e-06 
0.05 1.576 0 0.0 1e-06 
3.0 1.576 0 0.0 1e-06 
0.05 1.577 0 0.0 1e-06 
3.0 1.577 0 0.0 1e-06 
0.05 1.578 0 0.0 1e-06 
3.0 1.578 0 0.0 1e-06 
0.05 1.579 0 0.0 1e-06 
3.0 1.579 0 0.0 1e-06 
0.05 1.58 0 0.0 1e-06 
3.0 1.58 0 0.0 1e-06 
0.05 1.581 0 0.0 1e-06 
3.0 1.581 0 0.0 1e-06 
0.05 1.582 0 0.0 1e-06 
3.0 1.582 0 0.0 1e-06 
0.05 1.583 0 0.0 1e-06 
3.0 1.583 0 0.0 1e-06 
0.05 1.584 0 0.0 1e-06 
3.0 1.584 0 0.0 1e-06 
0.05 1.585 0 0.0 1e-06 
3.0 1.585 0 0.0 1e-06 
0.05 1.586 0 0.0 1e-06 
3.0 1.586 0 0.0 1e-06 
0.05 1.587 0 0.0 1e-06 
3.0 1.587 0 0.0 1e-06 
0.05 1.588 0 0.0 1e-06 
3.0 1.588 0 0.0 1e-06 
0.05 1.589 0 0.0 1e-06 
3.0 1.589 0 0.0 1e-06 
0.05 1.59 0 0.0 1e-06 
3.0 1.59 0 0.0 1e-06 
0.05 1.591 0 0.0 1e-06 
3.0 1.591 0 0.0 1e-06 
0.05 1.592 0 0.0 1e-06 
3.0 1.592 0 0.0 1e-06 
0.05 1.593 0 0.0 1e-06 
3.0 1.593 0 0.0 1e-06 
0.05 1.594 0 0.0 1e-06 
3.0 1.594 0 0.0 1e-06 
0.05 1.595 0 0.0 1e-06 
3.0 1.595 0 0.0 1e-06 
0.05 1.596 0 0.0 1e-06 
3.0 1.596 0 0.0 1e-06 
0.05 1.597 0 0.0 1e-06 
3.0 1.597 0 0.0 1e-06 
0.05 1.598 0 0.0 1e-06 
3.0 1.598 0 0.0 1e-06 
0.05 1.599 0 0.0 1e-06 
3.0 1.599 0 0.0 1e-06 
0.05 1.6 0 0.0 1e-06 
3.0 1.6 0 0.0 1e-06 
0.05 1.601 0 0.0 1e-06 
3.0 1.601 0 0.0 1e-06 
0.05 1.602 0 0.0 1e-06 
3.0 1.602 0 0.0 1e-06 
0.05 1.603 0 0.0 1e-06 
3.0 1.603 0 0.0 1e-06 
0.05 1.604 0 0.0 1e-06 
3.0 1.604 0 0.0 1e-06 
0.05 1.605 0 0.0 1e-06 
3.0 1.605 0 0.0 1e-06 
0.05 1.606 0 0.0 1e-06 
3.0 1.606 0 0.0 1e-06 
0.05 1.607 0 0.0 1e-06 
3.0 1.607 0 0.0 1e-06 
0.05 1.608 0 0.0 1e-06 
3.0 1.608 0 0.0 1e-06 
0.05 1.609 0 0.0 1e-06 
3.0 1.609 0 0.0 1e-06 
0.05 1.61 0 0.0 1e-06 
3.0 1.61 0 0.0 1e-06 
0.05 1.611 0 0.0 1e-06 
3.0 1.611 0 0.0 1e-06 
0.05 1.612 0 0.0 1e-06 
3.0 1.612 0 0.0 1e-06 
0.05 1.613 0 0.0 1e-06 
3.0 1.613 0 0.0 1e-06 
0.05 1.614 0 0.0 1e-06 
3.0 1.614 0 0.0 1e-06 
0.05 1.615 0 0.0 1e-06 
3.0 1.615 0 0.0 1e-06 
0.05 1.616 0 0.0 1e-06 
3.0 1.616 0 0.0 1e-06 
0.05 1.617 0 0.0 1e-06 
3.0 1.617 0 0.0 1e-06 
0.05 1.618 0 0.0 1e-06 
3.0 1.618 0 0.0 1e-06 
0.05 1.619 0 0.0 1e-06 
3.0 1.619 0 0.0 1e-06 
0.05 1.62 0 0.0 1e-06 
3.0 1.62 0 0.0 1e-06 
0.05 1.621 0 0.0 1e-06 
3.0 1.621 0 0.0 1e-06 
0.05 1.622 0 0.0 1e-06 
3.0 1.622 0 0.0 1e-06 
0.05 1.623 0 0.0 1e-06 
3.0 1.623 0 0.0 1e-06 
0.05 1.624 0 0.0 1e-06 
3.0 1.624 0 0.0 1e-06 
0.05 1.625 0 0.0 1e-06 
3.0 1.625 0 0.0 1e-06 
0.05 1.626 0 0.0 1e-06 
3.0 1.626 0 0.0 1e-06 
0.05 1.627 0 0.0 1e-06 
3.0 1.627 0 0.0 1e-06 
0.05 1.628 0 0.0 1e-06 
3.0 1.628 0 0.0 1e-06 
0.05 1.629 0 0.0 1e-06 
3.0 1.629 0 0.0 1e-06 
0.05 1.63 0 0.0 1e-06 
3.0 1.63 0 0.0 1e-06 
0.05 1.631 0 0.0 1e-06 
3.0 1.631 0 0.0 1e-06 
0.05 1.632 0 0.0 1e-06 
3.0 1.632 0 0.0 1e-06 
0.05 1.633 0 0.0 1e-06 
3.0 1.633 0 0.0 1e-06 
0.05 1.634 0 0.0 1e-06 
3.0 1.634 0 0.0 1e-06 
0.05 1.635 0 0.0 1e-06 
3.0 1.635 0 0.0 1e-06 
0.05 1.636 0 0.0 1e-06 
3.0 1.636 0 0.0 1e-06 
0.05 1.637 0 0.0 1e-06 
3.0 1.637 0 0.0 1e-06 
0.05 1.638 0 0.0 1e-06 
3.0 1.638 0 0.0 1e-06 
0.05 1.639 0 0.0 1e-06 
3.0 1.639 0 0.0 1e-06 
0.05 1.64 0 0.0 1e-06 
3.0 1.64 0 0.0 1e-06 
0.05 1.641 0 0.0 1e-06 
3.0 1.641 0 0.0 1e-06 
0.05 1.642 0 0.0 1e-06 
3.0 1.642 0 0.0 1e-06 
0.05 1.643 0 0.0 1e-06 
3.0 1.643 0 0.0 1e-06 
0.05 1.644 0 0.0 1e-06 
3.0 1.644 0 0.0 1e-06 
0.05 1.645 0 0.0 1e-06 
3.0 1.645 0 0.0 1e-06 
0.05 1.646 0 0.0 1e-06 
3.0 1.646 0 0.0 1e-06 
0.05 1.647 0 0.0 1e-06 
3.0 1.647 0 0.0 1e-06 
0.05 1.648 0 0.0 1e-06 
3.0 1.648 0 0.0 1e-06 
0.05 1.649 0 0.0 1e-06 
3.0 1.649 0 0.0 1e-06 
0.05 1.65 0 0.0 1e-06 
3.0 1.65 0 0.0 1e-06 
0.05 1.651 0 0.0 1e-06 
3.0 1.651 0 0.0 1e-06 
0.05 1.652 0 0.0 1e-06 
3.0 1.652 0 0.0 1e-06 
0.05 1.653 0 0.0 1e-06 
3.0 1.653 0 0.0 1e-06 
0.05 1.654 0 0.0 1e-06 
3.0 1.654 0 0.0 1e-06 
0.05 1.655 0 0.0 1e-06 
3.0 1.655 0 0.0 1e-06 
0.05 1.656 0 0.0 1e-06 
3.0 1.656 0 0.0 1e-06 
0.05 1.657 0 0.0 1e-06 
3.0 1.657 0 0.0 1e-06 
0.05 1.658 0 0.0 1e-06 
3.0 1.658 0 0.0 1e-06 
0.05 1.659 0 0.0 1e-06 
3.0 1.659 0 0.0 1e-06 
0.05 1.66 0 0.0 1e-06 
3.0 1.66 0 0.0 1e-06 
0.05 1.661 0 0.0 1e-06 
3.0 1.661 0 0.0 1e-06 
0.05 1.662 0 0.0 1e-06 
3.0 1.662 0 0.0 1e-06 
0.05 1.663 0 0.0 1e-06 
3.0 1.663 0 0.0 1e-06 
0.05 1.664 0 0.0 1e-06 
3.0 1.664 0 0.0 1e-06 
0.05 1.665 0 0.0 1e-06 
3.0 1.665 0 0.0 1e-06 
0.05 1.666 0 0.0 1e-06 
3.0 1.666 0 0.0 1e-06 
0.05 1.667 0 0.0 1e-06 
3.0 1.667 0 0.0 1e-06 
0.05 1.668 0 0.0 1e-06 
3.0 1.668 0 0.0 1e-06 
0.05 1.669 0 0.0 1e-06 
3.0 1.669 0 0.0 1e-06 
0.05 1.67 0 0.0 1e-06 
3.0 1.67 0 0.0 1e-06 
0.05 1.671 0 0.0 1e-06 
3.0 1.671 0 0.0 1e-06 
0.05 1.672 0 0.0 1e-06 
3.0 1.672 0 0.0 1e-06 
0.05 1.673 0 0.0 1e-06 
3.0 1.673 0 0.0 1e-06 
0.05 1.674 0 0.0 1e-06 
3.0 1.674 0 0.0 1e-06 
0.05 1.675 0 0.0 1e-06 
3.0 1.675 0 0.0 1e-06 
0.05 1.676 0 0.0 1e-06 
3.0 1.676 0 0.0 1e-06 
0.05 1.677 0 0.0 1e-06 
3.0 1.677 0 0.0 1e-06 
0.05 1.678 0 0.0 1e-06 
3.0 1.678 0 0.0 1e-06 
0.05 1.679 0 0.0 1e-06 
3.0 1.679 0 0.0 1e-06 
0.05 1.68 0 0.0 1e-06 
3.0 1.68 0 0.0 1e-06 
0.05 1.681 0 0.0 1e-06 
3.0 1.681 0 0.0 1e-06 
0.05 1.682 0 0.0 1e-06 
3.0 1.682 0 0.0 1e-06 
0.05 1.683 0 0.0 1e-06 
3.0 1.683 0 0.0 1e-06 
0.05 1.684 0 0.0 1e-06 
3.0 1.684 0 0.0 1e-06 
0.05 1.685 0 0.0 1e-06 
3.0 1.685 0 0.0 1e-06 
0.05 1.686 0 0.0 1e-06 
3.0 1.686 0 0.0 1e-06 
0.05 1.687 0 0.0 1e-06 
3.0 1.687 0 0.0 1e-06 
0.05 1.688 0 0.0 1e-06 
3.0 1.688 0 0.0 1e-06 
0.05 1.689 0 0.0 1e-06 
3.0 1.689 0 0.0 1e-06 
0.05 1.69 0 0.0 1e-06 
3.0 1.69 0 0.0 1e-06 
0.05 1.691 0 0.0 1e-06 
3.0 1.691 0 0.0 1e-06 
0.05 1.692 0 0.0 1e-06 
3.0 1.692 0 0.0 1e-06 
0.05 1.693 0 0.0 1e-06 
3.0 1.693 0 0.0 1e-06 
0.05 1.694 0 0.0 1e-06 
3.0 1.694 0 0.0 1e-06 
0.05 1.695 0 0.0 1e-06 
3.0 1.695 0 0.0 1e-06 
0.05 1.696 0 0.0 1e-06 
3.0 1.696 0 0.0 1e-06 
0.05 1.697 0 0.0 1e-06 
3.0 1.697 0 0.0 1e-06 
0.05 1.698 0 0.0 1e-06 
3.0 1.698 0 0.0 1e-06 
0.05 1.699 0 0.0 1e-06 
3.0 1.699 0 0.0 1e-06 
0.05 1.7 0 0.0 1e-06 
3.0 1.7 0 0.0 1e-06 
0.05 1.701 0 0.0 1e-06 
3.0 1.701 0 0.0 1e-06 
0.05 1.702 0 0.0 1e-06 
3.0 1.702 0 0.0 1e-06 
0.05 1.703 0 0.0 1e-06 
3.0 1.703 0 0.0 1e-06 
0.05 1.704 0 0.0 1e-06 
3.0 1.704 0 0.0 1e-06 
0.05 1.705 0 0.0 1e-06 
3.0 1.705 0 0.0 1e-06 
0.05 1.706 0 0.0 1e-06 
3.0 1.706 0 0.0 1e-06 
0.05 1.707 0 0.0 1e-06 
3.0 1.707 0 0.0 1e-06 
0.05 1.708 0 0.0 1e-06 
3.0 1.708 0 0.0 1e-06 
0.05 1.709 0 0.0 1e-06 
3.0 1.709 0 0.0 1e-06 
0.05 1.71 0 0.0 1e-06 
3.0 1.71 0 0.0 1e-06 
0.05 1.711 0 0.0 1e-06 
3.0 1.711 0 0.0 1e-06 
0.05 1.712 0 0.0 1e-06 
3.0 1.712 0 0.0 1e-06 
0.05 1.713 0 0.0 1e-06 
3.0 1.713 0 0.0 1e-06 
0.05 1.714 0 0.0 1e-06 
3.0 1.714 0 0.0 1e-06 
0.05 1.715 0 0.0 1e-06 
3.0 1.715 0 0.0 1e-06 
0.05 1.716 0 0.0 1e-06 
3.0 1.716 0 0.0 1e-06 
0.05 1.717 0 0.0 1e-06 
3.0 1.717 0 0.0 1e-06 
0.05 1.718 0 0.0 1e-06 
3.0 1.718 0 0.0 1e-06 
0.05 1.719 0 0.0 1e-06 
3.0 1.719 0 0.0 1e-06 
0.05 1.72 0 0.0 1e-06 
3.0 1.72 0 0.0 1e-06 
0.05 1.721 0 0.0 1e-06 
3.0 1.721 0 0.0 1e-06 
0.05 1.722 0 0.0 1e-06 
3.0 1.722 0 0.0 1e-06 
0.05 1.723 0 0.0 1e-06 
3.0 1.723 0 0.0 1e-06 
0.05 1.724 0 0.0 1e-06 
3.0 1.724 0 0.0 1e-06 
0.05 1.725 0 0.0 1e-06 
3.0 1.725 0 0.0 1e-06 
0.05 1.726 0 0.0 1e-06 
3.0 1.726 0 0.0 1e-06 
0.05 1.727 0 0.0 1e-06 
3.0 1.727 0 0.0 1e-06 
0.05 1.728 0 0.0 1e-06 
3.0 1.728 0 0.0 1e-06 
0.05 1.729 0 0.0 1e-06 
3.0 1.729 0 0.0 1e-06 
0.05 1.73 0 0.0 1e-06 
3.0 1.73 0 0.0 1e-06 
0.05 1.731 0 0.0 1e-06 
3.0 1.731 0 0.0 1e-06 
0.05 1.732 0 0.0 1e-06 
3.0 1.732 0 0.0 1e-06 
0.05 1.733 0 0.0 1e-06 
3.0 1.733 0 0.0 1e-06 
0.05 1.734 0 0.0 1e-06 
3.0 1.734 0 0.0 1e-06 
0.05 1.735 0 0.0 1e-06 
3.0 1.735 0 0.0 1e-06 
0.05 1.736 0 0.0 1e-06 
3.0 1.736 0 0.0 1e-06 
0.05 1.737 0 0.0 1e-06 
3.0 1.737 0 0.0 1e-06 
0.05 1.738 0 0.0 1e-06 
3.0 1.738 0 0.0 1e-06 
0.05 1.739 0 0.0 1e-06 
3.0 1.739 0 0.0 1e-06 
0.05 1.74 0 0.0 1e-06 
3.0 1.74 0 0.0 1e-06 
0.05 1.741 0 0.0 1e-06 
3.0 1.741 0 0.0 1e-06 
0.05 1.742 0 0.0 1e-06 
3.0 1.742 0 0.0 1e-06 
0.05 1.743 0 0.0 1e-06 
3.0 1.743 0 0.0 1e-06 
0.05 1.744 0 0.0 1e-06 
3.0 1.744 0 0.0 1e-06 
0.05 1.745 0 0.0 1e-06 
3.0 1.745 0 0.0 1e-06 
0.05 1.746 0 0.0 1e-06 
3.0 1.746 0 0.0 1e-06 
0.05 1.747 0 0.0 1e-06 
3.0 1.747 0 0.0 1e-06 
0.05 1.748 0 0.0 1e-06 
3.0 1.748 0 0.0 1e-06 
0.05 1.749 0 0.0 1e-06 
3.0 1.749 0 0.0 1e-06 
0.05 1.75 0 0.0 1e-06 
3.0 1.75 0 0.0 1e-06 
0.05 1.751 0 0.0 1e-06 
3.0 1.751 0 0.0 1e-06 
0.05 1.752 0 0.0 1e-06 
3.0 1.752 0 0.0 1e-06 
0.05 1.753 0 0.0 1e-06 
3.0 1.753 0 0.0 1e-06 
0.05 1.754 0 0.0 1e-06 
3.0 1.754 0 0.0 1e-06 
0.05 1.755 0 0.0 1e-06 
3.0 1.755 0 0.0 1e-06 
0.05 1.756 0 0.0 1e-06 
3.0 1.756 0 0.0 1e-06 
0.05 1.757 0 0.0 1e-06 
3.0 1.757 0 0.0 1e-06 
0.05 1.758 0 0.0 1e-06 
3.0 1.758 0 0.0 1e-06 
0.05 1.759 0 0.0 1e-06 
3.0 1.759 0 0.0 1e-06 
0.05 1.76 0 0.0 1e-06 
3.0 1.76 0 0.0 1e-06 
0.05 1.761 0 0.0 1e-06 
3.0 1.761 0 0.0 1e-06 
0.05 1.762 0 0.0 1e-06 
3.0 1.762 0 0.0 1e-06 
0.05 1.763 0 0.0 1e-06 
3.0 1.763 0 0.0 1e-06 
0.05 1.764 0 0.0 1e-06 
3.0 1.764 0 0.0 1e-06 
0.05 1.765 0 0.0 1e-06 
3.0 1.765 0 0.0 1e-06 
0.05 1.766 0 0.0 1e-06 
3.0 1.766 0 0.0 1e-06 
0.05 1.767 0 0.0 1e-06 
3.0 1.767 0 0.0 1e-06 
0.05 1.768 0 0.0 1e-06 
3.0 1.768 0 0.0 1e-06 
0.05 1.769 0 0.0 1e-06 
3.0 1.769 0 0.0 1e-06 
0.05 1.77 0 0.0 1e-06 
3.0 1.77 0 0.0 1e-06 
0.05 1.771 0 0.0 1e-06 
3.0 1.771 0 0.0 1e-06 
0.05 1.772 0 0.0 1e-06 
3.0 1.772 0 0.0 1e-06 
0.05 1.773 0 0.0 1e-06 
3.0 1.773 0 0.0 1e-06 
0.05 1.774 0 0.0 1e-06 
3.0 1.774 0 0.0 1e-06 
0.05 1.775 0 0.0 1e-06 
3.0 1.775 0 0.0 1e-06 
0.05 1.776 0 0.0 1e-06 
3.0 1.776 0 0.0 1e-06 
0.05 1.777 0 0.0 1e-06 
3.0 1.777 0 0.0 1e-06 
0.05 1.778 0 0.0 1e-06 
3.0 1.778 0 0.0 1e-06 
0.05 1.779 0 0.0 1e-06 
3.0 1.779 0 0.0 1e-06 
0.05 1.78 0 0.0 1e-06 
3.0 1.78 0 0.0 1e-06 
0.05 1.781 0 0.0 1e-06 
3.0 1.781 0 0.0 1e-06 
0.05 1.782 0 0.0 1e-06 
3.0 1.782 0 0.0 1e-06 
0.05 1.783 0 0.0 1e-06 
3.0 1.783 0 0.0 1e-06 
0.05 1.784 0 0.0 1e-06 
3.0 1.784 0 0.0 1e-06 
0.05 1.785 0 0.0 1e-06 
3.0 1.785 0 0.0 1e-06 
0.05 1.786 0 0.0 1e-06 
3.0 1.786 0 0.0 1e-06 
0.05 1.787 0 0.0 1e-06 
3.0 1.787 0 0.0 1e-06 
0.05 1.788 0 0.0 1e-06 
3.0 1.788 0 0.0 1e-06 
0.05 1.789 0 0.0 1e-06 
3.0 1.789 0 0.0 1e-06 
0.05 1.79 0 0.0 1e-06 
3.0 1.79 0 0.0 1e-06 
0.05 1.791 0 0.0 1e-06 
3.0 1.791 0 0.0 1e-06 
0.05 1.792 0 0.0 1e-06 
3.0 1.792 0 0.0 1e-06 
0.05 1.793 0 0.0 1e-06 
3.0 1.793 0 0.0 1e-06 
0.05 1.794 0 0.0 1e-06 
3.0 1.794 0 0.0 1e-06 
0.05 1.795 0 0.0 1e-06 
3.0 1.795 0 0.0 1e-06 
0.05 1.796 0 0.0 1e-06 
3.0 1.796 0 0.0 1e-06 
0.05 1.797 0 0.0 1e-06 
3.0 1.797 0 0.0 1e-06 
0.05 1.798 0 0.0 1e-06 
3.0 1.798 0 0.0 1e-06 
0.05 1.799 0 0.0 1e-06 
3.0 1.799 0 0.0 1e-06 
0.05 1.8 0 0.0 1e-06 
3.0 1.8 0 0.0 1e-06 
0.05 1.801 0 0.0 1e-06 
3.0 1.801 0 0.0 1e-06 
0.05 1.802 0 0.0 1e-06 
3.0 1.802 0 0.0 1e-06 
0.05 1.803 0 0.0 1e-06 
3.0 1.803 0 0.0 1e-06 
0.05 1.804 0 0.0 1e-06 
3.0 1.804 0 0.0 1e-06 
0.05 1.805 0 0.0 1e-06 
3.0 1.805 0 0.0 1e-06 
0.05 1.806 0 0.0 1e-06 
3.0 1.806 0 0.0 1e-06 
0.05 1.807 0 0.0 1e-06 
3.0 1.807 0 0.0 1e-06 
0.05 1.808 0 0.0 1e-06 
3.0 1.808 0 0.0 1e-06 
0.05 1.809 0 0.0 1e-06 
3.0 1.809 0 0.0 1e-06 
0.05 1.81 0 0.0 1e-06 
3.0 1.81 0 0.0 1e-06 
0.05 1.811 0 0.0 1e-06 
3.0 1.811 0 0.0 1e-06 
0.05 1.812 0 0.0 1e-06 
3.0 1.812 0 0.0 1e-06 
0.05 1.813 0 0.0 1e-06 
3.0 1.813 0 0.0 1e-06 
0.05 1.814 0 0.0 1e-06 
3.0 1.814 0 0.0 1e-06 
0.05 1.815 0 0.0 1e-06 
3.0 1.815 0 0.0 1e-06 
0.05 1.816 0 0.0 1e-06 
3.0 1.816 0 0.0 1e-06 
0.05 1.817 0 0.0 1e-06 
3.0 1.817 0 0.0 1e-06 
0.05 1.818 0 0.0 1e-06 
3.0 1.818 0 0.0 1e-06 
0.05 1.819 0 0.0 1e-06 
3.0 1.819 0 0.0 1e-06 
0.05 1.82 0 0.0 1e-06 
3.0 1.82 0 0.0 1e-06 
0.05 1.821 0 0.0 1e-06 
3.0 1.821 0 0.0 1e-06 
0.05 1.822 0 0.0 1e-06 
3.0 1.822 0 0.0 1e-06 
0.05 1.823 0 0.0 1e-06 
3.0 1.823 0 0.0 1e-06 
0.05 1.824 0 0.0 1e-06 
3.0 1.824 0 0.0 1e-06 
0.05 1.825 0 0.0 1e-06 
3.0 1.825 0 0.0 1e-06 
0.05 1.826 0 0.0 1e-06 
3.0 1.826 0 0.0 1e-06 
0.05 1.827 0 0.0 1e-06 
3.0 1.827 0 0.0 1e-06 
0.05 1.828 0 0.0 1e-06 
3.0 1.828 0 0.0 1e-06 
0.05 1.829 0 0.0 1e-06 
3.0 1.829 0 0.0 1e-06 
0.05 1.83 0 0.0 1e-06 
3.0 1.83 0 0.0 1e-06 
0.05 1.831 0 0.0 1e-06 
3.0 1.831 0 0.0 1e-06 
0.05 1.832 0 0.0 1e-06 
3.0 1.832 0 0.0 1e-06 
0.05 1.833 0 0.0 1e-06 
3.0 1.833 0 0.0 1e-06 
0.05 1.834 0 0.0 1e-06 
3.0 1.834 0 0.0 1e-06 
0.05 1.835 0 0.0 1e-06 
3.0 1.835 0 0.0 1e-06 
0.05 1.836 0 0.0 1e-06 
3.0 1.836 0 0.0 1e-06 
0.05 1.837 0 0.0 1e-06 
3.0 1.837 0 0.0 1e-06 
0.05 1.838 0 0.0 1e-06 
3.0 1.838 0 0.0 1e-06 
0.05 1.839 0 0.0 1e-06 
3.0 1.839 0 0.0 1e-06 
0.05 1.84 0 0.0 1e-06 
3.0 1.84 0 0.0 1e-06 
0.05 1.841 0 0.0 1e-06 
3.0 1.841 0 0.0 1e-06 
0.05 1.842 0 0.0 1e-06 
3.0 1.842 0 0.0 1e-06 
0.05 1.843 0 0.0 1e-06 
3.0 1.843 0 0.0 1e-06 
0.05 1.844 0 0.0 1e-06 
3.0 1.844 0 0.0 1e-06 
0.05 1.845 0 0.0 1e-06 
3.0 1.845 0 0.0 1e-06 
0.05 1.846 0 0.0 1e-06 
3.0 1.846 0 0.0 1e-06 
0.05 1.847 0 0.0 1e-06 
3.0 1.847 0 0.0 1e-06 
0.05 1.848 0 0.0 1e-06 
3.0 1.848 0 0.0 1e-06 
0.05 1.849 0 0.0 1e-06 
3.0 1.849 0 0.0 1e-06 
0.05 1.85 0 0.0 1e-06 
3.0 1.85 0 0.0 1e-06 
0.05 1.851 0 0.0 1e-06 
3.0 1.851 0 0.0 1e-06 
0.05 1.852 0 0.0 1e-06 
3.0 1.852 0 0.0 1e-06 
0.05 1.853 0 0.0 1e-06 
3.0 1.853 0 0.0 1e-06 
0.05 1.854 0 0.0 1e-06 
3.0 1.854 0 0.0 1e-06 
0.05 1.855 0 0.0 1e-06 
3.0 1.855 0 0.0 1e-06 
0.05 1.856 0 0.0 1e-06 
3.0 1.856 0 0.0 1e-06 
0.05 1.857 0 0.0 1e-06 
3.0 1.857 0 0.0 1e-06 
0.05 1.858 0 0.0 1e-06 
3.0 1.858 0 0.0 1e-06 
0.05 1.859 0 0.0 1e-06 
3.0 1.859 0 0.0 1e-06 
0.05 1.86 0 0.0 1e-06 
3.0 1.86 0 0.0 1e-06 
0.05 1.861 0 0.0 1e-06 
3.0 1.861 0 0.0 1e-06 
0.05 1.862 0 0.0 1e-06 
3.0 1.862 0 0.0 1e-06 
0.05 1.863 0 0.0 1e-06 
3.0 1.863 0 0.0 1e-06 
0.05 1.864 0 0.0 1e-06 
3.0 1.864 0 0.0 1e-06 
0.05 1.865 0 0.0 1e-06 
3.0 1.865 0 0.0 1e-06 
0.05 1.866 0 0.0 1e-06 
3.0 1.866 0 0.0 1e-06 
0.05 1.867 0 0.0 1e-06 
3.0 1.867 0 0.0 1e-06 
0.05 1.868 0 0.0 1e-06 
3.0 1.868 0 0.0 1e-06 
0.05 1.869 0 0.0 1e-06 
3.0 1.869 0 0.0 1e-06 
0.05 1.87 0 0.0 1e-06 
3.0 1.87 0 0.0 1e-06 
0.05 1.871 0 0.0 1e-06 
3.0 1.871 0 0.0 1e-06 
0.05 1.872 0 0.0 1e-06 
3.0 1.872 0 0.0 1e-06 
0.05 1.873 0 0.0 1e-06 
3.0 1.873 0 0.0 1e-06 
0.05 1.874 0 0.0 1e-06 
3.0 1.874 0 0.0 1e-06 
0.05 1.875 0 0.0 1e-06 
3.0 1.875 0 0.0 1e-06 
0.05 1.876 0 0.0 1e-06 
3.0 1.876 0 0.0 1e-06 
0.05 1.877 0 0.0 1e-06 
3.0 1.877 0 0.0 1e-06 
0.05 1.878 0 0.0 1e-06 
3.0 1.878 0 0.0 1e-06 
0.05 1.879 0 0.0 1e-06 
3.0 1.879 0 0.0 1e-06 
0.05 1.88 0 0.0 1e-06 
3.0 1.88 0 0.0 1e-06 
0.05 1.881 0 0.0 1e-06 
3.0 1.881 0 0.0 1e-06 
0.05 1.882 0 0.0 1e-06 
3.0 1.882 0 0.0 1e-06 
0.05 1.883 0 0.0 1e-06 
3.0 1.883 0 0.0 1e-06 
0.05 1.884 0 0.0 1e-06 
3.0 1.884 0 0.0 1e-06 
0.05 1.885 0 0.0 1e-06 
3.0 1.885 0 0.0 1e-06 
0.05 1.886 0 0.0 1e-06 
3.0 1.886 0 0.0 1e-06 
0.05 1.887 0 0.0 1e-06 
3.0 1.887 0 0.0 1e-06 
0.05 1.888 0 0.0 1e-06 
3.0 1.888 0 0.0 1e-06 
0.05 1.889 0 0.0 1e-06 
3.0 1.889 0 0.0 1e-06 
0.05 1.89 0 0.0 1e-06 
3.0 1.89 0 0.0 1e-06 
0.05 1.891 0 0.0 1e-06 
3.0 1.891 0 0.0 1e-06 
0.05 1.892 0 0.0 1e-06 
3.0 1.892 0 0.0 1e-06 
0.05 1.893 0 0.0 1e-06 
3.0 1.893 0 0.0 1e-06 
0.05 1.894 0 0.0 1e-06 
3.0 1.894 0 0.0 1e-06 
0.05 1.895 0 0.0 1e-06 
3.0 1.895 0 0.0 1e-06 
0.05 1.896 0 0.0 1e-06 
3.0 1.896 0 0.0 1e-06 
0.05 1.897 0 0.0 1e-06 
3.0 1.897 0 0.0 1e-06 
0.05 1.898 0 0.0 1e-06 
3.0 1.898 0 0.0 1e-06 
0.05 1.899 0 0.0 1e-06 
3.0 1.899 0 0.0 1e-06 
0.05 1.9 0 0.0 1e-06 
3.0 1.9 0 0.0 1e-06 
0.05 1.901 0 0.0 1e-06 
3.0 1.901 0 0.0 1e-06 
0.05 1.902 0 0.0 1e-06 
3.0 1.902 0 0.0 1e-06 
0.05 1.903 0 0.0 1e-06 
3.0 1.903 0 0.0 1e-06 
0.05 1.904 0 0.0 1e-06 
3.0 1.904 0 0.0 1e-06 
0.05 1.905 0 0.0 1e-06 
3.0 1.905 0 0.0 1e-06 
0.05 1.906 0 0.0 1e-06 
3.0 1.906 0 0.0 1e-06 
0.05 1.907 0 0.0 1e-06 
3.0 1.907 0 0.0 1e-06 
0.05 1.908 0 0.0 1e-06 
3.0 1.908 0 0.0 1e-06 
0.05 1.909 0 0.0 1e-06 
3.0 1.909 0 0.0 1e-06 
0.05 1.91 0 0.0 1e-06 
3.0 1.91 0 0.0 1e-06 
0.05 1.911 0 0.0 1e-06 
3.0 1.911 0 0.0 1e-06 
0.05 1.912 0 0.0 1e-06 
3.0 1.912 0 0.0 1e-06 
0.05 1.913 0 0.0 1e-06 
3.0 1.913 0 0.0 1e-06 
0.05 1.914 0 0.0 1e-06 
3.0 1.914 0 0.0 1e-06 
0.05 1.915 0 0.0 1e-06 
3.0 1.915 0 0.0 1e-06 
0.05 1.916 0 0.0 1e-06 
3.0 1.916 0 0.0 1e-06 
0.05 1.917 0 0.0 1e-06 
3.0 1.917 0 0.0 1e-06 
0.05 1.918 0 0.0 1e-06 
3.0 1.918 0 0.0 1e-06 
0.05 1.919 0 0.0 1e-06 
3.0 1.919 0 0.0 1e-06 
0.05 1.92 0 0.0 1e-06 
3.0 1.92 0 0.0 1e-06 
0.05 1.921 0 0.0 1e-06 
3.0 1.921 0 0.0 1e-06 
0.05 1.922 0 0.0 1e-06 
3.0 1.922 0 0.0 1e-06 
0.05 1.923 0 0.0 1e-06 
3.0 1.923 0 0.0 1e-06 
0.05 1.924 0 0.0 1e-06 
3.0 1.924 0 0.0 1e-06 
0.05 1.925 0 0.0 1e-06 
3.0 1.925 0 0.0 1e-06 
0.05 1.926 0 0.0 1e-06 
3.0 1.926 0 0.0 1e-06 
0.05 1.927 0 0.0 1e-06 
3.0 1.927 0 0.0 1e-06 
0.05 1.928 0 0.0 1e-06 
3.0 1.928 0 0.0 1e-06 
0.05 1.929 0 0.0 1e-06 
3.0 1.929 0 0.0 1e-06 
0.05 1.93 0 0.0 1e-06 
3.0 1.93 0 0.0 1e-06 
0.05 1.931 0 0.0 1e-06 
3.0 1.931 0 0.0 1e-06 
0.05 1.932 0 0.0 1e-06 
3.0 1.932 0 0.0 1e-06 
0.05 1.933 0 0.0 1e-06 
3.0 1.933 0 0.0 1e-06 
0.05 1.934 0 0.0 1e-06 
3.0 1.934 0 0.0 1e-06 
0.05 1.935 0 0.0 1e-06 
3.0 1.935 0 0.0 1e-06 
0.05 1.936 0 0.0 1e-06 
3.0 1.936 0 0.0 1e-06 
0.05 1.937 0 0.0 1e-06 
3.0 1.937 0 0.0 1e-06 
0.05 1.938 0 0.0 1e-06 
3.0 1.938 0 0.0 1e-06 
0.05 1.939 0 0.0 1e-06 
3.0 1.939 0 0.0 1e-06 
0.05 1.94 0 0.0 1e-06 
3.0 1.94 0 0.0 1e-06 
0.05 1.941 0 0.0 1e-06 
3.0 1.941 0 0.0 1e-06 
0.05 1.942 0 0.0 1e-06 
3.0 1.942 0 0.0 1e-06 
0.05 1.943 0 0.0 1e-06 
3.0 1.943 0 0.0 1e-06 
0.05 1.944 0 0.0 1e-06 
3.0 1.944 0 0.0 1e-06 
0.05 1.945 0 0.0 1e-06 
3.0 1.945 0 0.0 1e-06 
0.05 1.946 0 0.0 1e-06 
3.0 1.946 0 0.0 1e-06 
0.05 1.947 0 0.0 1e-06 
3.0 1.947 0 0.0 1e-06 
0.05 1.948 0 0.0 1e-06 
3.0 1.948 0 0.0 1e-06 
0.05 1.949 0 0.0 1e-06 
3.0 1.949 0 0.0 1e-06 
0.05 1.95 0 0.0 1e-06 
3.0 1.95 0 0.0 1e-06 
0.05 1.951 0 0.0 1e-06 
3.0 1.951 0 0.0 1e-06 
0.05 1.952 0 0.0 1e-06 
3.0 1.952 0 0.0 1e-06 
0.05 1.953 0 0.0 1e-06 
3.0 1.953 0 0.0 1e-06 
0.05 1.954 0 0.0 1e-06 
3.0 1.954 0 0.0 1e-06 
0.05 1.955 0 0.0 1e-06 
3.0 1.955 0 0.0 1e-06 
0.05 1.956 0 0.0 1e-06 
3.0 1.956 0 0.0 1e-06 
0.05 1.957 0 0.0 1e-06 
3.0 1.957 0 0.0 1e-06 
0.05 1.958 0 0.0 1e-06 
3.0 1.958 0 0.0 1e-06 
0.05 1.959 0 0.0 1e-06 
3.0 1.959 0 0.0 1e-06 
0.05 1.96 0 0.0 1e-06 
3.0 1.96 0 0.0 1e-06 
0.05 1.961 0 0.0 1e-06 
3.0 1.961 0 0.0 1e-06 
0.05 1.962 0 0.0 1e-06 
3.0 1.962 0 0.0 1e-06 
0.05 1.963 0 0.0 1e-06 
3.0 1.963 0 0.0 1e-06 
0.05 1.964 0 0.0 1e-06 
3.0 1.964 0 0.0 1e-06 
0.05 1.965 0 0.0 1e-06 
3.0 1.965 0 0.0 1e-06 
0.05 1.966 0 0.0 1e-06 
3.0 1.966 0 0.0 1e-06 
0.05 1.967 0 0.0 1e-06 
3.0 1.967 0 0.0 1e-06 
0.05 1.968 0 0.0 1e-06 
3.0 1.968 0 0.0 1e-06 
0.05 1.969 0 0.0 1e-06 
3.0 1.969 0 0.0 1e-06 
0.05 1.97 0 0.0 1e-06 
3.0 1.97 0 0.0 1e-06 
0.05 1.971 0 0.0 1e-06 
3.0 1.971 0 0.0 1e-06 
0.05 1.972 0 0.0 1e-06 
3.0 1.972 0 0.0 1e-06 
0.05 1.973 0 0.0 1e-06 
3.0 1.973 0 0.0 1e-06 
0.05 1.974 0 0.0 1e-06 
3.0 1.974 0 0.0 1e-06 
0.05 1.975 0 0.0 1e-06 
3.0 1.975 0 0.0 1e-06 
0.05 1.976 0 0.0 1e-06 
3.0 1.976 0 0.0 1e-06 
0.05 1.977 0 0.0 1e-06 
3.0 1.977 0 0.0 1e-06 
0.05 1.978 0 0.0 1e-06 
3.0 1.978 0 0.0 1e-06 
0.05 1.979 0 0.0 1e-06 
3.0 1.979 0 0.0 1e-06 
0.05 1.98 0 0.0 1e-06 
3.0 1.98 0 0.0 1e-06 
0.05 1.981 0 0.0 1e-06 
3.0 1.981 0 0.0 1e-06 
0.05 1.982 0 0.0 1e-06 
3.0 1.982 0 0.0 1e-06 
0.05 1.983 0 0.0 1e-06 
3.0 1.983 0 0.0 1e-06 
0.05 1.984 0 0.0 1e-06 
3.0 1.984 0 0.0 1e-06 
0.05 1.985 0 0.0 1e-06 
3.0 1.985 0 0.0 1e-06 
0.05 1.986 0 0.0 1e-06 
3.0 1.986 0 0.0 1e-06 
0.05 1.987 0 0.0 1e-06 
3.0 1.987 0 0.0 1e-06 
0.05 1.988 0 0.0 1e-06 
3.0 1.988 0 0.0 1e-06 
0.05 1.989 0 0.0 1e-06 
3.0 1.989 0 0.0 1e-06 
0.05 1.99 0 0.0 1e-06 
3.0 1.99 0 0.0 1e-06 
0.05 1.991 0 0.0 1e-06 
3.0 1.991 0 0.0 1e-06 
0.05 1.992 0 0.0 1e-06 
3.0 1.992 0 0.0 1e-06 
0.05 1.993 0 0.0 1e-06 
3.0 1.993 0 0.0 1e-06 
0.05 1.994 0 0.0 1e-06 
3.0 1.994 0 0.0 1e-06 
0.05 1.995 0 0.0 1e-06 
3.0 1.995 0 0.0 1e-06 
0.05 1.996 0 0.0 1e-06 
3.0 1.996 0 0.0 1e-06 
0.05 1.997 0 0.0 1e-06 
3.0 1.997 0 0.0 1e-06 
0.05 1.998 0 0.0 1e-06 
3.0 1.998 0 0.0 1e-06 
0.05 1.999 0 0.0 1e-06 
3.0 1.999 0 0.0 1e-06 
0.05 2.0 0 0.0 1e-06 
3.0 2.0 0 0.0 1e-06 
0.05 2.001 0 0.0 1e-06 
3.0 2.001 0 0.0 1e-06 
0.05 2.002 0 0.0 1e-06 
3.0 2.002 0 0.0 1e-06 
0.05 2.003 0 0.0 1e-06 
3.0 2.003 0 0.0 1e-06 
0.05 2.004 0 0.0 1e-06 
3.0 2.004 0 0.0 1e-06 
0.05 2.005 0 0.0 1e-06 
3.0 2.005 0 0.0 1e-06 
0.05 2.006 0 0.0 1e-06 
3.0 2.006 0 0.0 1e-06 
0.05 2.007 0 0.0 1e-06 
3.0 2.007 0 0.0 1e-06 
0.05 2.008 0 0.0 1e-06 
3.0 2.008 0 0.0 1e-06 
0.05 2.009 0 0.0 1e-06 
3.0 2.009 0 0.0 1e-06 
0.05 2.01 0 0.0 1e-06 
3.0 2.01 0 0.0 1e-06 
0.05 2.011 0 0.0 1e-06 
3.0 2.011 0 0.0 1e-06 
0.05 2.012 0 0.0 1e-06 
3.0 2.012 0 0.0 1e-06 
0.05 2.013 0 0.0 1e-06 
3.0 2.013 0 0.0 1e-06 
0.05 2.014 0 0.0 1e-06 
3.0 2.014 0 0.0 1e-06 
0.05 2.015 0 0.0 1e-06 
3.0 2.015 0 0.0 1e-06 
0.05 2.016 0 0.0 1e-06 
3.0 2.016 0 0.0 1e-06 
0.05 2.017 0 0.0 1e-06 
3.0 2.017 0 0.0 1e-06 
0.05 2.018 0 0.0 1e-06 
3.0 2.018 0 0.0 1e-06 
0.05 2.019 0 0.0 1e-06 
3.0 2.019 0 0.0 1e-06 
0.05 2.02 0 0.0 1e-06 
3.0 2.02 0 0.0 1e-06 
0.05 2.021 0 0.0 1e-06 
3.0 2.021 0 0.0 1e-06 
0.05 2.022 0 0.0 1e-06 
3.0 2.022 0 0.0 1e-06 
0.05 2.023 0 0.0 1e-06 
3.0 2.023 0 0.0 1e-06 
0.05 2.024 0 0.0 1e-06 
3.0 2.024 0 0.0 1e-06 
0.05 2.025 0 0.0 1e-06 
3.0 2.025 0 0.0 1e-06 
0.05 2.026 0 0.0 1e-06 
3.0 2.026 0 0.0 1e-06 
0.05 2.027 0 0.0 1e-06 
3.0 2.027 0 0.0 1e-06 
0.05 2.028 0 0.0 1e-06 
3.0 2.028 0 0.0 1e-06 
0.05 2.029 0 0.0 1e-06 
3.0 2.029 0 0.0 1e-06 
0.05 2.03 0 0.0 1e-06 
3.0 2.03 0 0.0 1e-06 
0.05 2.031 0 0.0 1e-06 
3.0 2.031 0 0.0 1e-06 
0.05 2.032 0 0.0 1e-06 
3.0 2.032 0 0.0 1e-06 
0.05 2.033 0 0.0 1e-06 
3.0 2.033 0 0.0 1e-06 
0.05 2.034 0 0.0 1e-06 
3.0 2.034 0 0.0 1e-06 
0.05 2.035 0 0.0 1e-06 
3.0 2.035 0 0.0 1e-06 
0.05 2.036 0 0.0 1e-06 
3.0 2.036 0 0.0 1e-06 
0.05 2.037 0 0.0 1e-06 
3.0 2.037 0 0.0 1e-06 
0.05 2.038 0 0.0 1e-06 
3.0 2.038 0 0.0 1e-06 
0.05 2.039 0 0.0 1e-06 
3.0 2.039 0 0.0 1e-06 
0.05 2.04 0 0.0 1e-06 
3.0 2.04 0 0.0 1e-06 
0.05 2.041 0 0.0 1e-06 
3.0 2.041 0 0.0 1e-06 
0.05 2.042 0 0.0 1e-06 
3.0 2.042 0 0.0 1e-06 
0.05 2.043 0 0.0 1e-06 
3.0 2.043 0 0.0 1e-06 
0.05 2.044 0 0.0 1e-06 
3.0 2.044 0 0.0 1e-06 
0.05 2.045 0 0.0 1e-06 
3.0 2.045 0 0.0 1e-06 
0.05 2.046 0 0.0 1e-06 
3.0 2.046 0 0.0 1e-06 
0.05 2.047 0 0.0 1e-06 
3.0 2.047 0 0.0 1e-06 
0.05 2.048 0 0.0 1e-06 
3.0 2.048 0 0.0 1e-06 
0.05 2.049 0 0.0 1e-06 
3.0 2.049 0 0.0 1e-06 
0.05 2.05 0 0.0 1e-06 
3.0 2.05 0 0.0 1e-06 
0.05 2.051 0 0.0 1e-06 
3.0 2.051 0 0.0 1e-06 
0.05 2.052 0 0.0 1e-06 
3.0 2.052 0 0.0 1e-06 
0.05 2.053 0 0.0 1e-06 
3.0 2.053 0 0.0 1e-06 
0.05 2.054 0 0.0 1e-06 
3.0 2.054 0 0.0 1e-06 
0.05 2.055 0 0.0 1e-06 
3.0 2.055 0 0.0 1e-06 
0.05 2.056 0 0.0 1e-06 
3.0 2.056 0 0.0 1e-06 
0.05 2.057 0 0.0 1e-06 
3.0 2.057 0 0.0 1e-06 
0.05 2.058 0 0.0 1e-06 
3.0 2.058 0 0.0 1e-06 
0.05 2.059 0 0.0 1e-06 
3.0 2.059 0 0.0 1e-06 
0.05 2.06 0 0.0 1e-06 
3.0 2.06 0 0.0 1e-06 
0.05 2.061 0 0.0 1e-06 
3.0 2.061 0 0.0 1e-06 
0.05 2.062 0 0.0 1e-06 
3.0 2.062 0 0.0 1e-06 
0.05 2.063 0 0.0 1e-06 
3.0 2.063 0 0.0 1e-06 
0.05 2.064 0 0.0 1e-06 
3.0 2.064 0 0.0 1e-06 
0.05 2.065 0 0.0 1e-06 
3.0 2.065 0 0.0 1e-06 
0.05 2.066 0 0.0 1e-06 
3.0 2.066 0 0.0 1e-06 
0.05 2.067 0 0.0 1e-06 
3.0 2.067 0 0.0 1e-06 
0.05 2.068 0 0.0 1e-06 
3.0 2.068 0 0.0 1e-06 
0.05 2.069 0 0.0 1e-06 
3.0 2.069 0 0.0 1e-06 
0.05 2.07 0 0.0 1e-06 
3.0 2.07 0 0.0 1e-06 
0.05 2.071 0 0.0 1e-06 
3.0 2.071 0 0.0 1e-06 
0.05 2.072 0 0.0 1e-06 
3.0 2.072 0 0.0 1e-06 
0.05 2.073 0 0.0 1e-06 
3.0 2.073 0 0.0 1e-06 
0.05 2.074 0 0.0 1e-06 
3.0 2.074 0 0.0 1e-06 
0.05 2.075 0 0.0 1e-06 
3.0 2.075 0 0.0 1e-06 
0.05 2.076 0 0.0 1e-06 
3.0 2.076 0 0.0 1e-06 
0.05 2.077 0 0.0 1e-06 
3.0 2.077 0 0.0 1e-06 
0.05 2.078 0 0.0 1e-06 
3.0 2.078 0 0.0 1e-06 
0.05 2.079 0 0.0 1e-06 
3.0 2.079 0 0.0 1e-06 
0.05 2.08 0 0.0 1e-06 
3.0 2.08 0 0.0 1e-06 
0.05 2.081 0 0.0 1e-06 
3.0 2.081 0 0.0 1e-06 
0.05 2.082 0 0.0 1e-06 
3.0 2.082 0 0.0 1e-06 
0.05 2.083 0 0.0 1e-06 
3.0 2.083 0 0.0 1e-06 
0.05 2.084 0 0.0 1e-06 
3.0 2.084 0 0.0 1e-06 
0.05 2.085 0 0.0 1e-06 
3.0 2.085 0 0.0 1e-06 
0.05 2.086 0 0.0 1e-06 
3.0 2.086 0 0.0 1e-06 
0.05 2.087 0 0.0 1e-06 
3.0 2.087 0 0.0 1e-06 
0.05 2.088 0 0.0 1e-06 
3.0 2.088 0 0.0 1e-06 
0.05 2.089 0 0.0 1e-06 
3.0 2.089 0 0.0 1e-06 
0.05 2.09 0 0.0 1e-06 
3.0 2.09 0 0.0 1e-06 
0.05 2.091 0 0.0 1e-06 
3.0 2.091 0 0.0 1e-06 
0.05 2.092 0 0.0 1e-06 
3.0 2.092 0 0.0 1e-06 
0.05 2.093 0 0.0 1e-06 
3.0 2.093 0 0.0 1e-06 
0.05 2.094 0 0.0 1e-06 
3.0 2.094 0 0.0 1e-06 
0.05 2.095 0 0.0 1e-06 
3.0 2.095 0 0.0 1e-06 
0.05 2.096 0 0.0 1e-06 
3.0 2.096 0 0.0 1e-06 
0.05 2.097 0 0.0 1e-06 
3.0 2.097 0 0.0 1e-06 
0.05 2.098 0 0.0 1e-06 
3.0 2.098 0 0.0 1e-06 
0.05 2.099 0 0.0 1e-06 
3.0 2.099 0 0.0 1e-06 
0.05 2.1 0 0.0 1e-06 
3.0 2.1 0 0.0 1e-06 
0.05 2.101 0 0.0 1e-06 
3.0 2.101 0 0.0 1e-06 
0.05 2.102 0 0.0 1e-06 
3.0 2.102 0 0.0 1e-06 
0.05 2.103 0 0.0 1e-06 
3.0 2.103 0 0.0 1e-06 
0.05 2.104 0 0.0 1e-06 
3.0 2.104 0 0.0 1e-06 
0.05 2.105 0 0.0 1e-06 
3.0 2.105 0 0.0 1e-06 
0.05 2.106 0 0.0 1e-06 
3.0 2.106 0 0.0 1e-06 
0.05 2.107 0 0.0 1e-06 
3.0 2.107 0 0.0 1e-06 
0.05 2.108 0 0.0 1e-06 
3.0 2.108 0 0.0 1e-06 
0.05 2.109 0 0.0 1e-06 
3.0 2.109 0 0.0 1e-06 
0.05 2.11 0 0.0 1e-06 
3.0 2.11 0 0.0 1e-06 
0.05 2.111 0 0.0 1e-06 
3.0 2.111 0 0.0 1e-06 
0.05 2.112 0 0.0 1e-06 
3.0 2.112 0 0.0 1e-06 
0.05 2.113 0 0.0 1e-06 
3.0 2.113 0 0.0 1e-06 
0.05 2.114 0 0.0 1e-06 
3.0 2.114 0 0.0 1e-06 
0.05 2.115 0 0.0 1e-06 
3.0 2.115 0 0.0 1e-06 
0.05 2.116 0 0.0 1e-06 
3.0 2.116 0 0.0 1e-06 
0.05 2.117 0 0.0 1e-06 
3.0 2.117 0 0.0 1e-06 
0.05 2.118 0 0.0 1e-06 
3.0 2.118 0 0.0 1e-06 
0.05 2.119 0 0.0 1e-06 
3.0 2.119 0 0.0 1e-06 
0.05 2.12 0 0.0 1e-06 
3.0 2.12 0 0.0 1e-06 
0.05 2.121 0 0.0 1e-06 
3.0 2.121 0 0.0 1e-06 
0.05 2.122 0 0.0 1e-06 
3.0 2.122 0 0.0 1e-06 
0.05 2.123 0 0.0 1e-06 
3.0 2.123 0 0.0 1e-06 
0.05 2.124 0 0.0 1e-06 
3.0 2.124 0 0.0 1e-06 
0.05 2.125 0 0.0 1e-06 
3.0 2.125 0 0.0 1e-06 
0.05 2.126 0 0.0 1e-06 
3.0 2.126 0 0.0 1e-06 
0.05 2.127 0 0.0 1e-06 
3.0 2.127 0 0.0 1e-06 
0.05 2.128 0 0.0 1e-06 
3.0 2.128 0 0.0 1e-06 
0.05 2.129 0 0.0 1e-06 
3.0 2.129 0 0.0 1e-06 
0.05 2.13 0 0.0 1e-06 
3.0 2.13 0 0.0 1e-06 
0.05 2.131 0 0.0 1e-06 
3.0 2.131 0 0.0 1e-06 
0.05 2.132 0 0.0 1e-06 
3.0 2.132 0 0.0 1e-06 
0.05 2.133 0 0.0 1e-06 
3.0 2.133 0 0.0 1e-06 
0.05 2.134 0 0.0 1e-06 
3.0 2.134 0 0.0 1e-06 
0.05 2.135 0 0.0 1e-06 
3.0 2.135 0 0.0 1e-06 
0.05 2.136 0 0.0 1e-06 
3.0 2.136 0 0.0 1e-06 
0.05 2.137 0 0.0 1e-06 
3.0 2.137 0 0.0 1e-06 
0.05 2.138 0 0.0 1e-06 
3.0 2.138 0 0.0 1e-06 
0.05 2.139 0 0.0 1e-06 
3.0 2.139 0 0.0 1e-06 
0.05 2.14 0 0.0 1e-06 
3.0 2.14 0 0.0 1e-06 
0.05 2.141 0 0.0 1e-06 
3.0 2.141 0 0.0 1e-06 
0.05 2.142 0 0.0 1e-06 
3.0 2.142 0 0.0 1e-06 
0.05 2.143 0 0.0 1e-06 
3.0 2.143 0 0.0 1e-06 
0.05 2.144 0 0.0 1e-06 
3.0 2.144 0 0.0 1e-06 
0.05 2.145 0 0.0 1e-06 
3.0 2.145 0 0.0 1e-06 
0.05 2.146 0 0.0 1e-06 
3.0 2.146 0 0.0 1e-06 
0.05 2.147 0 0.0 1e-06 
3.0 2.147 0 0.0 1e-06 
0.05 2.148 0 0.0 1e-06 
3.0 2.148 0 0.0 1e-06 
0.05 2.149 0 0.0 1e-06 
3.0 2.149 0 0.0 1e-06 
0.05 2.15 0 0.0 1e-06 
3.0 2.15 0 0.0 1e-06 
0.05 2.151 0 0.0 1e-06 
3.0 2.151 0 0.0 1e-06 
0.05 2.152 0 0.0 1e-06 
3.0 2.152 0 0.0 1e-06 
0.05 2.153 0 0.0 1e-06 
3.0 2.153 0 0.0 1e-06 
0.05 2.154 0 0.0 1e-06 
3.0 2.154 0 0.0 1e-06 
0.05 2.155 0 0.0 1e-06 
3.0 2.155 0 0.0 1e-06 
0.05 2.156 0 0.0 1e-06 
3.0 2.156 0 0.0 1e-06 
0.05 2.157 0 0.0 1e-06 
3.0 2.157 0 0.0 1e-06 
0.05 2.158 0 0.0 1e-06 
3.0 2.158 0 0.0 1e-06 
0.05 2.159 0 0.0 1e-06 
3.0 2.159 0 0.0 1e-06 
0.05 2.16 0 0.0 1e-06 
3.0 2.16 0 0.0 1e-06 
0.05 2.161 0 0.0 1e-06 
3.0 2.161 0 0.0 1e-06 
0.05 2.162 0 0.0 1e-06 
3.0 2.162 0 0.0 1e-06 
0.05 2.163 0 0.0 1e-06 
3.0 2.163 0 0.0 1e-06 
0.05 2.164 0 0.0 1e-06 
3.0 2.164 0 0.0 1e-06 
0.05 2.165 0 0.0 1e-06 
3.0 2.165 0 0.0 1e-06 
0.05 2.166 0 0.0 1e-06 
3.0 2.166 0 0.0 1e-06 
0.05 2.167 0 0.0 1e-06 
3.0 2.167 0 0.0 1e-06 
0.05 2.168 0 0.0 1e-06 
3.0 2.168 0 0.0 1e-06 
0.05 2.169 0 0.0 1e-06 
3.0 2.169 0 0.0 1e-06 
0.05 2.17 0 0.0 1e-06 
3.0 2.17 0 0.0 1e-06 
0.05 2.171 0 0.0 1e-06 
3.0 2.171 0 0.0 1e-06 
0.05 2.172 0 0.0 1e-06 
3.0 2.172 0 0.0 1e-06 
0.05 2.173 0 0.0 1e-06 
3.0 2.173 0 0.0 1e-06 
0.05 2.174 0 0.0 1e-06 
3.0 2.174 0 0.0 1e-06 
0.05 2.175 0 0.0 1e-06 
3.0 2.175 0 0.0 1e-06 
0.05 2.176 0 0.0 1e-06 
3.0 2.176 0 0.0 1e-06 
0.05 2.177 0 0.0 1e-06 
3.0 2.177 0 0.0 1e-06 
0.05 2.178 0 0.0 1e-06 
3.0 2.178 0 0.0 1e-06 
0.05 2.179 0 0.0 1e-06 
3.0 2.179 0 0.0 1e-06 
0.05 2.18 0 0.0 1e-06 
3.0 2.18 0 0.0 1e-06 
0.05 2.181 0 0.0 1e-06 
3.0 2.181 0 0.0 1e-06 
0.05 2.182 0 0.0 1e-06 
3.0 2.182 0 0.0 1e-06 
0.05 2.183 0 0.0 1e-06 
3.0 2.183 0 0.0 1e-06 
0.05 2.184 0 0.0 1e-06 
3.0 2.184 0 0.0 1e-06 
0.05 2.185 0 0.0 1e-06 
3.0 2.185 0 0.0 1e-06 
0.05 2.186 0 0.0 1e-06 
3.0 2.186 0 0.0 1e-06 
0.05 2.187 0 0.0 1e-06 
3.0 2.187 0 0.0 1e-06 
0.05 2.188 0 0.0 1e-06 
3.0 2.188 0 0.0 1e-06 
0.05 2.189 0 0.0 1e-06 
3.0 2.189 0 0.0 1e-06 
0.05 2.19 0 0.0 1e-06 
3.0 2.19 0 0.0 1e-06 
0.05 2.191 0 0.0 1e-06 
3.0 2.191 0 0.0 1e-06 
0.05 2.192 0 0.0 1e-06 
3.0 2.192 0 0.0 1e-06 
0.05 2.193 0 0.0 1e-06 
3.0 2.193 0 0.0 1e-06 
0.05 2.194 0 0.0 1e-06 
3.0 2.194 0 0.0 1e-06 
0.05 2.195 0 0.0 1e-06 
3.0 2.195 0 0.0 1e-06 
0.05 2.196 0 0.0 1e-06 
3.0 2.196 0 0.0 1e-06 
0.05 2.197 0 0.0 1e-06 
3.0 2.197 0 0.0 1e-06 
0.05 2.198 0 0.0 1e-06 
3.0 2.198 0 0.0 1e-06 
0.05 2.199 0 0.0 1e-06 
3.0 2.199 0 0.0 1e-06 
0.05 2.2 0 0.0 1e-06 
3.0 2.2 0 0.0 1e-06 
0.05 2.201 0 0.0 1e-06 
3.0 2.201 0 0.0 1e-06 
0.05 2.202 0 0.0 1e-06 
3.0 2.202 0 0.0 1e-06 
0.05 2.203 0 0.0 1e-06 
3.0 2.203 0 0.0 1e-06 
0.05 2.204 0 0.0 1e-06 
3.0 2.204 0 0.0 1e-06 
0.05 2.205 0 0.0 1e-06 
3.0 2.205 0 0.0 1e-06 
0.05 2.206 0 0.0 1e-06 
3.0 2.206 0 0.0 1e-06 
0.05 2.207 0 0.0 1e-06 
3.0 2.207 0 0.0 1e-06 
0.05 2.208 0 0.0 1e-06 
3.0 2.208 0 0.0 1e-06 
0.05 2.209 0 0.0 1e-06 
3.0 2.209 0 0.0 1e-06 
0.05 2.21 0 0.0 1e-06 
3.0 2.21 0 0.0 1e-06 
0.05 2.211 0 0.0 1e-06 
3.0 2.211 0 0.0 1e-06 
0.05 2.212 0 0.0 1e-06 
3.0 2.212 0 0.0 1e-06 
0.05 2.213 0 0.0 1e-06 
3.0 2.213 0 0.0 1e-06 
0.05 2.214 0 0.0 1e-06 
3.0 2.214 0 0.0 1e-06 
0.05 2.215 0 0.0 1e-06 
3.0 2.215 0 0.0 1e-06 
0.05 2.216 0 0.0 1e-06 
3.0 2.216 0 0.0 1e-06 
0.05 2.217 0 0.0 1e-06 
3.0 2.217 0 0.0 1e-06 
0.05 2.218 0 0.0 1e-06 
3.0 2.218 0 0.0 1e-06 
0.05 2.219 0 0.0 1e-06 
3.0 2.219 0 0.0 1e-06 
0.05 2.22 0 0.0 1e-06 
3.0 2.22 0 0.0 1e-06 
0.05 2.221 0 0.0 1e-06 
3.0 2.221 0 0.0 1e-06 
0.05 2.222 0 0.0 1e-06 
3.0 2.222 0 0.0 1e-06 
0.05 2.223 0 0.0 1e-06 
3.0 2.223 0 0.0 1e-06 
0.05 2.224 0 0.0 1e-06 
3.0 2.224 0 0.0 1e-06 
0.05 2.225 0 0.0 1e-06 
3.0 2.225 0 0.0 1e-06 
0.05 2.226 0 0.0 1e-06 
3.0 2.226 0 0.0 1e-06 
0.05 2.227 0 0.0 1e-06 
3.0 2.227 0 0.0 1e-06 
0.05 2.228 0 0.0 1e-06 
3.0 2.228 0 0.0 1e-06 
0.05 2.229 0 0.0 1e-06 
3.0 2.229 0 0.0 1e-06 
0.05 2.23 0 0.0 1e-06 
3.0 2.23 0 0.0 1e-06 
0.05 2.231 0 0.0 1e-06 
3.0 2.231 0 0.0 1e-06 
0.05 2.232 0 0.0 1e-06 
3.0 2.232 0 0.0 1e-06 
0.05 2.233 0 0.0 1e-06 
3.0 2.233 0 0.0 1e-06 
0.05 2.234 0 0.0 1e-06 
3.0 2.234 0 0.0 1e-06 
0.05 2.235 0 0.0 1e-06 
3.0 2.235 0 0.0 1e-06 
0.05 2.236 0 0.0 1e-06 
3.0 2.236 0 0.0 1e-06 
0.05 2.237 0 0.0 1e-06 
3.0 2.237 0 0.0 1e-06 
0.05 2.238 0 0.0 1e-06 
3.0 2.238 0 0.0 1e-06 
0.05 2.239 0 0.0 1e-06 
3.0 2.239 0 0.0 1e-06 
0.05 2.24 0 0.0 1e-06 
3.0 2.24 0 0.0 1e-06 
0.05 2.241 0 0.0 1e-06 
3.0 2.241 0 0.0 1e-06 
0.05 2.242 0 0.0 1e-06 
3.0 2.242 0 0.0 1e-06 
0.05 2.243 0 0.0 1e-06 
3.0 2.243 0 0.0 1e-06 
0.05 2.244 0 0.0 1e-06 
3.0 2.244 0 0.0 1e-06 
0.05 2.245 0 0.0 1e-06 
3.0 2.245 0 0.0 1e-06 
0.05 2.246 0 0.0 1e-06 
3.0 2.246 0 0.0 1e-06 
0.05 2.247 0 0.0 1e-06 
3.0 2.247 0 0.0 1e-06 
0.05 2.248 0 0.0 1e-06 
3.0 2.248 0 0.0 1e-06 
0.05 2.249 0 0.0 1e-06 
3.0 2.249 0 0.0 1e-06 
0.05 2.25 0 0.0 1e-06 
3.0 2.25 0 0.0 1e-06 
0.05 2.251 0 0.0 1e-06 
3.0 2.251 0 0.0 1e-06 
0.05 2.252 0 0.0 1e-06 
3.0 2.252 0 0.0 1e-06 
0.05 2.253 0 0.0 1e-06 
3.0 2.253 0 0.0 1e-06 
0.05 2.254 0 0.0 1e-06 
3.0 2.254 0 0.0 1e-06 
0.05 2.255 0 0.0 1e-06 
3.0 2.255 0 0.0 1e-06 
0.05 2.256 0 0.0 1e-06 
3.0 2.256 0 0.0 1e-06 
0.05 2.257 0 0.0 1e-06 
3.0 2.257 0 0.0 1e-06 
0.05 2.258 0 0.0 1e-06 
3.0 2.258 0 0.0 1e-06 
0.05 2.259 0 0.0 1e-06 
3.0 2.259 0 0.0 1e-06 
0.05 2.26 0 0.0 1e-06 
3.0 2.26 0 0.0 1e-06 
0.05 2.261 0 0.0 1e-06 
3.0 2.261 0 0.0 1e-06 
0.05 2.262 0 0.0 1e-06 
3.0 2.262 0 0.0 1e-06 
0.05 2.263 0 0.0 1e-06 
3.0 2.263 0 0.0 1e-06 
0.05 2.264 0 0.0 1e-06 
3.0 2.264 0 0.0 1e-06 
0.05 2.265 0 0.0 1e-06 
3.0 2.265 0 0.0 1e-06 
0.05 2.266 0 0.0 1e-06 
3.0 2.266 0 0.0 1e-06 
0.05 2.267 0 0.0 1e-06 
3.0 2.267 0 0.0 1e-06 
0.05 2.268 0 0.0 1e-06 
3.0 2.268 0 0.0 1e-06 
0.05 2.269 0 0.0 1e-06 
3.0 2.269 0 0.0 1e-06 
0.05 2.27 0 0.0 1e-06 
3.0 2.27 0 0.0 1e-06 
0.05 2.271 0 0.0 1e-06 
3.0 2.271 0 0.0 1e-06 
0.05 2.272 0 0.0 1e-06 
3.0 2.272 0 0.0 1e-06 
0.05 2.273 0 0.0 1e-06 
3.0 2.273 0 0.0 1e-06 
0.05 2.274 0 0.0 1e-06 
3.0 2.274 0 0.0 1e-06 
0.05 2.275 0 0.0 1e-06 
3.0 2.275 0 0.0 1e-06 
0.05 2.276 0 0.0 1e-06 
3.0 2.276 0 0.0 1e-06 
0.05 2.277 0 0.0 1e-06 
3.0 2.277 0 0.0 1e-06 
0.05 2.278 0 0.0 1e-06 
3.0 2.278 0 0.0 1e-06 
0.05 2.279 0 0.0 1e-06 
3.0 2.279 0 0.0 1e-06 
0.05 2.28 0 0.0 1e-06 
3.0 2.28 0 0.0 1e-06 
0.05 2.281 0 0.0 1e-06 
3.0 2.281 0 0.0 1e-06 
0.05 2.282 0 0.0 1e-06 
3.0 2.282 0 0.0 1e-06 
0.05 2.283 0 0.0 1e-06 
3.0 2.283 0 0.0 1e-06 
0.05 2.284 0 0.0 1e-06 
3.0 2.284 0 0.0 1e-06 
0.05 2.285 0 0.0 1e-06 
3.0 2.285 0 0.0 1e-06 
0.05 2.286 0 0.0 1e-06 
3.0 2.286 0 0.0 1e-06 
0.05 2.287 0 0.0 1e-06 
3.0 2.287 0 0.0 1e-06 
0.05 2.288 0 0.0 1e-06 
3.0 2.288 0 0.0 1e-06 
0.05 2.289 0 0.0 1e-06 
3.0 2.289 0 0.0 1e-06 
0.05 2.29 0 0.0 1e-06 
3.0 2.29 0 0.0 1e-06 
0.05 2.291 0 0.0 1e-06 
3.0 2.291 0 0.0 1e-06 
0.05 2.292 0 0.0 1e-06 
3.0 2.292 0 0.0 1e-06 
0.05 2.293 0 0.0 1e-06 
3.0 2.293 0 0.0 1e-06 
0.05 2.294 0 0.0 1e-06 
3.0 2.294 0 0.0 1e-06 
0.05 2.295 0 0.0 1e-06 
3.0 2.295 0 0.0 1e-06 
0.05 2.296 0 0.0 1e-06 
3.0 2.296 0 0.0 1e-06 
0.05 2.297 0 0.0 1e-06 
3.0 2.297 0 0.0 1e-06 
0.05 2.298 0 0.0 1e-06 
3.0 2.298 0 0.0 1e-06 
0.05 2.299 0 0.0 1e-06 
3.0 2.299 0 0.0 1e-06 
0.05 2.3 0 0.0 1e-06 
3.0 2.3 0 0.0 1e-06 
0.05 2.301 0 0.0 1e-06 
3.0 2.301 0 0.0 1e-06 
0.05 2.302 0 0.0 1e-06 
3.0 2.302 0 0.0 1e-06 
0.05 2.303 0 0.0 1e-06 
3.0 2.303 0 0.0 1e-06 
0.05 2.304 0 0.0 1e-06 
3.0 2.304 0 0.0 1e-06 
0.05 2.305 0 0.0 1e-06 
3.0 2.305 0 0.0 1e-06 
0.05 2.306 0 0.0 1e-06 
3.0 2.306 0 0.0 1e-06 
0.05 2.307 0 0.0 1e-06 
3.0 2.307 0 0.0 1e-06 
0.05 2.308 0 0.0 1e-06 
3.0 2.308 0 0.0 1e-06 
0.05 2.309 0 0.0 1e-06 
3.0 2.309 0 0.0 1e-06 
0.05 2.31 0 0.0 1e-06 
3.0 2.31 0 0.0 1e-06 
0.05 2.311 0 0.0 1e-06 
3.0 2.311 0 0.0 1e-06 
0.05 2.312 0 0.0 1e-06 
3.0 2.312 0 0.0 1e-06 
0.05 2.313 0 0.0 1e-06 
3.0 2.313 0 0.0 1e-06 
0.05 2.314 0 0.0 1e-06 
3.0 2.314 0 0.0 1e-06 
0.05 2.315 0 0.0 1e-06 
3.0 2.315 0 0.0 1e-06 
0.05 2.316 0 0.0 1e-06 
3.0 2.316 0 0.0 1e-06 
0.05 2.317 0 0.0 1e-06 
3.0 2.317 0 0.0 1e-06 
0.05 2.318 0 0.0 1e-06 
3.0 2.318 0 0.0 1e-06 
0.05 2.319 0 0.0 1e-06 
3.0 2.319 0 0.0 1e-06 
0.05 2.32 0 0.0 1e-06 
3.0 2.32 0 0.0 1e-06 
0.05 2.321 0 0.0 1e-06 
3.0 2.321 0 0.0 1e-06 
0.05 2.322 0 0.0 1e-06 
3.0 2.322 0 0.0 1e-06 
0.05 2.323 0 0.0 1e-06 
3.0 2.323 0 0.0 1e-06 
0.05 2.324 0 0.0 1e-06 
3.0 2.324 0 0.0 1e-06 
0.05 2.325 0 0.0 1e-06 
3.0 2.325 0 0.0 1e-06 
0.05 2.326 0 0.0 1e-06 
3.0 2.326 0 0.0 1e-06 
0.05 2.327 0 0.0 1e-06 
3.0 2.327 0 0.0 1e-06 
0.05 2.328 0 0.0 1e-06 
3.0 2.328 0 0.0 1e-06 
0.05 2.329 0 0.0 1e-06 
3.0 2.329 0 0.0 1e-06 
0.05 2.33 0 0.0 1e-06 
3.0 2.33 0 0.0 1e-06 
0.05 2.331 0 0.0 1e-06 
3.0 2.331 0 0.0 1e-06 
0.05 2.332 0 0.0 1e-06 
3.0 2.332 0 0.0 1e-06 
0.05 2.333 0 0.0 1e-06 
3.0 2.333 0 0.0 1e-06 
0.05 2.334 0 0.0 1e-06 
3.0 2.334 0 0.0 1e-06 
0.05 2.335 0 0.0 1e-06 
3.0 2.335 0 0.0 1e-06 
0.05 2.336 0 0.0 1e-06 
3.0 2.336 0 0.0 1e-06 
0.05 2.337 0 0.0 1e-06 
3.0 2.337 0 0.0 1e-06 
0.05 2.338 0 0.0 1e-06 
3.0 2.338 0 0.0 1e-06 
0.05 2.339 0 0.0 1e-06 
3.0 2.339 0 0.0 1e-06 
0.05 2.34 0 0.0 1e-06 
3.0 2.34 0 0.0 1e-06 
0.05 2.341 0 0.0 1e-06 
3.0 2.341 0 0.0 1e-06 
0.05 2.342 0 0.0 1e-06 
3.0 2.342 0 0.0 1e-06 
0.05 2.343 0 0.0 1e-06 
3.0 2.343 0 0.0 1e-06 
0.05 2.344 0 0.0 1e-06 
3.0 2.344 0 0.0 1e-06 
0.05 2.345 0 0.0 1e-06 
3.0 2.345 0 0.0 1e-06 
0.05 2.346 0 0.0 1e-06 
3.0 2.346 0 0.0 1e-06 
0.05 2.347 0 0.0 1e-06 
3.0 2.347 0 0.0 1e-06 
0.05 2.348 0 0.0 1e-06 
3.0 2.348 0 0.0 1e-06 
0.05 2.349 0 0.0 1e-06 
3.0 2.349 0 0.0 1e-06 
0.05 2.35 0 0.0 1e-06 
3.0 2.35 0 0.0 1e-06 
0.05 2.351 0 0.0 1e-06 
3.0 2.351 0 0.0 1e-06 
0.05 2.352 0 0.0 1e-06 
3.0 2.352 0 0.0 1e-06 
0.05 2.353 0 0.0 1e-06 
3.0 2.353 0 0.0 1e-06 
0.05 2.354 0 0.0 1e-06 
3.0 2.354 0 0.0 1e-06 
0.05 2.355 0 0.0 1e-06 
3.0 2.355 0 0.0 1e-06 
0.05 2.356 0 0.0 1e-06 
3.0 2.356 0 0.0 1e-06 
0.05 2.357 0 0.0 1e-06 
3.0 2.357 0 0.0 1e-06 
0.05 2.358 0 0.0 1e-06 
3.0 2.358 0 0.0 1e-06 
0.05 2.359 0 0.0 1e-06 
3.0 2.359 0 0.0 1e-06 
0.05 2.36 0 0.0 1e-06 
3.0 2.36 0 0.0 1e-06 
0.05 2.361 0 0.0 1e-06 
3.0 2.361 0 0.0 1e-06 
0.05 2.362 0 0.0 1e-06 
3.0 2.362 0 0.0 1e-06 
0.05 2.363 0 0.0 1e-06 
3.0 2.363 0 0.0 1e-06 
0.05 2.364 0 0.0 1e-06 
3.0 2.364 0 0.0 1e-06 
0.05 2.365 0 0.0 1e-06 
3.0 2.365 0 0.0 1e-06 
0.05 2.366 0 0.0 1e-06 
3.0 2.366 0 0.0 1e-06 
0.05 2.367 0 0.0 1e-06 
3.0 2.367 0 0.0 1e-06 
0.05 2.368 0 0.0 1e-06 
3.0 2.368 0 0.0 1e-06 
0.05 2.369 0 0.0 1e-06 
3.0 2.369 0 0.0 1e-06 
0.05 2.37 0 0.0 1e-06 
3.0 2.37 0 0.0 1e-06 
0.05 2.371 0 0.0 1e-06 
3.0 2.371 0 0.0 1e-06 
0.05 2.372 0 0.0 1e-06 
3.0 2.372 0 0.0 1e-06 
0.05 2.373 0 0.0 1e-06 
3.0 2.373 0 0.0 1e-06 
0.05 2.374 0 0.0 1e-06 
3.0 2.374 0 0.0 1e-06 
0.05 2.375 0 0.0 1e-06 
3.0 2.375 0 0.0 1e-06 
0.05 2.376 0 0.0 1e-06 
3.0 2.376 0 0.0 1e-06 
0.05 2.377 0 0.0 1e-06 
3.0 2.377 0 0.0 1e-06 
0.05 2.378 0 0.0 1e-06 
3.0 2.378 0 0.0 1e-06 
0.05 2.379 0 0.0 1e-06 
3.0 2.379 0 0.0 1e-06 
0.05 2.38 0 0.0 1e-06 
3.0 2.38 0 0.0 1e-06 
0.05 2.381 0 0.0 1e-06 
3.0 2.381 0 0.0 1e-06 
0.05 2.382 0 0.0 1e-06 
3.0 2.382 0 0.0 1e-06 
0.05 2.383 0 0.0 1e-06 
3.0 2.383 0 0.0 1e-06 
0.05 2.384 0 0.0 1e-06 
3.0 2.384 0 0.0 1e-06 
0.05 2.385 0 0.0 1e-06 
3.0 2.385 0 0.0 1e-06 
0.05 2.386 0 0.0 1e-06 
3.0 2.386 0 0.0 1e-06 
0.05 2.387 0 0.0 1e-06 
3.0 2.387 0 0.0 1e-06 
0.05 2.388 0 0.0 1e-06 
3.0 2.388 0 0.0 1e-06 
0.05 2.389 0 0.0 1e-06 
3.0 2.389 0 0.0 1e-06 
0.05 2.39 0 0.0 1e-06 
3.0 2.39 0 0.0 1e-06 
0.05 2.391 0 0.0 1e-06 
3.0 2.391 0 0.0 1e-06 
0.05 2.392 0 0.0 1e-06 
3.0 2.392 0 0.0 1e-06 
0.05 2.393 0 0.0 1e-06 
3.0 2.393 0 0.0 1e-06 
0.05 2.394 0 0.0 1e-06 
3.0 2.394 0 0.0 1e-06 
0.05 2.395 0 0.0 1e-06 
3.0 2.395 0 0.0 1e-06 
0.05 2.396 0 0.0 1e-06 
3.0 2.396 0 0.0 1e-06 
0.05 2.397 0 0.0 1e-06 
3.0 2.397 0 0.0 1e-06 
0.05 2.398 0 0.0 1e-06 
3.0 2.398 0 0.0 1e-06 
0.05 2.399 0 0.0 1e-06 
3.0 2.399 0 0.0 1e-06 
0.05 2.4 0 0.0 1e-06 
3.0 2.4 0 0.0 1e-06 
0.05 2.401 0 0.0 1e-06 
3.0 2.401 0 0.0 1e-06 
0.05 2.402 0 0.0 1e-06 
3.0 2.402 0 0.0 1e-06 
0.05 2.403 0 0.0 1e-06 
3.0 2.403 0 0.0 1e-06 
0.05 2.404 0 0.0 1e-06 
3.0 2.404 0 0.0 1e-06 
0.05 2.405 0 0.0 1e-06 
3.0 2.405 0 0.0 1e-06 
0.05 2.406 0 0.0 1e-06 
3.0 2.406 0 0.0 1e-06 
0.05 2.407 0 0.0 1e-06 
3.0 2.407 0 0.0 1e-06 
0.05 2.408 0 0.0 1e-06 
3.0 2.408 0 0.0 1e-06 
0.05 2.409 0 0.0 1e-06 
3.0 2.409 0 0.0 1e-06 
0.05 2.41 0 0.0 1e-06 
3.0 2.41 0 0.0 1e-06 
0.05 2.411 0 0.0 1e-06 
3.0 2.411 0 0.0 1e-06 
0.05 2.412 0 0.0 1e-06 
3.0 2.412 0 0.0 1e-06 
0.05 2.413 0 0.0 1e-06 
3.0 2.413 0 0.0 1e-06 
0.05 2.414 0 0.0 1e-06 
3.0 2.414 0 0.0 1e-06 
0.05 2.415 0 0.0 1e-06 
3.0 2.415 0 0.0 1e-06 
0.05 2.416 0 0.0 1e-06 
3.0 2.416 0 0.0 1e-06 
0.05 2.417 0 0.0 1e-06 
3.0 2.417 0 0.0 1e-06 
0.05 2.418 0 0.0 1e-06 
3.0 2.418 0 0.0 1e-06 
0.05 2.419 0 0.0 1e-06 
3.0 2.419 0 0.0 1e-06 
0.05 2.42 0 0.0 1e-06 
3.0 2.42 0 0.0 1e-06 
0.05 2.421 0 0.0 1e-06 
3.0 2.421 0 0.0 1e-06 
0.05 2.422 0 0.0 1e-06 
3.0 2.422 0 0.0 1e-06 
0.05 2.423 0 0.0 1e-06 
3.0 2.423 0 0.0 1e-06 
0.05 2.424 0 0.0 1e-06 
3.0 2.424 0 0.0 1e-06 
0.05 2.425 0 0.0 1e-06 
3.0 2.425 0 0.0 1e-06 
0.05 2.426 0 0.0 1e-06 
3.0 2.426 0 0.0 1e-06 
0.05 2.427 0 0.0 1e-06 
3.0 2.427 0 0.0 1e-06 
0.05 2.428 0 0.0 1e-06 
3.0 2.428 0 0.0 1e-06 
0.05 2.429 0 0.0 1e-06 
3.0 2.429 0 0.0 1e-06 
0.05 2.43 0 0.0 1e-06 
3.0 2.43 0 0.0 1e-06 
0.05 2.431 0 0.0 1e-06 
3.0 2.431 0 0.0 1e-06 
0.05 2.432 0 0.0 1e-06 
3.0 2.432 0 0.0 1e-06 
0.05 2.433 0 0.0 1e-06 
3.0 2.433 0 0.0 1e-06 
0.05 2.434 0 0.0 1e-06 
3.0 2.434 0 0.0 1e-06 
0.05 2.435 0 0.0 1e-06 
3.0 2.435 0 0.0 1e-06 
0.05 2.436 0 0.0 1e-06 
3.0 2.436 0 0.0 1e-06 
0.05 2.437 0 0.0 1e-06 
3.0 2.437 0 0.0 1e-06 
0.05 2.438 0 0.0 1e-06 
3.0 2.438 0 0.0 1e-06 
0.05 2.439 0 0.0 1e-06 
3.0 2.439 0 0.0 1e-06 
0.05 2.44 0 0.0 1e-06 
3.0 2.44 0 0.0 1e-06 
0.05 2.441 0 0.0 1e-06 
3.0 2.441 0 0.0 1e-06 
0.05 2.442 0 0.0 1e-06 
3.0 2.442 0 0.0 1e-06 
0.05 2.443 0 0.0 1e-06 
3.0 2.443 0 0.0 1e-06 
0.05 2.444 0 0.0 1e-06 
3.0 2.444 0 0.0 1e-06 
0.05 2.445 0 0.0 1e-06 
3.0 2.445 0 0.0 1e-06 
0.05 2.446 0 0.0 1e-06 
3.0 2.446 0 0.0 1e-06 
0.05 2.447 0 0.0 1e-06 
3.0 2.447 0 0.0 1e-06 
0.05 2.448 0 0.0 1e-06 
3.0 2.448 0 0.0 1e-06 
0.05 2.449 0 0.0 1e-06 
3.0 2.449 0 0.0 1e-06 
0.05 2.45 0 0.0 1e-06 
3.0 2.45 0 0.0 1e-06 
0.05 2.451 0 0.0 1e-06 
3.0 2.451 0 0.0 1e-06 
0.05 2.452 0 0.0 1e-06 
3.0 2.452 0 0.0 1e-06 
0.05 2.453 0 0.0 1e-06 
3.0 2.453 0 0.0 1e-06 
0.05 2.454 0 0.0 1e-06 
3.0 2.454 0 0.0 1e-06 
0.05 2.455 0 0.0 1e-06 
3.0 2.455 0 0.0 1e-06 
0.05 2.456 0 0.0 1e-06 
3.0 2.456 0 0.0 1e-06 
0.05 2.457 0 0.0 1e-06 
3.0 2.457 0 0.0 1e-06 
0.05 2.458 0 0.0 1e-06 
3.0 2.458 0 0.0 1e-06 
0.05 2.459 0 0.0 1e-06 
3.0 2.459 0 0.0 1e-06 
0.05 2.46 0 0.0 1e-06 
3.0 2.46 0 0.0 1e-06 
0.05 2.461 0 0.0 1e-06 
3.0 2.461 0 0.0 1e-06 
0.05 2.462 0 0.0 1e-06 
3.0 2.462 0 0.0 1e-06 
0.05 2.463 0 0.0 1e-06 
3.0 2.463 0 0.0 1e-06 
0.05 2.464 0 0.0 1e-06 
3.0 2.464 0 0.0 1e-06 
0.05 2.465 0 0.0 1e-06 
3.0 2.465 0 0.0 1e-06 
0.05 2.466 0 0.0 1e-06 
3.0 2.466 0 0.0 1e-06 
0.05 2.467 0 0.0 1e-06 
3.0 2.467 0 0.0 1e-06 
0.05 2.468 0 0.0 1e-06 
3.0 2.468 0 0.0 1e-06 
0.05 2.469 0 0.0 1e-06 
3.0 2.469 0 0.0 1e-06 
0.05 2.47 0 0.0 1e-06 
3.0 2.47 0 0.0 1e-06 
0.05 2.471 0 0.0 1e-06 
3.0 2.471 0 0.0 1e-06 
0.05 2.472 0 0.0 1e-06 
3.0 2.472 0 0.0 1e-06 
0.05 2.473 0 0.0 1e-06 
3.0 2.473 0 0.0 1e-06 
0.05 2.474 0 0.0 1e-06 
3.0 2.474 0 0.0 1e-06 
0.05 2.475 0 0.0 1e-06 
3.0 2.475 0 0.0 1e-06 
0.05 2.476 0 0.0 1e-06 
3.0 2.476 0 0.0 1e-06 
0.05 2.477 0 0.0 1e-06 
3.0 2.477 0 0.0 1e-06 
0.05 2.478 0 0.0 1e-06 
3.0 2.478 0 0.0 1e-06 
0.05 2.479 0 0.0 1e-06 
3.0 2.479 0 0.0 1e-06 
0.05 2.48 0 0.0 1e-06 
3.0 2.48 0 0.0 1e-06 
0.05 2.481 0 0.0 1e-06 
3.0 2.481 0 0.0 1e-06 
0.05 2.482 0 0.0 1e-06 
3.0 2.482 0 0.0 1e-06 
0.05 2.483 0 0.0 1e-06 
3.0 2.483 0 0.0 1e-06 
0.05 2.484 0 0.0 1e-06 
3.0 2.484 0 0.0 1e-06 
0.05 2.485 0 0.0 1e-06 
3.0 2.485 0 0.0 1e-06 
0.05 2.486 0 0.0 1e-06 
3.0 2.486 0 0.0 1e-06 
0.05 2.487 0 0.0 1e-06 
3.0 2.487 0 0.0 1e-06 
0.05 2.488 0 0.0 1e-06 
3.0 2.488 0 0.0 1e-06 
0.05 2.489 0 0.0 1e-06 
3.0 2.489 0 0.0 1e-06 
0.05 2.49 0 0.0 1e-06 
3.0 2.49 0 0.0 1e-06 
0.05 2.491 0 0.0 1e-06 
3.0 2.491 0 0.0 1e-06 
0.05 2.492 0 0.0 1e-06 
3.0 2.492 0 0.0 1e-06 
0.05 2.493 0 0.0 1e-06 
3.0 2.493 0 0.0 1e-06 
0.05 2.494 0 0.0 1e-06 
3.0 2.494 0 0.0 1e-06 
0.05 2.495 0 0.0 1e-06 
3.0 2.495 0 0.0 1e-06 
0.05 2.496 0 0.0 1e-06 
3.0 2.496 0 0.0 1e-06 
0.05 2.497 0 0.0 1e-06 
3.0 2.497 0 0.0 1e-06 
0.05 2.498 0 0.0 1e-06 
3.0 2.498 0 0.0 1e-06 
0.05 2.499 0 0.0 1e-06 
3.0 2.499 0 0.0 1e-06 
0.05 2.5 0 0.0 1e-06 
3.0 2.5 0 0.0 1e-06 
0.05 2.501 0 0.0 1e-06 
3.0 2.501 0 0.0 1e-06 
0.05 2.502 0 0.0 1e-06 
3.0 2.502 0 0.0 1e-06 
0.05 2.503 0 0.0 1e-06 
3.0 2.503 0 0.0 1e-06 
0.05 2.504 0 0.0 1e-06 
3.0 2.504 0 0.0 1e-06 
0.05 2.505 0 0.0 1e-06 
3.0 2.505 0 0.0 1e-06 
0.05 2.506 0 0.0 1e-06 
3.0 2.506 0 0.0 1e-06 
0.05 2.507 0 0.0 1e-06 
3.0 2.507 0 0.0 1e-06 
0.05 2.508 0 0.0 1e-06 
3.0 2.508 0 0.0 1e-06 
0.05 2.509 0 0.0 1e-06 
3.0 2.509 0 0.0 1e-06 
0.05 2.51 0 0.0 1e-06 
3.0 2.51 0 0.0 1e-06 
0.05 2.511 0 0.0 1e-06 
3.0 2.511 0 0.0 1e-06 
0.05 2.512 0 0.0 1e-06 
3.0 2.512 0 0.0 1e-06 
0.05 2.513 0 0.0 1e-06 
3.0 2.513 0 0.0 1e-06 
0.05 2.514 0 0.0 1e-06 
3.0 2.514 0 0.0 1e-06 
0.05 2.515 0 0.0 1e-06 
3.0 2.515 0 0.0 1e-06 
0.05 2.516 0 0.0 1e-06 
3.0 2.516 0 0.0 1e-06 
0.05 2.517 0 0.0 1e-06 
3.0 2.517 0 0.0 1e-06 
0.05 2.518 0 0.0 1e-06 
3.0 2.518 0 0.0 1e-06 
0.05 2.519 0 0.0 1e-06 
3.0 2.519 0 0.0 1e-06 
0.05 2.52 0 0.0 1e-06 
3.0 2.52 0 0.0 1e-06 
0.05 2.521 0 0.0 1e-06 
3.0 2.521 0 0.0 1e-06 
0.05 2.522 0 0.0 1e-06 
3.0 2.522 0 0.0 1e-06 
0.05 2.523 0 0.0 1e-06 
3.0 2.523 0 0.0 1e-06 
0.05 2.524 0 0.0 1e-06 
3.0 2.524 0 0.0 1e-06 
0.05 2.525 0 0.0 1e-06 
3.0 2.525 0 0.0 1e-06 
0.05 2.526 0 0.0 1e-06 
3.0 2.526 0 0.0 1e-06 
0.05 2.527 0 0.0 1e-06 
3.0 2.527 0 0.0 1e-06 
0.05 2.528 0 0.0 1e-06 
3.0 2.528 0 0.0 1e-06 
0.05 2.529 0 0.0 1e-06 
3.0 2.529 0 0.0 1e-06 
0.05 2.53 0 0.0 1e-06 
3.0 2.53 0 0.0 1e-06 
0.05 2.531 0 0.0 1e-06 
3.0 2.531 0 0.0 1e-06 
0.05 2.532 0 0.0 1e-06 
3.0 2.532 0 0.0 1e-06 
0.05 2.533 0 0.0 1e-06 
3.0 2.533 0 0.0 1e-06 
0.05 2.534 0 0.0 1e-06 
3.0 2.534 0 0.0 1e-06 
0.05 2.535 0 0.0 1e-06 
3.0 2.535 0 0.0 1e-06 
0.05 2.536 0 0.0 1e-06 
3.0 2.536 0 0.0 1e-06 
0.05 2.537 0 0.0 1e-06 
3.0 2.537 0 0.0 1e-06 
0.05 2.538 0 0.0 1e-06 
3.0 2.538 0 0.0 1e-06 
0.05 2.539 0 0.0 1e-06 
3.0 2.539 0 0.0 1e-06 
0.05 2.54 0 0.0 1e-06 
3.0 2.54 0 0.0 1e-06 
0.05 2.541 0 0.0 1e-06 
3.0 2.541 0 0.0 1e-06 
0.05 2.542 0 0.0 1e-06 
3.0 2.542 0 0.0 1e-06 
0.05 2.543 0 0.0 1e-06 
3.0 2.543 0 0.0 1e-06 
0.05 2.544 0 0.0 1e-06 
3.0 2.544 0 0.0 1e-06 
0.05 2.545 0 0.0 1e-06 
3.0 2.545 0 0.0 1e-06 
0.05 2.546 0 0.0 1e-06 
3.0 2.546 0 0.0 1e-06 
0.05 2.547 0 0.0 1e-06 
3.0 2.547 0 0.0 1e-06 
0.05 2.548 0 0.0 1e-06 
3.0 2.548 0 0.0 1e-06 
0.05 2.549 0 0.0 1e-06 
3.0 2.549 0 0.0 1e-06 
0.05 2.55 0 0.0 1e-06 
3.0 2.55 0 0.0 1e-06 
0.05 2.551 0 0.0 1e-06 
3.0 2.551 0 0.0 1e-06 
0.05 2.552 0 0.0 1e-06 
3.0 2.552 0 0.0 1e-06 
0.05 2.553 0 0.0 1e-06 
3.0 2.553 0 0.0 1e-06 
0.05 2.554 0 0.0 1e-06 
3.0 2.554 0 0.0 1e-06 
0.05 2.555 0 0.0 1e-06 
3.0 2.555 0 0.0 1e-06 
0.05 2.556 0 0.0 1e-06 
3.0 2.556 0 0.0 1e-06 
0.05 2.557 0 0.0 1e-06 
3.0 2.557 0 0.0 1e-06 
0.05 2.558 0 0.0 1e-06 
3.0 2.558 0 0.0 1e-06 
0.05 2.559 0 0.0 1e-06 
3.0 2.559 0 0.0 1e-06 
0.05 2.56 0 0.0 1e-06 
3.0 2.56 0 0.0 1e-06 
0.05 2.561 0 0.0 1e-06 
3.0 2.561 0 0.0 1e-06 
0.05 2.562 0 0.0 1e-06 
3.0 2.562 0 0.0 1e-06 
0.05 2.563 0 0.0 1e-06 
3.0 2.563 0 0.0 1e-06 
0.05 2.564 0 0.0 1e-06 
3.0 2.564 0 0.0 1e-06 
0.05 2.565 0 0.0 1e-06 
3.0 2.565 0 0.0 1e-06 
0.05 2.566 0 0.0 1e-06 
3.0 2.566 0 0.0 1e-06 
0.05 2.567 0 0.0 1e-06 
3.0 2.567 0 0.0 1e-06 
0.05 2.568 0 0.0 1e-06 
3.0 2.568 0 0.0 1e-06 
0.05 2.569 0 0.0 1e-06 
3.0 2.569 0 0.0 1e-06 
0.05 2.57 0 0.0 1e-06 
3.0 2.57 0 0.0 1e-06 
0.05 2.571 0 0.0 1e-06 
3.0 2.571 0 0.0 1e-06 
0.05 2.572 0 0.0 1e-06 
3.0 2.572 0 0.0 1e-06 
0.05 2.573 0 0.0 1e-06 
3.0 2.573 0 0.0 1e-06 
0.05 2.574 0 0.0 1e-06 
3.0 2.574 0 0.0 1e-06 
0.05 2.575 0 0.0 1e-06 
3.0 2.575 0 0.0 1e-06 
0.05 2.576 0 0.0 1e-06 
3.0 2.576 0 0.0 1e-06 
0.05 2.577 0 0.0 1e-06 
3.0 2.577 0 0.0 1e-06 
0.05 2.578 0 0.0 1e-06 
3.0 2.578 0 0.0 1e-06 
0.05 2.579 0 0.0 1e-06 
3.0 2.579 0 0.0 1e-06 
0.05 2.58 0 0.0 1e-06 
3.0 2.58 0 0.0 1e-06 
0.05 2.581 0 0.0 1e-06 
3.0 2.581 0 0.0 1e-06 
0.05 2.582 0 0.0 1e-06 
3.0 2.582 0 0.0 1e-06 
0.05 2.583 0 0.0 1e-06 
3.0 2.583 0 0.0 1e-06 
0.05 2.584 0 0.0 1e-06 
3.0 2.584 0 0.0 1e-06 
0.05 2.585 0 0.0 1e-06 
3.0 2.585 0 0.0 1e-06 
0.05 2.586 0 0.0 1e-06 
3.0 2.586 0 0.0 1e-06 
0.05 2.587 0 0.0 1e-06 
3.0 2.587 0 0.0 1e-06 
0.05 2.588 0 0.0 1e-06 
3.0 2.588 0 0.0 1e-06 
0.05 2.589 0 0.0 1e-06 
3.0 2.589 0 0.0 1e-06 
0.05 2.59 0 0.0 1e-06 
3.0 2.59 0 0.0 1e-06 
0.05 2.591 0 0.0 1e-06 
3.0 2.591 0 0.0 1e-06 
0.05 2.592 0 0.0 1e-06 
3.0 2.592 0 0.0 1e-06 
0.05 2.593 0 0.0 1e-06 
3.0 2.593 0 0.0 1e-06 
0.05 2.594 0 0.0 1e-06 
3.0 2.594 0 0.0 1e-06 
0.05 2.595 0 0.0 1e-06 
3.0 2.595 0 0.0 1e-06 
0.05 2.596 0 0.0 1e-06 
3.0 2.596 0 0.0 1e-06 
0.05 2.597 0 0.0 1e-06 
3.0 2.597 0 0.0 1e-06 
0.05 2.598 0 0.0 1e-06 
3.0 2.598 0 0.0 1e-06 
0.05 2.599 0 0.0 1e-06 
3.0 2.599 0 0.0 1e-06 
0.05 2.6 0 0.0 1e-06 
3.0 2.6 0 0.0 1e-06 
0.05 2.601 0 0.0 1e-06 
3.0 2.601 0 0.0 1e-06 
0.05 2.602 0 0.0 1e-06 
3.0 2.602 0 0.0 1e-06 
0.05 2.603 0 0.0 1e-06 
3.0 2.603 0 0.0 1e-06 
0.05 2.604 0 0.0 1e-06 
3.0 2.604 0 0.0 1e-06 
0.05 2.605 0 0.0 1e-06 
3.0 2.605 0 0.0 1e-06 
0.05 2.606 0 0.0 1e-06 
3.0 2.606 0 0.0 1e-06 
0.05 2.607 0 0.0 1e-06 
3.0 2.607 0 0.0 1e-06 
0.05 2.608 0 0.0 1e-06 
3.0 2.608 0 0.0 1e-06 
0.05 2.609 0 0.0 1e-06 
3.0 2.609 0 0.0 1e-06 
0.05 2.61 0 0.0 1e-06 
3.0 2.61 0 0.0 1e-06 
0.05 2.611 0 0.0 1e-06 
3.0 2.611 0 0.0 1e-06 
0.05 2.612 0 0.0 1e-06 
3.0 2.612 0 0.0 1e-06 
0.05 2.613 0 0.0 1e-06 
3.0 2.613 0 0.0 1e-06 
0.05 2.614 0 0.0 1e-06 
3.0 2.614 0 0.0 1e-06 
0.05 2.615 0 0.0 1e-06 
3.0 2.615 0 0.0 1e-06 
0.05 2.616 0 0.0 1e-06 
3.0 2.616 0 0.0 1e-06 
0.05 2.617 0 0.0 1e-06 
3.0 2.617 0 0.0 1e-06 
0.05 2.618 0 0.0 1e-06 
3.0 2.618 0 0.0 1e-06 
0.05 2.619 0 0.0 1e-06 
3.0 2.619 0 0.0 1e-06 
0.05 2.62 0 0.0 1e-06 
3.0 2.62 0 0.0 1e-06 
0.05 2.621 0 0.0 1e-06 
3.0 2.621 0 0.0 1e-06 
0.05 2.622 0 0.0 1e-06 
3.0 2.622 0 0.0 1e-06 
0.05 2.623 0 0.0 1e-06 
3.0 2.623 0 0.0 1e-06 
0.05 2.624 0 0.0 1e-06 
3.0 2.624 0 0.0 1e-06 
0.05 2.625 0 0.0 1e-06 
3.0 2.625 0 0.0 1e-06 
0.05 2.626 0 0.0 1e-06 
3.0 2.626 0 0.0 1e-06 
0.05 2.627 0 0.0 1e-06 
3.0 2.627 0 0.0 1e-06 
0.05 2.628 0 0.0 1e-06 
3.0 2.628 0 0.0 1e-06 
0.05 2.629 0 0.0 1e-06 
3.0 2.629 0 0.0 1e-06 
0.05 2.63 0 0.0 1e-06 
3.0 2.63 0 0.0 1e-06 
0.05 2.631 0 0.0 1e-06 
3.0 2.631 0 0.0 1e-06 
0.05 2.632 0 0.0 1e-06 
3.0 2.632 0 0.0 1e-06 
0.05 2.633 0 0.0 1e-06 
3.0 2.633 0 0.0 1e-06 
0.05 2.634 0 0.0 1e-06 
3.0 2.634 0 0.0 1e-06 
0.05 2.635 0 0.0 1e-06 
3.0 2.635 0 0.0 1e-06 
0.05 2.636 0 0.0 1e-06 
3.0 2.636 0 0.0 1e-06 
0.05 2.637 0 0.0 1e-06 
3.0 2.637 0 0.0 1e-06 
0.05 2.638 0 0.0 1e-06 
3.0 2.638 0 0.0 1e-06 
0.05 2.639 0 0.0 1e-06 
3.0 2.639 0 0.0 1e-06 
0.05 2.64 0 0.0 1e-06 
3.0 2.64 0 0.0 1e-06 
0.05 2.641 0 0.0 1e-06 
3.0 2.641 0 0.0 1e-06 
0.05 2.642 0 0.0 1e-06 
3.0 2.642 0 0.0 1e-06 
0.05 2.643 0 0.0 1e-06 
3.0 2.643 0 0.0 1e-06 
0.05 2.644 0 0.0 1e-06 
3.0 2.644 0 0.0 1e-06 
0.05 2.645 0 0.0 1e-06 
3.0 2.645 0 0.0 1e-06 
0.05 2.646 0 0.0 1e-06 
3.0 2.646 0 0.0 1e-06 
0.05 2.647 0 0.0 1e-06 
3.0 2.647 0 0.0 1e-06 
0.05 2.648 0 0.0 1e-06 
3.0 2.648 0 0.0 1e-06 
0.05 2.649 0 0.0 1e-06 
3.0 2.649 0 0.0 1e-06 
0.05 2.65 0 0.0 1e-06 
3.0 2.65 0 0.0 1e-06 
0.05 2.651 0 0.0 1e-06 
3.0 2.651 0 0.0 1e-06 
0.05 2.652 0 0.0 1e-06 
3.0 2.652 0 0.0 1e-06 
0.05 2.653 0 0.0 1e-06 
3.0 2.653 0 0.0 1e-06 
0.05 2.654 0 0.0 1e-06 
3.0 2.654 0 0.0 1e-06 
0.05 2.655 0 0.0 1e-06 
3.0 2.655 0 0.0 1e-06 
0.05 2.656 0 0.0 1e-06 
3.0 2.656 0 0.0 1e-06 
0.05 2.657 0 0.0 1e-06 
3.0 2.657 0 0.0 1e-06 
0.05 2.658 0 0.0 1e-06 
3.0 2.658 0 0.0 1e-06 
0.05 2.659 0 0.0 1e-06 
3.0 2.659 0 0.0 1e-06 
0.05 2.66 0 0.0 1e-06 
3.0 2.66 0 0.0 1e-06 
0.05 2.661 0 0.0 1e-06 
3.0 2.661 0 0.0 1e-06 
0.05 2.662 0 0.0 1e-06 
3.0 2.662 0 0.0 1e-06 
0.05 2.663 0 0.0 1e-06 
3.0 2.663 0 0.0 1e-06 
0.05 2.664 0 0.0 1e-06 
3.0 2.664 0 0.0 1e-06 
0.05 2.665 0 0.0 1e-06 
3.0 2.665 0 0.0 1e-06 
0.05 2.666 0 0.0 1e-06 
3.0 2.666 0 0.0 1e-06 
0.05 2.667 0 0.0 1e-06 
3.0 2.667 0 0.0 1e-06 
0.05 2.668 0 0.0 1e-06 
3.0 2.668 0 0.0 1e-06 
0.05 2.669 0 0.0 1e-06 
3.0 2.669 0 0.0 1e-06 
0.05 2.67 0 0.0 1e-06 
3.0 2.67 0 0.0 1e-06 
0.05 2.671 0 0.0 1e-06 
3.0 2.671 0 0.0 1e-06 
0.05 2.672 0 0.0 1e-06 
3.0 2.672 0 0.0 1e-06 
0.05 2.673 0 0.0 1e-06 
3.0 2.673 0 0.0 1e-06 
0.05 2.674 0 0.0 1e-06 
3.0 2.674 0 0.0 1e-06 
0.05 2.675 0 0.0 1e-06 
3.0 2.675 0 0.0 1e-06 
0.05 2.676 0 0.0 1e-06 
3.0 2.676 0 0.0 1e-06 
0.05 2.677 0 0.0 1e-06 
3.0 2.677 0 0.0 1e-06 
0.05 2.678 0 0.0 1e-06 
3.0 2.678 0 0.0 1e-06 
0.05 2.679 0 0.0 1e-06 
3.0 2.679 0 0.0 1e-06 
0.05 2.68 0 0.0 1e-06 
3.0 2.68 0 0.0 1e-06 
0.05 2.681 0 0.0 1e-06 
3.0 2.681 0 0.0 1e-06 
0.05 2.682 0 0.0 1e-06 
3.0 2.682 0 0.0 1e-06 
0.05 2.683 0 0.0 1e-06 
3.0 2.683 0 0.0 1e-06 
0.05 2.684 0 0.0 1e-06 
3.0 2.684 0 0.0 1e-06 
0.05 2.685 0 0.0 1e-06 
3.0 2.685 0 0.0 1e-06 
0.05 2.686 0 0.0 1e-06 
3.0 2.686 0 0.0 1e-06 
0.05 2.687 0 0.0 1e-06 
3.0 2.687 0 0.0 1e-06 
0.05 2.688 0 0.0 1e-06 
3.0 2.688 0 0.0 1e-06 
0.05 2.689 0 0.0 1e-06 
3.0 2.689 0 0.0 1e-06 
0.05 2.69 0 0.0 1e-06 
3.0 2.69 0 0.0 1e-06 
0.05 2.691 0 0.0 1e-06 
3.0 2.691 0 0.0 1e-06 
0.05 2.692 0 0.0 1e-06 
3.0 2.692 0 0.0 1e-06 
0.05 2.693 0 0.0 1e-06 
3.0 2.693 0 0.0 1e-06 
0.05 2.694 0 0.0 1e-06 
3.0 2.694 0 0.0 1e-06 
0.05 2.695 0 0.0 1e-06 
3.0 2.695 0 0.0 1e-06 
0.05 2.696 0 0.0 1e-06 
3.0 2.696 0 0.0 1e-06 
0.05 2.697 0 0.0 1e-06 
3.0 2.697 0 0.0 1e-06 
0.05 2.698 0 0.0 1e-06 
3.0 2.698 0 0.0 1e-06 
0.05 2.699 0 0.0 1e-06 
3.0 2.699 0 0.0 1e-06 
0.05 2.7 0 0.0 1e-06 
3.0 2.7 0 0.0 1e-06 
0.05 2.701 0 0.0 1e-06 
3.0 2.701 0 0.0 1e-06 
0.05 2.702 0 0.0 1e-06 
3.0 2.702 0 0.0 1e-06 
0.05 2.703 0 0.0 1e-06 
3.0 2.703 0 0.0 1e-06 
0.05 2.704 0 0.0 1e-06 
3.0 2.704 0 0.0 1e-06 
0.05 2.705 0 0.0 1e-06 
3.0 2.705 0 0.0 1e-06 
0.05 2.706 0 0.0 1e-06 
3.0 2.706 0 0.0 1e-06 
0.05 2.707 0 0.0 1e-06 
3.0 2.707 0 0.0 1e-06 
0.05 2.708 0 0.0 1e-06 
3.0 2.708 0 0.0 1e-06 
0.05 2.709 0 0.0 1e-06 
3.0 2.709 0 0.0 1e-06 
0.05 2.71 0 0.0 1e-06 
3.0 2.71 0 0.0 1e-06 
0.05 2.711 0 0.0 1e-06 
3.0 2.711 0 0.0 1e-06 
0.05 2.712 0 0.0 1e-06 
3.0 2.712 0 0.0 1e-06 
0.05 2.713 0 0.0 1e-06 
3.0 2.713 0 0.0 1e-06 
0.05 2.714 0 0.0 1e-06 
3.0 2.714 0 0.0 1e-06 
0.05 2.715 0 0.0 1e-06 
3.0 2.715 0 0.0 1e-06 
0.05 2.716 0 0.0 1e-06 
3.0 2.716 0 0.0 1e-06 
0.05 2.717 0 0.0 1e-06 
3.0 2.717 0 0.0 1e-06 
0.05 2.718 0 0.0 1e-06 
3.0 2.718 0 0.0 1e-06 
0.05 2.719 0 0.0 1e-06 
3.0 2.719 0 0.0 1e-06 
0.05 2.72 0 0.0 1e-06 
3.0 2.72 0 0.0 1e-06 
0.05 2.721 0 0.0 1e-06 
3.0 2.721 0 0.0 1e-06 
0.05 2.722 0 0.0 1e-06 
3.0 2.722 0 0.0 1e-06 
0.05 2.723 0 0.0 1e-06 
3.0 2.723 0 0.0 1e-06 
0.05 2.724 0 0.0 1e-06 
3.0 2.724 0 0.0 1e-06 
0.05 2.725 0 0.0 1e-06 
3.0 2.725 0 0.0 1e-06 
0.05 2.726 0 0.0 1e-06 
3.0 2.726 0 0.0 1e-06 
0.05 2.727 0 0.0 1e-06 
3.0 2.727 0 0.0 1e-06 
0.05 2.728 0 0.0 1e-06 
3.0 2.728 0 0.0 1e-06 
0.05 2.729 0 0.0 1e-06 
3.0 2.729 0 0.0 1e-06 
0.05 2.73 0 0.0 1e-06 
3.0 2.73 0 0.0 1e-06 
0.05 2.731 0 0.0 1e-06 
3.0 2.731 0 0.0 1e-06 
0.05 2.732 0 0.0 1e-06 
3.0 2.732 0 0.0 1e-06 
0.05 2.733 0 0.0 1e-06 
3.0 2.733 0 0.0 1e-06 
0.05 2.734 0 0.0 1e-06 
3.0 2.734 0 0.0 1e-06 
0.05 2.735 0 0.0 1e-06 
3.0 2.735 0 0.0 1e-06 
0.05 2.736 0 0.0 1e-06 
3.0 2.736 0 0.0 1e-06 
0.05 2.737 0 0.0 1e-06 
3.0 2.737 0 0.0 1e-06 
0.05 2.738 0 0.0 1e-06 
3.0 2.738 0 0.0 1e-06 
0.05 2.739 0 0.0 1e-06 
3.0 2.739 0 0.0 1e-06 
0.05 2.74 0 0.0 1e-06 
3.0 2.74 0 0.0 1e-06 
0.05 2.741 0 0.0 1e-06 
3.0 2.741 0 0.0 1e-06 
0.05 2.742 0 0.0 1e-06 
3.0 2.742 0 0.0 1e-06 
0.05 2.743 0 0.0 1e-06 
3.0 2.743 0 0.0 1e-06 
0.05 2.744 0 0.0 1e-06 
3.0 2.744 0 0.0 1e-06 
0.05 2.745 0 0.0 1e-06 
3.0 2.745 0 0.0 1e-06 
0.05 2.746 0 0.0 1e-06 
3.0 2.746 0 0.0 1e-06 
0.05 2.747 0 0.0 1e-06 
3.0 2.747 0 0.0 1e-06 
0.05 2.748 0 0.0 1e-06 
3.0 2.748 0 0.0 1e-06 
0.05 2.749 0 0.0 1e-06 
3.0 2.749 0 0.0 1e-06 
0.05 2.75 0 0.0 1e-06 
3.0 2.75 0 0.0 1e-06 
0.05 2.751 0 0.0 1e-06 
3.0 2.751 0 0.0 1e-06 
0.05 2.752 0 0.0 1e-06 
3.0 2.752 0 0.0 1e-06 
0.05 2.753 0 0.0 1e-06 
3.0 2.753 0 0.0 1e-06 
0.05 2.754 0 0.0 1e-06 
3.0 2.754 0 0.0 1e-06 
0.05 2.755 0 0.0 1e-06 
3.0 2.755 0 0.0 1e-06 
0.05 2.756 0 0.0 1e-06 
3.0 2.756 0 0.0 1e-06 
0.05 2.757 0 0.0 1e-06 
3.0 2.757 0 0.0 1e-06 
0.05 2.758 0 0.0 1e-06 
3.0 2.758 0 0.0 1e-06 
0.05 2.759 0 0.0 1e-06 
3.0 2.759 0 0.0 1e-06 
0.05 2.76 0 0.0 1e-06 
3.0 2.76 0 0.0 1e-06 
0.05 2.761 0 0.0 1e-06 
3.0 2.761 0 0.0 1e-06 
0.05 2.762 0 0.0 1e-06 
3.0 2.762 0 0.0 1e-06 
0.05 2.763 0 0.0 1e-06 
3.0 2.763 0 0.0 1e-06 
0.05 2.764 0 0.0 1e-06 
3.0 2.764 0 0.0 1e-06 
0.05 2.765 0 0.0 1e-06 
3.0 2.765 0 0.0 1e-06 
0.05 2.766 0 0.0 1e-06 
3.0 2.766 0 0.0 1e-06 
0.05 2.767 0 0.0 1e-06 
3.0 2.767 0 0.0 1e-06 
0.05 2.768 0 0.0 1e-06 
3.0 2.768 0 0.0 1e-06 
0.05 2.769 0 0.0 1e-06 
3.0 2.769 0 0.0 1e-06 
0.05 2.77 0 0.0 1e-06 
3.0 2.77 0 0.0 1e-06 
0.05 2.771 0 0.0 1e-06 
3.0 2.771 0 0.0 1e-06 
0.05 2.772 0 0.0 1e-06 
3.0 2.772 0 0.0 1e-06 
0.05 2.773 0 0.0 1e-06 
3.0 2.773 0 0.0 1e-06 
0.05 2.774 0 0.0 1e-06 
3.0 2.774 0 0.0 1e-06 
0.05 2.775 0 0.0 1e-06 
3.0 2.775 0 0.0 1e-06 
0.05 2.776 0 0.0 1e-06 
3.0 2.776 0 0.0 1e-06 
0.05 2.777 0 0.0 1e-06 
3.0 2.777 0 0.0 1e-06 
0.05 2.778 0 0.0 1e-06 
3.0 2.778 0 0.0 1e-06 
0.05 2.779 0 0.0 1e-06 
3.0 2.779 0 0.0 1e-06 
0.05 2.78 0 0.0 1e-06 
3.0 2.78 0 0.0 1e-06 
0.05 2.781 0 0.0 1e-06 
3.0 2.781 0 0.0 1e-06 
0.05 2.782 0 0.0 1e-06 
3.0 2.782 0 0.0 1e-06 
0.05 2.783 0 0.0 1e-06 
3.0 2.783 0 0.0 1e-06 
0.05 2.784 0 0.0 1e-06 
3.0 2.784 0 0.0 1e-06 
0.05 2.785 0 0.0 1e-06 
3.0 2.785 0 0.0 1e-06 
0.05 2.786 0 0.0 1e-06 
3.0 2.786 0 0.0 1e-06 
0.05 2.787 0 0.0 1e-06 
3.0 2.787 0 0.0 1e-06 
0.05 2.788 0 0.0 1e-06 
3.0 2.788 0 0.0 1e-06 
0.05 2.789 0 0.0 1e-06 
3.0 2.789 0 0.0 1e-06 
0.05 2.79 0 0.0 1e-06 
3.0 2.79 0 0.0 1e-06 
0.05 2.791 0 0.0 1e-06 
3.0 2.791 0 0.0 1e-06 
0.05 2.792 0 0.0 1e-06 
3.0 2.792 0 0.0 1e-06 
0.05 2.793 0 0.0 1e-06 
3.0 2.793 0 0.0 1e-06 
0.05 2.794 0 0.0 1e-06 
3.0 2.794 0 0.0 1e-06 
0.05 2.795 0 0.0 1e-06 
3.0 2.795 0 0.0 1e-06 
0.05 2.796 0 0.0 1e-06 
3.0 2.796 0 0.0 1e-06 
0.05 2.797 0 0.0 1e-06 
3.0 2.797 0 0.0 1e-06 
0.05 2.798 0 0.0 1e-06 
3.0 2.798 0 0.0 1e-06 
0.05 2.799 0 0.0 1e-06 
3.0 2.799 0 0.0 1e-06 
0.05 2.8 0 0.0 1e-06 
3.0 2.8 0 0.0 1e-06 
0.05 2.801 0 0.0 1e-06 
3.0 2.801 0 0.0 1e-06 
0.05 2.802 0 0.0 1e-06 
3.0 2.802 0 0.0 1e-06 
0.05 2.803 0 0.0 1e-06 
3.0 2.803 0 0.0 1e-06 
0.05 2.804 0 0.0 1e-06 
3.0 2.804 0 0.0 1e-06 
0.05 2.805 0 0.0 1e-06 
3.0 2.805 0 0.0 1e-06 
0.05 2.806 0 0.0 1e-06 
3.0 2.806 0 0.0 1e-06 
0.05 2.807 0 0.0 1e-06 
3.0 2.807 0 0.0 1e-06 
0.05 2.808 0 0.0 1e-06 
3.0 2.808 0 0.0 1e-06 
0.05 2.809 0 0.0 1e-06 
3.0 2.809 0 0.0 1e-06 
0.05 2.81 0 0.0 1e-06 
3.0 2.81 0 0.0 1e-06 
0.05 2.811 0 0.0 1e-06 
3.0 2.811 0 0.0 1e-06 
0.05 2.812 0 0.0 1e-06 
3.0 2.812 0 0.0 1e-06 
0.05 2.813 0 0.0 1e-06 
3.0 2.813 0 0.0 1e-06 
0.05 2.814 0 0.0 1e-06 
3.0 2.814 0 0.0 1e-06 
0.05 2.815 0 0.0 1e-06 
3.0 2.815 0 0.0 1e-06 
0.05 2.816 0 0.0 1e-06 
3.0 2.816 0 0.0 1e-06 
0.05 2.817 0 0.0 1e-06 
3.0 2.817 0 0.0 1e-06 
0.05 2.818 0 0.0 1e-06 
3.0 2.818 0 0.0 1e-06 
0.05 2.819 0 0.0 1e-06 
3.0 2.819 0 0.0 1e-06 
0.05 2.82 0 0.0 1e-06 
3.0 2.82 0 0.0 1e-06 
0.05 2.821 0 0.0 1e-06 
3.0 2.821 0 0.0 1e-06 
0.05 2.822 0 0.0 1e-06 
3.0 2.822 0 0.0 1e-06 
0.05 2.823 0 0.0 1e-06 
3.0 2.823 0 0.0 1e-06 
0.05 2.824 0 0.0 1e-06 
3.0 2.824 0 0.0 1e-06 
0.05 2.825 0 0.0 1e-06 
3.0 2.825 0 0.0 1e-06 
0.05 2.826 0 0.0 1e-06 
3.0 2.826 0 0.0 1e-06 
0.05 2.827 0 0.0 1e-06 
3.0 2.827 0 0.0 1e-06 
0.05 2.828 0 0.0 1e-06 
3.0 2.828 0 0.0 1e-06 
0.05 2.829 0 0.0 1e-06 
3.0 2.829 0 0.0 1e-06 
0.05 2.83 0 0.0 1e-06 
3.0 2.83 0 0.0 1e-06 
0.05 2.831 0 0.0 1e-06 
3.0 2.831 0 0.0 1e-06 
0.05 2.832 0 0.0 1e-06 
3.0 2.832 0 0.0 1e-06 
0.05 2.833 0 0.0 1e-06 
3.0 2.833 0 0.0 1e-06 
0.05 2.834 0 0.0 1e-06 
3.0 2.834 0 0.0 1e-06 
0.05 2.835 0 0.0 1e-06 
3.0 2.835 0 0.0 1e-06 
0.05 2.836 0 0.0 1e-06 
3.0 2.836 0 0.0 1e-06 
0.05 2.837 0 0.0 1e-06 
3.0 2.837 0 0.0 1e-06 
0.05 2.838 0 0.0 1e-06 
3.0 2.838 0 0.0 1e-06 
0.05 2.839 0 0.0 1e-06 
3.0 2.839 0 0.0 1e-06 
0.05 2.84 0 0.0 1e-06 
3.0 2.84 0 0.0 1e-06 
0.05 2.841 0 0.0 1e-06 
3.0 2.841 0 0.0 1e-06 
0.05 2.842 0 0.0 1e-06 
3.0 2.842 0 0.0 1e-06 
0.05 2.843 0 0.0 1e-06 
3.0 2.843 0 0.0 1e-06 
0.05 2.844 0 0.0 1e-06 
3.0 2.844 0 0.0 1e-06 
0.05 2.845 0 0.0 1e-06 
3.0 2.845 0 0.0 1e-06 
0.05 2.846 0 0.0 1e-06 
3.0 2.846 0 0.0 1e-06 
0.05 2.847 0 0.0 1e-06 
3.0 2.847 0 0.0 1e-06 
0.05 2.848 0 0.0 1e-06 
3.0 2.848 0 0.0 1e-06 
0.05 2.849 0 0.0 1e-06 
3.0 2.849 0 0.0 1e-06 
0.05 2.85 0 0.0 1e-06 
3.0 2.85 0 0.0 1e-06 
0.05 2.851 0 0.0 1e-06 
3.0 2.851 0 0.0 1e-06 
0.05 2.852 0 0.0 1e-06 
3.0 2.852 0 0.0 1e-06 
0.05 2.853 0 0.0 1e-06 
3.0 2.853 0 0.0 1e-06 
0.05 2.854 0 0.0 1e-06 
3.0 2.854 0 0.0 1e-06 
0.05 2.855 0 0.0 1e-06 
3.0 2.855 0 0.0 1e-06 
0.05 2.856 0 0.0 1e-06 
3.0 2.856 0 0.0 1e-06 
0.05 2.857 0 0.0 1e-06 
3.0 2.857 0 0.0 1e-06 
0.05 2.858 0 0.0 1e-06 
3.0 2.858 0 0.0 1e-06 
0.05 2.859 0 0.0 1e-06 
3.0 2.859 0 0.0 1e-06 
0.05 2.86 0 0.0 1e-06 
3.0 2.86 0 0.0 1e-06 
0.05 2.861 0 0.0 1e-06 
3.0 2.861 0 0.0 1e-06 
0.05 2.862 0 0.0 1e-06 
3.0 2.862 0 0.0 1e-06 
0.05 2.863 0 0.0 1e-06 
3.0 2.863 0 0.0 1e-06 
0.05 2.864 0 0.0 1e-06 
3.0 2.864 0 0.0 1e-06 
0.05 2.865 0 0.0 1e-06 
3.0 2.865 0 0.0 1e-06 
0.05 2.866 0 0.0 1e-06 
3.0 2.866 0 0.0 1e-06 
0.05 2.867 0 0.0 1e-06 
3.0 2.867 0 0.0 1e-06 
0.05 2.868 0 0.0 1e-06 
3.0 2.868 0 0.0 1e-06 
0.05 2.869 0 0.0 1e-06 
3.0 2.869 0 0.0 1e-06 
0.05 2.87 0 0.0 1e-06 
3.0 2.87 0 0.0 1e-06 
0.05 2.871 0 0.0 1e-06 
3.0 2.871 0 0.0 1e-06 
0.05 2.872 0 0.0 1e-06 
3.0 2.872 0 0.0 1e-06 
0.05 2.873 0 0.0 1e-06 
3.0 2.873 0 0.0 1e-06 
0.05 2.874 0 0.0 1e-06 
3.0 2.874 0 0.0 1e-06 
0.05 2.875 0 0.0 1e-06 
3.0 2.875 0 0.0 1e-06 
0.05 2.876 0 0.0 1e-06 
3.0 2.876 0 0.0 1e-06 
0.05 2.877 0 0.0 1e-06 
3.0 2.877 0 0.0 1e-06 
0.05 2.878 0 0.0 1e-06 
3.0 2.878 0 0.0 1e-06 
0.05 2.879 0 0.0 1e-06 
3.0 2.879 0 0.0 1e-06 
0.05 2.88 0 0.0 1e-06 
3.0 2.88 0 0.0 1e-06 
0.05 2.881 0 0.0 1e-06 
3.0 2.881 0 0.0 1e-06 
0.05 2.882 0 0.0 1e-06 
3.0 2.882 0 0.0 1e-06 
0.05 2.883 0 0.0 1e-06 
3.0 2.883 0 0.0 1e-06 
0.05 2.884 0 0.0 1e-06 
3.0 2.884 0 0.0 1e-06 
0.05 2.885 0 0.0 1e-06 
3.0 2.885 0 0.0 1e-06 
0.05 2.886 0 0.0 1e-06 
3.0 2.886 0 0.0 1e-06 
0.05 2.887 0 0.0 1e-06 
3.0 2.887 0 0.0 1e-06 
0.05 2.888 0 0.0 1e-06 
3.0 2.888 0 0.0 1e-06 
0.05 2.889 0 0.0 1e-06 
3.0 2.889 0 0.0 1e-06 
0.05 2.89 0 0.0 1e-06 
3.0 2.89 0 0.0 1e-06 
0.05 2.891 0 0.0 1e-06 
3.0 2.891 0 0.0 1e-06 
0.05 2.892 0 0.0 1e-06 
3.0 2.892 0 0.0 1e-06 
0.05 2.893 0 0.0 1e-06 
3.0 2.893 0 0.0 1e-06 
0.05 2.894 0 0.0 1e-06 
3.0 2.894 0 0.0 1e-06 
0.05 2.895 0 0.0 1e-06 
3.0 2.895 0 0.0 1e-06 
0.05 2.896 0 0.0 1e-06 
3.0 2.896 0 0.0 1e-06 
0.05 2.897 0 0.0 1e-06 
3.0 2.897 0 0.0 1e-06 
0.05 2.898 0 0.0 1e-06 
3.0 2.898 0 0.0 1e-06 
0.05 2.899 0 0.0 1e-06 
3.0 2.899 0 0.0 1e-06 
0.05 2.9 0 0.0 1e-06 
3.0 2.9 0 0.0 1e-06 
0.05 2.901 0 0.0 1e-06 
3.0 2.901 0 0.0 1e-06 
0.05 2.902 0 0.0 1e-06 
3.0 2.902 0 0.0 1e-06 
0.05 2.903 0 0.0 1e-06 
3.0 2.903 0 0.0 1e-06 
0.05 2.904 0 0.0 1e-06 
3.0 2.904 0 0.0 1e-06 
0.05 2.905 0 0.0 1e-06 
3.0 2.905 0 0.0 1e-06 
0.05 2.906 0 0.0 1e-06 
3.0 2.906 0 0.0 1e-06 
0.05 2.907 0 0.0 1e-06 
3.0 2.907 0 0.0 1e-06 
0.05 2.908 0 0.0 1e-06 
3.0 2.908 0 0.0 1e-06 
0.05 2.909 0 0.0 1e-06 
3.0 2.909 0 0.0 1e-06 
0.05 2.91 0 0.0 1e-06 
3.0 2.91 0 0.0 1e-06 
0.05 2.911 0 0.0 1e-06 
3.0 2.911 0 0.0 1e-06 
0.05 2.912 0 0.0 1e-06 
3.0 2.912 0 0.0 1e-06 
0.05 2.913 0 0.0 1e-06 
3.0 2.913 0 0.0 1e-06 
0.05 2.914 0 0.0 1e-06 
3.0 2.914 0 0.0 1e-06 
0.05 2.915 0 0.0 1e-06 
3.0 2.915 0 0.0 1e-06 
0.05 2.916 0 0.0 1e-06 
3.0 2.916 0 0.0 1e-06 
0.05 2.917 0 0.0 1e-06 
3.0 2.917 0 0.0 1e-06 
0.05 2.918 0 0.0 1e-06 
3.0 2.918 0 0.0 1e-06 
0.05 2.919 0 0.0 1e-06 
3.0 2.919 0 0.0 1e-06 
0.05 2.92 0 0.0 1e-06 
3.0 2.92 0 0.0 1e-06 
0.05 2.921 0 0.0 1e-06 
3.0 2.921 0 0.0 1e-06 
0.05 2.922 0 0.0 1e-06 
3.0 2.922 0 0.0 1e-06 
0.05 2.923 0 0.0 1e-06 
3.0 2.923 0 0.0 1e-06 
0.05 2.924 0 0.0 1e-06 
3.0 2.924 0 0.0 1e-06 
0.05 2.925 0 0.0 1e-06 
3.0 2.925 0 0.0 1e-06 
0.05 2.926 0 0.0 1e-06 
3.0 2.926 0 0.0 1e-06 
0.05 2.927 0 0.0 1e-06 
3.0 2.927 0 0.0 1e-06 
0.05 2.928 0 0.0 1e-06 
3.0 2.928 0 0.0 1e-06 
0.05 2.929 0 0.0 1e-06 
3.0 2.929 0 0.0 1e-06 
0.05 2.93 0 0.0 1e-06 
3.0 2.93 0 0.0 1e-06 
0.05 2.931 0 0.0 1e-06 
3.0 2.931 0 0.0 1e-06 
0.05 2.932 0 0.0 1e-06 
3.0 2.932 0 0.0 1e-06 
0.05 2.933 0 0.0 1e-06 
3.0 2.933 0 0.0 1e-06 
0.05 2.934 0 0.0 1e-06 
3.0 2.934 0 0.0 1e-06 
0.05 2.935 0 0.0 1e-06 
3.0 2.935 0 0.0 1e-06 
0.05 2.936 0 0.0 1e-06 
3.0 2.936 0 0.0 1e-06 
0.05 2.937 0 0.0 1e-06 
3.0 2.937 0 0.0 1e-06 
0.05 2.938 0 0.0 1e-06 
3.0 2.938 0 0.0 1e-06 
0.05 2.939 0 0.0 1e-06 
3.0 2.939 0 0.0 1e-06 
0.05 2.94 0 0.0 1e-06 
3.0 2.94 0 0.0 1e-06 
0.05 2.941 0 0.0 1e-06 
3.0 2.941 0 0.0 1e-06 
0.05 2.942 0 0.0 1e-06 
3.0 2.942 0 0.0 1e-06 
0.05 2.943 0 0.0 1e-06 
3.0 2.943 0 0.0 1e-06 
0.05 2.944 0 0.0 1e-06 
3.0 2.944 0 0.0 1e-06 
0.05 2.945 0 0.0 1e-06 
3.0 2.945 0 0.0 1e-06 
0.05 2.946 0 0.0 1e-06 
3.0 2.946 0 0.0 1e-06 
0.05 2.947 0 0.0 1e-06 
3.0 2.947 0 0.0 1e-06 
0.05 2.948 0 0.0 1e-06 
3.0 2.948 0 0.0 1e-06 
0.05 2.949 0 0.0 1e-06 
3.0 2.949 0 0.0 1e-06 
0.05 2.95 0 0.0 1e-06 
3.0 2.95 0 0.0 1e-06 
0.05 2.951 0 0.0 1e-06 
3.0 2.951 0 0.0 1e-06 
0.05 2.952 0 0.0 1e-06 
3.0 2.952 0 0.0 1e-06 
0.05 2.953 0 0.0 1e-06 
3.0 2.953 0 0.0 1e-06 
0.05 2.954 0 0.0 1e-06 
3.0 2.954 0 0.0 1e-06 
0.05 2.955 0 0.0 1e-06 
3.0 2.955 0 0.0 1e-06 
0.05 2.956 0 0.0 1e-06 
3.0 2.956 0 0.0 1e-06 
0.05 2.957 0 0.0 1e-06 
3.0 2.957 0 0.0 1e-06 
0.05 2.958 0 0.0 1e-06 
3.0 2.958 0 0.0 1e-06 
0.05 2.959 0 0.0 1e-06 
3.0 2.959 0 0.0 1e-06 
0.05 2.96 0 0.0 1e-06 
3.0 2.96 0 0.0 1e-06 
0.05 2.961 0 0.0 1e-06 
3.0 2.961 0 0.0 1e-06 
0.05 2.962 0 0.0 1e-06 
3.0 2.962 0 0.0 1e-06 
0.05 2.963 0 0.0 1e-06 
3.0 2.963 0 0.0 1e-06 
0.05 2.964 0 0.0 1e-06 
3.0 2.964 0 0.0 1e-06 
0.05 2.965 0 0.0 1e-06 
3.0 2.965 0 0.0 1e-06 
0.05 2.966 0 0.0 1e-06 
3.0 2.966 0 0.0 1e-06 
0.05 2.967 0 0.0 1e-06 
3.0 2.967 0 0.0 1e-06 
0.05 2.968 0 0.0 1e-06 
3.0 2.968 0 0.0 1e-06 
0.05 2.969 0 0.0 1e-06 
3.0 2.969 0 0.0 1e-06 
0.05 2.97 0 0.0 1e-06 
3.0 2.97 0 0.0 1e-06 
0.05 2.971 0 0.0 1e-06 
3.0 2.971 0 0.0 1e-06 
0.05 2.972 0 0.0 1e-06 
3.0 2.972 0 0.0 1e-06 
0.05 2.973 0 0.0 1e-06 
3.0 2.973 0 0.0 1e-06 
0.05 2.974 0 0.0 1e-06 
3.0 2.974 0 0.0 1e-06 
0.05 2.975 0 0.0 1e-06 
3.0 2.975 0 0.0 1e-06 
0.05 2.976 0 0.0 1e-06 
3.0 2.976 0 0.0 1e-06 
0.05 2.977 0 0.0 1e-06 
3.0 2.977 0 0.0 1e-06 
0.05 2.978 0 0.0 1e-06 
3.0 2.978 0 0.0 1e-06 
0.05 2.979 0 0.0 1e-06 
3.0 2.979 0 0.0 1e-06 
0.05 2.98 0 0.0 1e-06 
3.0 2.98 0 0.0 1e-06 
0.05 2.981 0 0.0 1e-06 
3.0 2.981 0 0.0 1e-06 
0.05 2.982 0 0.0 1e-06 
3.0 2.982 0 0.0 1e-06 
0.05 2.983 0 0.0 1e-06 
3.0 2.983 0 0.0 1e-06 
0.05 2.984 0 0.0 1e-06 
3.0 2.984 0 0.0 1e-06 
0.05 2.985 0 0.0 1e-06 
3.0 2.985 0 0.0 1e-06 
0.05 2.986 0 0.0 1e-06 
3.0 2.986 0 0.0 1e-06 
0.05 2.987 0 0.0 1e-06 
3.0 2.987 0 0.0 1e-06 
0.05 2.988 0 0.0 1e-06 
3.0 2.988 0 0.0 1e-06 
0.05 2.989 0 0.0 1e-06 
3.0 2.989 0 0.0 1e-06 
0.05 2.99 0 0.0 1e-06 
3.0 2.99 0 0.0 1e-06 
0.05 2.991 0 0.0 1e-06 
3.0 2.991 0 0.0 1e-06 
0.05 2.992 0 0.0 1e-06 
3.0 2.992 0 0.0 1e-06 
0.05 2.993 0 0.0 1e-06 
3.0 2.993 0 0.0 1e-06 
0.05 2.994 0 0.0 1e-06 
3.0 2.994 0 0.0 1e-06 
0.05 2.995 0 0.0 1e-06 
3.0 2.995 0 0.0 1e-06 
0.05 2.996 0 0.0 1e-06 
3.0 2.996 0 0.0 1e-06 
0.05 2.997 0 0.0 1e-06 
3.0 2.997 0 0.0 1e-06 
0.05 2.998 0 0.0 1e-06 
3.0 2.998 0 0.0 1e-06 
0.05 2.999 0 0.0 1e-06 
3.0 2.999 0 0.0 1e-06 
0.05 3.0 0 0.0 1e-06 
3.0 3.0 0 0.0 1e-06 
0.05 3.001 0 0.0 1e-06 
3.0 3.001 0 0.0 1e-06 
0.05 3.002 0 0.0 1e-06 
3.0 3.002 0 0.0 1e-06 
0.05 3.003 0 0.0 1e-06 
3.0 3.003 0 0.0 1e-06 
0.05 3.004 0 0.0 1e-06 
3.0 3.004 0 0.0 1e-06 
0.05 3.005 0 0.0 1e-06 
3.0 3.005 0 0.0 1e-06 
0.05 3.006 0 0.0 1e-06 
3.0 3.006 0 0.0 1e-06 
0.05 3.007 0 0.0 1e-06 
3.0 3.007 0 0.0 1e-06 
0.05 3.008 0 0.0 1e-06 
3.0 3.008 0 0.0 1e-06 
0.05 3.009 0 0.0 1e-06 
3.0 3.009 0 0.0 1e-06 
0.05 3.01 0 0.0 1e-06 
3.0 3.01 0 0.0 1e-06 
0.05 3.011 0 0.0 1e-06 
3.0 3.011 0 0.0 1e-06 
0.05 3.012 0 0.0 1e-06 
3.0 3.012 0 0.0 1e-06 
0.05 3.013 0 0.0 1e-06 
3.0 3.013 0 0.0 1e-06 
0.05 3.014 0 0.0 1e-06 
3.0 3.014 0 0.0 1e-06 
0.05 3.015 0 0.0 1e-06 
3.0 3.015 0 0.0 1e-06 
0.05 3.016 0 0.0 1e-06 
3.0 3.016 0 0.0 1e-06 
0.05 3.017 0 0.0 1e-06 
3.0 3.017 0 0.0 1e-06 
0.05 3.018 0 0.0 1e-06 
3.0 3.018 0 0.0 1e-06 
0.05 3.019 0 0.0 1e-06 
3.0 3.019 0 0.0 1e-06 
0.05 3.02 0 0.0 1e-06 
3.0 3.02 0 0.0 1e-06 
0.05 3.021 0 0.0 1e-06 
3.0 3.021 0 0.0 1e-06 
0.05 3.022 0 0.0 1e-06 
3.0 3.022 0 0.0 1e-06 
0.05 3.023 0 0.0 1e-06 
3.0 3.023 0 0.0 1e-06 
0.05 3.024 0 0.0 1e-06 
3.0 3.024 0 0.0 1e-06 
0.05 3.025 0 0.0 1e-06 
3.0 3.025 0 0.0 1e-06 
0.05 3.026 0 0.0 1e-06 
3.0 3.026 0 0.0 1e-06 
0.05 3.027 0 0.0 1e-06 
3.0 3.027 0 0.0 1e-06 
0.05 3.028 0 0.0 1e-06 
3.0 3.028 0 0.0 1e-06 
0.05 3.029 0 0.0 1e-06 
3.0 3.029 0 0.0 1e-06 
0.05 3.03 0 0.0 1e-06 
3.0 3.03 0 0.0 1e-06 
0.05 3.031 0 0.0 1e-06 
3.0 3.031 0 0.0 1e-06 
0.05 3.032 0 0.0 1e-06 
3.0 3.032 0 0.0 1e-06 
0.05 3.033 0 0.0 1e-06 
3.0 3.033 0 0.0 1e-06 
0.05 3.034 0 0.0 1e-06 
3.0 3.034 0 0.0 1e-06 
0.05 3.035 0 0.0 1e-06 
3.0 3.035 0 0.0 1e-06 
0.05 3.036 0 0.0 1e-06 
3.0 3.036 0 0.0 1e-06 
0.05 3.037 0 0.0 1e-06 
3.0 3.037 0 0.0 1e-06 
0.05 3.038 0 0.0 1e-06 
3.0 3.038 0 0.0 1e-06 
0.05 3.039 0 0.0 1e-06 
3.0 3.039 0 0.0 1e-06 
0.05 3.04 0 0.0 1e-06 
3.0 3.04 0 0.0 1e-06 
0.05 3.041 0 0.0 1e-06 
3.0 3.041 0 0.0 1e-06 
0.05 3.042 0 0.0 1e-06 
3.0 3.042 0 0.0 1e-06 
0.05 3.043 0 0.0 1e-06 
3.0 3.043 0 0.0 1e-06 
0.05 3.044 0 0.0 1e-06 
3.0 3.044 0 0.0 1e-06 
0.05 3.045 0 0.0 1e-06 
3.0 3.045 0 0.0 1e-06 
0.05 3.046 0 0.0 1e-06 
3.0 3.046 0 0.0 1e-06 
0.05 3.047 0 0.0 1e-06 
3.0 3.047 0 0.0 1e-06 
0.05 3.048 0 0.0 1e-06 
3.0 3.048 0 0.0 1e-06 
0.05 3.049 0 0.0 1e-06 
3.0 3.049 0 0.0 1e-06 
0.05 3.05 0 0.0 1e-06 
3.0 3.05 0 0.0 1e-06 
0.05 3.051 0 0.0 1e-06 
3.0 3.051 0 0.0 1e-06 
0.05 3.052 0 0.0 1e-06 
3.0 3.052 0 0.0 1e-06 
0.05 3.053 0 0.0 1e-06 
3.0 3.053 0 0.0 1e-06 
0.05 3.054 0 0.0 1e-06 
3.0 3.054 0 0.0 1e-06 
0.05 3.055 0 0.0 1e-06 
3.0 3.055 0 0.0 1e-06 
0.05 3.056 0 0.0 1e-06 
3.0 3.056 0 0.0 1e-06 
0.05 3.057 0 0.0 1e-06 
3.0 3.057 0 0.0 1e-06 
0.05 3.058 0 0.0 1e-06 
3.0 3.058 0 0.0 1e-06 
0.05 3.059 0 0.0 1e-06 
3.0 3.059 0 0.0 1e-06 
0.05 3.06 0 0.0 1e-06 
3.0 3.06 0 0.0 1e-06 
0.05 3.061 0 0.0 1e-06 
3.0 3.061 0 0.0 1e-06 
0.05 3.062 0 0.0 1e-06 
3.0 3.062 0 0.0 1e-06 
0.05 3.063 0 0.0 1e-06 
3.0 3.063 0 0.0 1e-06 
0.05 3.064 0 0.0 1e-06 
3.0 3.064 0 0.0 1e-06 
0.05 3.065 0 0.0 1e-06 
3.0 3.065 0 0.0 1e-06 
0.05 3.066 0 0.0 1e-06 
3.0 3.066 0 0.0 1e-06 
0.05 3.067 0 0.0 1e-06 
3.0 3.067 0 0.0 1e-06 
0.05 3.068 0 0.0 1e-06 
3.0 3.068 0 0.0 1e-06 
0.05 3.069 0 0.0 1e-06 
3.0 3.069 0 0.0 1e-06 
0.05 3.07 0 0.0 1e-06 
3.0 3.07 0 0.0 1e-06 
0.05 3.071 0 0.0 1e-06 
3.0 3.071 0 0.0 1e-06 
0.05 3.072 0 0.0 1e-06 
3.0 3.072 0 0.0 1e-06 
0.05 3.073 0 0.0 1e-06 
3.0 3.073 0 0.0 1e-06 
0.05 3.074 0 0.0 1e-06 
3.0 3.074 0 0.0 1e-06 
0.05 3.075 0 0.0 1e-06 
3.0 3.075 0 0.0 1e-06 
0.05 3.076 0 0.0 1e-06 
3.0 3.076 0 0.0 1e-06 
0.05 3.077 0 0.0 1e-06 
3.0 3.077 0 0.0 1e-06 
0.05 3.078 0 0.0 1e-06 
3.0 3.078 0 0.0 1e-06 
0.05 3.079 0 0.0 1e-06 
3.0 3.079 0 0.0 1e-06 
0.05 3.08 0 0.0 1e-06 
3.0 3.08 0 0.0 1e-06 
0.05 3.081 0 0.0 1e-06 
3.0 3.081 0 0.0 1e-06 
0.05 3.082 0 0.0 1e-06 
3.0 3.082 0 0.0 1e-06 
0.05 3.083 0 0.0 1e-06 
3.0 3.083 0 0.0 1e-06 
0.05 3.084 0 0.0 1e-06 
3.0 3.084 0 0.0 1e-06 
0.05 3.085 0 0.0 1e-06 
3.0 3.085 0 0.0 1e-06 
0.05 3.086 0 0.0 1e-06 
3.0 3.086 0 0.0 1e-06 
0.05 3.087 0 0.0 1e-06 
3.0 3.087 0 0.0 1e-06 
0.05 3.088 0 0.0 1e-06 
3.0 3.088 0 0.0 1e-06 
0.05 3.089 0 0.0 1e-06 
3.0 3.089 0 0.0 1e-06 
0.05 3.09 0 0.0 1e-06 
3.0 3.09 0 0.0 1e-06 
0.05 3.091 0 0.0 1e-06 
3.0 3.091 0 0.0 1e-06 
0.05 3.092 0 0.0 1e-06 
3.0 3.092 0 0.0 1e-06 
0.05 3.093 0 0.0 1e-06 
3.0 3.093 0 0.0 1e-06 
0.05 3.094 0 0.0 1e-06 
3.0 3.094 0 0.0 1e-06 
0.05 3.095 0 0.0 1e-06 
3.0 3.095 0 0.0 1e-06 
0.05 3.096 0 0.0 1e-06 
3.0 3.096 0 0.0 1e-06 
0.05 3.097 0 0.0 1e-06 
3.0 3.097 0 0.0 1e-06 
0.05 3.098 0 0.0 1e-06 
3.0 3.098 0 0.0 1e-06 
0.05 3.099 0 0.0 1e-06 
3.0 3.099 0 0.0 1e-06 
0.05 3.1 0 0.0 1e-06 
3.0 3.1 0 0.0 1e-06 
0.05 3.101 0 0.0 1e-06 
3.0 3.101 0 0.0 1e-06 
0.05 3.102 0 0.0 1e-06 
3.0 3.102 0 0.0 1e-06 
0.05 3.103 0 0.0 1e-06 
3.0 3.103 0 0.0 1e-06 
0.05 3.104 0 0.0 1e-06 
3.0 3.104 0 0.0 1e-06 
0.05 3.105 0 0.0 1e-06 
3.0 3.105 0 0.0 1e-06 
0.05 3.106 0 0.0 1e-06 
3.0 3.106 0 0.0 1e-06 
0.05 3.107 0 0.0 1e-06 
3.0 3.107 0 0.0 1e-06 
0.05 3.108 0 0.0 1e-06 
3.0 3.108 0 0.0 1e-06 
0.05 3.109 0 0.0 1e-06 
3.0 3.109 0 0.0 1e-06 
0.05 3.11 0 0.0 1e-06 
3.0 3.11 0 0.0 1e-06 
0.05 3.111 0 0.0 1e-06 
3.0 3.111 0 0.0 1e-06 
0.05 3.112 0 0.0 1e-06 
3.0 3.112 0 0.0 1e-06 
0.05 3.113 0 0.0 1e-06 
3.0 3.113 0 0.0 1e-06 
0.05 3.114 0 0.0 1e-06 
3.0 3.114 0 0.0 1e-06 
0.05 3.115 0 0.0 1e-06 
3.0 3.115 0 0.0 1e-06 
0.05 3.116 0 0.0 1e-06 
3.0 3.116 0 0.0 1e-06 
0.05 3.117 0 0.0 1e-06 
3.0 3.117 0 0.0 1e-06 
0.05 3.118 0 0.0 1e-06 
3.0 3.118 0 0.0 1e-06 
0.05 3.119 0 0.0 1e-06 
3.0 3.119 0 0.0 1e-06 
0.05 3.12 0 0.0 1e-06 
3.0 3.12 0 0.0 1e-06 
0.05 3.121 0 0.0 1e-06 
3.0 3.121 0 0.0 1e-06 
0.05 3.122 0 0.0 1e-06 
3.0 3.122 0 0.0 1e-06 
0.05 3.123 0 0.0 1e-06 
3.0 3.123 0 0.0 1e-06 
0.05 3.124 0 0.0 1e-06 
3.0 3.124 0 0.0 1e-06 
0.05 3.125 0 0.0 1e-06 
3.0 3.125 0 0.0 1e-06 
0.05 3.126 0 0.0 1e-06 
3.0 3.126 0 0.0 1e-06 
0.05 3.127 0 0.0 1e-06 
3.0 3.127 0 0.0 1e-06 
0.05 3.128 0 0.0 1e-06 
3.0 3.128 0 0.0 1e-06 
0.05 3.129 0 0.0 1e-06 
3.0 3.129 0 0.0 1e-06 
0.05 3.13 0 0.0 1e-06 
3.0 3.13 0 0.0 1e-06 
0.05 3.131 0 0.0 1e-06 
3.0 3.131 0 0.0 1e-06 
0.05 3.132 0 0.0 1e-06 
3.0 3.132 0 0.0 1e-06 
0.05 3.133 0 0.0 1e-06 
3.0 3.133 0 0.0 1e-06 
0.05 3.134 0 0.0 1e-06 
3.0 3.134 0 0.0 1e-06 
0.05 3.135 0 0.0 1e-06 
3.0 3.135 0 0.0 1e-06 
0.05 3.136 0 0.0 1e-06 
3.0 3.136 0 0.0 1e-06 
0.05 3.137 0 0.0 1e-06 
3.0 3.137 0 0.0 1e-06 
0.05 3.138 0 0.0 1e-06 
3.0 3.138 0 0.0 1e-06 
0.05 3.139 0 0.0 1e-06 
3.0 3.139 0 0.0 1e-06 
0.05 3.14 0 0.0 1e-06 
3.0 3.14 0 0.0 1e-06 
0.05 3.141 0 0.0 1e-06 
3.0 3.141 0 0.0 1e-06 
0.05 3.142 0 0.0 1e-06 
3.0 3.142 0 0.0 1e-06 
0.05 3.143 0 0.0 1e-06 
3.0 3.143 0 0.0 1e-06 
0.05 3.144 0 0.0 1e-06 
3.0 3.144 0 0.0 1e-06 
0.05 3.145 0 0.0 1e-06 
3.0 3.145 0 0.0 1e-06 
0.05 3.146 0 0.0 1e-06 
3.0 3.146 0 0.0 1e-06 
0.05 3.147 0 0.0 1e-06 
3.0 3.147 0 0.0 1e-06 
0.05 3.148 0 0.0 1e-06 
3.0 3.148 0 0.0 1e-06 
0.05 3.149 0 0.0 1e-06 
3.0 3.149 0 0.0 1e-06 
0.05 3.15 0 0.0 1e-06 
3.0 3.15 0 0.0 1e-06 
0.05 3.151 0 0.0 1e-06 
3.0 3.151 0 0.0 1e-06 
0.05 3.152 0 0.0 1e-06 
3.0 3.152 0 0.0 1e-06 
0.05 3.153 0 0.0 1e-06 
3.0 3.153 0 0.0 1e-06 
0.05 3.154 0 0.0 1e-06 
3.0 3.154 0 0.0 1e-06 
0.05 3.155 0 0.0 1e-06 
3.0 3.155 0 0.0 1e-06 
0.05 3.156 0 0.0 1e-06 
3.0 3.156 0 0.0 1e-06 
0.05 3.157 0 0.0 1e-06 
3.0 3.157 0 0.0 1e-06 
0.05 3.158 0 0.0 1e-06 
3.0 3.158 0 0.0 1e-06 
0.05 3.159 0 0.0 1e-06 
3.0 3.159 0 0.0 1e-06 
0.05 3.16 0 0.0 1e-06 
3.0 3.16 0 0.0 1e-06 
0.05 3.161 0 0.0 1e-06 
3.0 3.161 0 0.0 1e-06 
0.05 3.162 0 0.0 1e-06 
3.0 3.162 0 0.0 1e-06 
0.05 3.163 0 0.0 1e-06 
3.0 3.163 0 0.0 1e-06 
0.05 3.164 0 0.0 1e-06 
3.0 3.164 0 0.0 1e-06 
0.05 3.165 0 0.0 1e-06 
3.0 3.165 0 0.0 1e-06 
0.05 3.166 0 0.0 1e-06 
3.0 3.166 0 0.0 1e-06 
0.05 3.167 0 0.0 1e-06 
3.0 3.167 0 0.0 1e-06 
0.05 3.168 0 0.0 1e-06 
3.0 3.168 0 0.0 1e-06 
0.05 3.169 0 0.0 1e-06 
3.0 3.169 0 0.0 1e-06 
0.05 3.17 0 0.0 1e-06 
3.0 3.17 0 0.0 1e-06 
0.05 3.171 0 0.0 1e-06 
3.0 3.171 0 0.0 1e-06 
0.05 3.172 0 0.0 1e-06 
3.0 3.172 0 0.0 1e-06 
0.05 3.173 0 0.0 1e-06 
3.0 3.173 0 0.0 1e-06 
0.05 3.174 0 0.0 1e-06 
3.0 3.174 0 0.0 1e-06 
0.05 3.175 0 0.0 1e-06 
3.0 3.175 0 0.0 1e-06 
0.05 3.176 0 0.0 1e-06 
3.0 3.176 0 0.0 1e-06 
0.05 3.177 0 0.0 1e-06 
3.0 3.177 0 0.0 1e-06 
0.05 3.178 0 0.0 1e-06 
3.0 3.178 0 0.0 1e-06 
0.05 3.179 0 0.0 1e-06 
3.0 3.179 0 0.0 1e-06 
0.05 3.18 0 0.0 1e-06 
3.0 3.18 0 0.0 1e-06 
0.05 3.181 0 0.0 1e-06 
3.0 3.181 0 0.0 1e-06 
0.05 3.182 0 0.0 1e-06 
3.0 3.182 0 0.0 1e-06 
0.05 3.183 0 0.0 1e-06 
3.0 3.183 0 0.0 1e-06 
0.05 3.184 0 0.0 1e-06 
3.0 3.184 0 0.0 1e-06 
0.05 3.185 0 0.0 1e-06 
3.0 3.185 0 0.0 1e-06 
0.05 3.186 0 0.0 1e-06 
3.0 3.186 0 0.0 1e-06 
0.05 3.187 0 0.0 1e-06 
3.0 3.187 0 0.0 1e-06 
0.05 3.188 0 0.0 1e-06 
3.0 3.188 0 0.0 1e-06 
0.05 3.189 0 0.0 1e-06 
3.0 3.189 0 0.0 1e-06 
0.05 3.19 0 0.0 1e-06 
3.0 3.19 0 0.0 1e-06 
0.05 3.191 0 0.0 1e-06 
3.0 3.191 0 0.0 1e-06 
0.05 3.192 0 0.0 1e-06 
3.0 3.192 0 0.0 1e-06 
0.05 3.193 0 0.0 1e-06 
3.0 3.193 0 0.0 1e-06 
0.05 3.194 0 0.0 1e-06 
3.0 3.194 0 0.0 1e-06 
0.05 3.195 0 0.0 1e-06 
3.0 3.195 0 0.0 1e-06 
0.05 3.196 0 0.0 1e-06 
3.0 3.196 0 0.0 1e-06 
0.05 3.197 0 0.0 1e-06 
3.0 3.197 0 0.0 1e-06 
0.05 3.198 0 0.0 1e-06 
3.0 3.198 0 0.0 1e-06 
0.05 3.199 0 0.0 1e-06 
3.0 3.199 0 0.0 1e-06 
0.05 3.2 0 0.0 1e-06 
3.0 3.2 0 0.0 1e-06 
0.05 3.201 0 0.0 1e-06 
3.0 3.201 0 0.0 1e-06 
0.05 3.202 0 0.0 1e-06 
3.0 3.202 0 0.0 1e-06 
0.05 3.203 0 0.0 1e-06 
3.0 3.203 0 0.0 1e-06 
0.05 3.204 0 0.0 1e-06 
3.0 3.204 0 0.0 1e-06 
0.05 3.205 0 0.0 1e-06 
3.0 3.205 0 0.0 1e-06 
0.05 3.206 0 0.0 1e-06 
3.0 3.206 0 0.0 1e-06 
0.05 3.207 0 0.0 1e-06 
3.0 3.207 0 0.0 1e-06 
0.05 3.208 0 0.0 1e-06 
3.0 3.208 0 0.0 1e-06 
0.05 3.209 0 0.0 1e-06 
3.0 3.209 0 0.0 1e-06 
0.05 3.21 0 0.0 1e-06 
3.0 3.21 0 0.0 1e-06 
0.05 3.211 0 0.0 1e-06 
3.0 3.211 0 0.0 1e-06 
0.05 3.212 0 0.0 1e-06 
3.0 3.212 0 0.0 1e-06 
0.05 3.213 0 0.0 1e-06 
3.0 3.213 0 0.0 1e-06 
0.05 3.214 0 0.0 1e-06 
3.0 3.214 0 0.0 1e-06 
0.05 3.215 0 0.0 1e-06 
3.0 3.215 0 0.0 1e-06 
0.05 3.216 0 0.0 1e-06 
3.0 3.216 0 0.0 1e-06 
0.05 3.217 0 0.0 1e-06 
3.0 3.217 0 0.0 1e-06 
0.05 3.218 0 0.0 1e-06 
3.0 3.218 0 0.0 1e-06 
0.05 3.219 0 0.0 1e-06 
3.0 3.219 0 0.0 1e-06 
0.05 3.22 0 0.0 1e-06 
3.0 3.22 0 0.0 1e-06 
0.05 3.221 0 0.0 1e-06 
3.0 3.221 0 0.0 1e-06 
0.05 3.222 0 0.0 1e-06 
3.0 3.222 0 0.0 1e-06 
0.05 3.223 0 0.0 1e-06 
3.0 3.223 0 0.0 1e-06 
0.05 3.224 0 0.0 1e-06 
3.0 3.224 0 0.0 1e-06 
0.05 3.225 0 0.0 1e-06 
3.0 3.225 0 0.0 1e-06 
0.05 3.226 0 0.0 1e-06 
3.0 3.226 0 0.0 1e-06 
0.05 3.227 0 0.0 1e-06 
3.0 3.227 0 0.0 1e-06 
0.05 3.228 0 0.0 1e-06 
3.0 3.228 0 0.0 1e-06 
0.05 3.229 0 0.0 1e-06 
3.0 3.229 0 0.0 1e-06 
0.05 3.23 0 0.0 1e-06 
3.0 3.23 0 0.0 1e-06 
0.05 3.231 0 0.0 1e-06 
3.0 3.231 0 0.0 1e-06 
0.05 3.232 0 0.0 1e-06 
3.0 3.232 0 0.0 1e-06 
0.05 3.233 0 0.0 1e-06 
3.0 3.233 0 0.0 1e-06 
0.05 3.234 0 0.0 1e-06 
3.0 3.234 0 0.0 1e-06 
0.05 3.235 0 0.0 1e-06 
3.0 3.235 0 0.0 1e-06 
0.05 3.236 0 0.0 1e-06 
3.0 3.236 0 0.0 1e-06 
0.05 3.237 0 0.0 1e-06 
3.0 3.237 0 0.0 1e-06 
0.05 3.238 0 0.0 1e-06 
3.0 3.238 0 0.0 1e-06 
0.05 3.239 0 0.0 1e-06 
3.0 3.239 0 0.0 1e-06 
0.05 3.24 0 0.0 1e-06 
3.0 3.24 0 0.0 1e-06 
0.05 3.241 0 0.0 1e-06 
3.0 3.241 0 0.0 1e-06 
0.05 3.242 0 0.0 1e-06 
3.0 3.242 0 0.0 1e-06 
0.05 3.243 0 0.0 1e-06 
3.0 3.243 0 0.0 1e-06 
0.05 3.244 0 0.0 1e-06 
3.0 3.244 0 0.0 1e-06 
0.05 3.245 0 0.0 1e-06 
3.0 3.245 0 0.0 1e-06 
0.05 3.246 0 0.0 1e-06 
3.0 3.246 0 0.0 1e-06 
0.05 3.247 0 0.0 1e-06 
3.0 3.247 0 0.0 1e-06 
0.05 3.248 0 0.0 1e-06 
3.0 3.248 0 0.0 1e-06 
0.05 3.249 0 0.0 1e-06 
3.0 3.249 0 0.0 1e-06 
0.05 3.25 0 0.0 1e-06 
3.0 3.25 0 0.0 1e-06 
0.05 3.251 0 0.0 1e-06 
3.0 3.251 0 0.0 1e-06 
0.05 3.252 0 0.0 1e-06 
3.0 3.252 0 0.0 1e-06 
0.05 3.253 0 0.0 1e-06 
3.0 3.253 0 0.0 1e-06 
0.05 3.254 0 0.0 1e-06 
3.0 3.254 0 0.0 1e-06 
0.05 3.255 0 0.0 1e-06 
3.0 3.255 0 0.0 1e-06 
0.05 3.256 0 0.0 1e-06 
3.0 3.256 0 0.0 1e-06 
0.05 3.257 0 0.0 1e-06 
3.0 3.257 0 0.0 1e-06 
0.05 3.258 0 0.0 1e-06 
3.0 3.258 0 0.0 1e-06 
0.05 3.259 0 0.0 1e-06 
3.0 3.259 0 0.0 1e-06 
0.05 3.26 0 0.0 1e-06 
3.0 3.26 0 0.0 1e-06 
0.05 3.261 0 0.0 1e-06 
3.0 3.261 0 0.0 1e-06 
0.05 3.262 0 0.0 1e-06 
3.0 3.262 0 0.0 1e-06 
0.05 3.263 0 0.0 1e-06 
3.0 3.263 0 0.0 1e-06 
0.05 3.264 0 0.0 1e-06 
3.0 3.264 0 0.0 1e-06 
0.05 3.265 0 0.0 1e-06 
3.0 3.265 0 0.0 1e-06 
0.05 3.266 0 0.0 1e-06 
3.0 3.266 0 0.0 1e-06 
0.05 3.267 0 0.0 1e-06 
3.0 3.267 0 0.0 1e-06 
0.05 3.268 0 0.0 1e-06 
3.0 3.268 0 0.0 1e-06 
0.05 3.269 0 0.0 1e-06 
3.0 3.269 0 0.0 1e-06 
0.05 3.27 0 0.0 1e-06 
3.0 3.27 0 0.0 1e-06 
0.05 3.271 0 0.0 1e-06 
3.0 3.271 0 0.0 1e-06 
0.05 3.272 0 0.0 1e-06 
3.0 3.272 0 0.0 1e-06 
0.05 3.273 0 0.0 1e-06 
3.0 3.273 0 0.0 1e-06 
0.05 3.274 0 0.0 1e-06 
3.0 3.274 0 0.0 1e-06 
0.05 3.275 0 0.0 1e-06 
3.0 3.275 0 0.0 1e-06 
0.05 3.276 0 0.0 1e-06 
3.0 3.276 0 0.0 1e-06 
0.05 3.277 0 0.0 1e-06 
3.0 3.277 0 0.0 1e-06 
0.05 3.278 0 0.0 1e-06 
3.0 3.278 0 0.0 1e-06 
0.05 3.279 0 0.0 1e-06 
3.0 3.279 0 0.0 1e-06 
0.05 3.28 0 0.0 1e-06 
3.0 3.28 0 0.0 1e-06 
0.05 3.281 0 0.0 1e-06 
3.0 3.281 0 0.0 1e-06 
0.05 3.282 0 0.0 1e-06 
3.0 3.282 0 0.0 1e-06 
0.05 3.283 0 0.0 1e-06 
3.0 3.283 0 0.0 1e-06 
0.05 3.284 0 0.0 1e-06 
3.0 3.284 0 0.0 1e-06 
0.05 3.285 0 0.0 1e-06 
3.0 3.285 0 0.0 1e-06 
0.05 3.286 0 0.0 1e-06 
3.0 3.286 0 0.0 1e-06 
0.05 3.287 0 0.0 1e-06 
3.0 3.287 0 0.0 1e-06 
0.05 3.288 0 0.0 1e-06 
3.0 3.288 0 0.0 1e-06 
0.05 3.289 0 0.0 1e-06 
3.0 3.289 0 0.0 1e-06 
0.05 3.29 0 0.0 1e-06 
3.0 3.29 0 0.0 1e-06 
0.05 3.291 0 0.0 1e-06 
3.0 3.291 0 0.0 1e-06 
0.05 3.292 0 0.0 1e-06 
3.0 3.292 0 0.0 1e-06 
0.05 3.293 0 0.0 1e-06 
3.0 3.293 0 0.0 1e-06 
0.05 3.294 0 0.0 1e-06 
3.0 3.294 0 0.0 1e-06 
0.05 3.295 0 0.0 1e-06 
3.0 3.295 0 0.0 1e-06 
0.05 3.296 0 0.0 1e-06 
3.0 3.296 0 0.0 1e-06 
0.05 3.297 0 0.0 1e-06 
3.0 3.297 0 0.0 1e-06 
0.05 3.298 0 0.0 1e-06 
3.0 3.298 0 0.0 1e-06 
0.05 3.299 0 0.0 1e-06 
3.0 3.299 0 0.0 1e-06 
0.05 3.3 0 0.0 1e-06 
3.0 3.3 0 0.0 1e-06 
0.05 3.301 0 0.0 1e-06 
3.0 3.301 0 0.0 1e-06 
0.05 3.302 0 0.0 1e-06 
3.0 3.302 0 0.0 1e-06 
0.05 3.303 0 0.0 1e-06 
3.0 3.303 0 0.0 1e-06 
0.05 3.304 0 0.0 1e-06 
3.0 3.304 0 0.0 1e-06 
0.05 3.305 0 0.0 1e-06 
3.0 3.305 0 0.0 1e-06 
0.05 3.306 0 0.0 1e-06 
3.0 3.306 0 0.0 1e-06 
0.05 3.307 0 0.0 1e-06 
3.0 3.307 0 0.0 1e-06 
0.05 3.308 0 0.0 1e-06 
3.0 3.308 0 0.0 1e-06 
0.05 3.309 0 0.0 1e-06 
3.0 3.309 0 0.0 1e-06 
0.05 3.31 0 0.0 1e-06 
3.0 3.31 0 0.0 1e-06 
0.05 3.311 0 0.0 1e-06 
3.0 3.311 0 0.0 1e-06 
0.05 3.312 0 0.0 1e-06 
3.0 3.312 0 0.0 1e-06 
0.05 3.313 0 0.0 1e-06 
3.0 3.313 0 0.0 1e-06 
0.05 3.314 0 0.0 1e-06 
3.0 3.314 0 0.0 1e-06 
0.05 3.315 0 0.0 1e-06 
3.0 3.315 0 0.0 1e-06 
0.05 3.316 0 0.0 1e-06 
3.0 3.316 0 0.0 1e-06 
0.05 3.317 0 0.0 1e-06 
3.0 3.317 0 0.0 1e-06 
0.05 3.318 0 0.0 1e-06 
3.0 3.318 0 0.0 1e-06 
0.05 3.319 0 0.0 1e-06 
3.0 3.319 0 0.0 1e-06 
0.05 3.32 0 0.0 1e-06 
3.0 3.32 0 0.0 1e-06 
0.05 3.321 0 0.0 1e-06 
3.0 3.321 0 0.0 1e-06 
0.05 3.322 0 0.0 1e-06 
3.0 3.322 0 0.0 1e-06 
0.05 3.323 0 0.0 1e-06 
3.0 3.323 0 0.0 1e-06 
0.05 3.324 0 0.0 1e-06 
3.0 3.324 0 0.0 1e-06 
0.05 3.325 0 0.0 1e-06 
3.0 3.325 0 0.0 1e-06 
0.05 3.326 0 0.0 1e-06 
3.0 3.326 0 0.0 1e-06 
0.05 3.327 0 0.0 1e-06 
3.0 3.327 0 0.0 1e-06 
0.05 3.328 0 0.0 1e-06 
3.0 3.328 0 0.0 1e-06 
0.05 3.329 0 0.0 1e-06 
3.0 3.329 0 0.0 1e-06 
0.05 3.33 0 0.0 1e-06 
3.0 3.33 0 0.0 1e-06 
0.05 3.331 0 0.0 1e-06 
3.0 3.331 0 0.0 1e-06 
0.05 3.332 0 0.0 1e-06 
3.0 3.332 0 0.0 1e-06 
0.05 3.333 0 0.0 1e-06 
3.0 3.333 0 0.0 1e-06 
0.05 3.334 0 0.0 1e-06 
3.0 3.334 0 0.0 1e-06 
0.05 3.335 0 0.0 1e-06 
3.0 3.335 0 0.0 1e-06 
0.05 3.336 0 0.0 1e-06 
3.0 3.336 0 0.0 1e-06 
0.05 3.337 0 0.0 1e-06 
3.0 3.337 0 0.0 1e-06 
0.05 3.338 0 0.0 1e-06 
3.0 3.338 0 0.0 1e-06 
0.05 3.339 0 0.0 1e-06 
3.0 3.339 0 0.0 1e-06 
0.05 3.34 0 0.0 1e-06 
3.0 3.34 0 0.0 1e-06 
0.05 3.341 0 0.0 1e-06 
3.0 3.341 0 0.0 1e-06 
0.05 3.342 0 0.0 1e-06 
3.0 3.342 0 0.0 1e-06 
0.05 3.343 0 0.0 1e-06 
3.0 3.343 0 0.0 1e-06 
0.05 3.344 0 0.0 1e-06 
3.0 3.344 0 0.0 1e-06 
0.05 3.345 0 0.0 1e-06 
3.0 3.345 0 0.0 1e-06 
0.05 3.346 0 0.0 1e-06 
3.0 3.346 0 0.0 1e-06 
0.05 3.347 0 0.0 1e-06 
3.0 3.347 0 0.0 1e-06 
0.05 3.348 0 0.0 1e-06 
3.0 3.348 0 0.0 1e-06 
0.05 3.349 0 0.0 1e-06 
3.0 3.349 0 0.0 1e-06 
0.05 3.35 0 0.0 1e-06 
3.0 3.35 0 0.0 1e-06 
0.05 3.351 0 0.0 1e-06 
3.0 3.351 0 0.0 1e-06 
0.05 3.352 0 0.0 1e-06 
3.0 3.352 0 0.0 1e-06 
0.05 3.353 0 0.0 1e-06 
3.0 3.353 0 0.0 1e-06 
0.05 3.354 0 0.0 1e-06 
3.0 3.354 0 0.0 1e-06 
0.05 3.355 0 0.0 1e-06 
3.0 3.355 0 0.0 1e-06 
0.05 3.356 0 0.0 1e-06 
3.0 3.356 0 0.0 1e-06 
0.05 3.357 0 0.0 1e-06 
3.0 3.357 0 0.0 1e-06 
0.05 3.358 0 0.0 1e-06 
3.0 3.358 0 0.0 1e-06 
0.05 3.359 0 0.0 1e-06 
3.0 3.359 0 0.0 1e-06 
0.05 3.36 0 0.0 1e-06 
3.0 3.36 0 0.0 1e-06 
0.05 3.361 0 0.0 1e-06 
3.0 3.361 0 0.0 1e-06 
0.05 3.362 0 0.0 1e-06 
3.0 3.362 0 0.0 1e-06 
0.05 3.363 0 0.0 1e-06 
3.0 3.363 0 0.0 1e-06 
0.05 3.364 0 0.0 1e-06 
3.0 3.364 0 0.0 1e-06 
0.05 3.365 0 0.0 1e-06 
3.0 3.365 0 0.0 1e-06 
0.05 3.366 0 0.0 1e-06 
3.0 3.366 0 0.0 1e-06 
0.05 3.367 0 0.0 1e-06 
3.0 3.367 0 0.0 1e-06 
0.05 3.368 0 0.0 1e-06 
3.0 3.368 0 0.0 1e-06 
0.05 3.369 0 0.0 1e-06 
3.0 3.369 0 0.0 1e-06 
0.05 3.37 0 0.0 1e-06 
3.0 3.37 0 0.0 1e-06 
0.05 3.371 0 0.0 1e-06 
3.0 3.371 0 0.0 1e-06 
0.05 3.372 0 0.0 1e-06 
3.0 3.372 0 0.0 1e-06 
0.05 3.373 0 0.0 1e-06 
3.0 3.373 0 0.0 1e-06 
0.05 3.374 0 0.0 1e-06 
3.0 3.374 0 0.0 1e-06 
0.05 3.375 0 0.0 1e-06 
3.0 3.375 0 0.0 1e-06 
0.05 3.376 0 0.0 1e-06 
3.0 3.376 0 0.0 1e-06 
0.05 3.377 0 0.0 1e-06 
3.0 3.377 0 0.0 1e-06 
0.05 3.378 0 0.0 1e-06 
3.0 3.378 0 0.0 1e-06 
0.05 3.379 0 0.0 1e-06 
3.0 3.379 0 0.0 1e-06 
0.05 3.38 0 0.0 1e-06 
3.0 3.38 0 0.0 1e-06 
0.05 3.381 0 0.0 1e-06 
3.0 3.381 0 0.0 1e-06 
0.05 3.382 0 0.0 1e-06 
3.0 3.382 0 0.0 1e-06 
0.05 3.383 0 0.0 1e-06 
3.0 3.383 0 0.0 1e-06 
0.05 3.384 0 0.0 1e-06 
3.0 3.384 0 0.0 1e-06 
0.05 3.385 0 0.0 1e-06 
3.0 3.385 0 0.0 1e-06 
0.05 3.386 0 0.0 1e-06 
3.0 3.386 0 0.0 1e-06 
0.05 3.387 0 0.0 1e-06 
3.0 3.387 0 0.0 1e-06 
0.05 3.388 0 0.0 1e-06 
3.0 3.388 0 0.0 1e-06 
0.05 3.389 0 0.0 1e-06 
3.0 3.389 0 0.0 1e-06 
0.05 3.39 0 0.0 1e-06 
3.0 3.39 0 0.0 1e-06 
0.05 3.391 0 0.0 1e-06 
3.0 3.391 0 0.0 1e-06 
0.05 3.392 0 0.0 1e-06 
3.0 3.392 0 0.0 1e-06 
0.05 3.393 0 0.0 1e-06 
3.0 3.393 0 0.0 1e-06 
0.05 3.394 0 0.0 1e-06 
3.0 3.394 0 0.0 1e-06 
0.05 3.395 0 0.0 1e-06 
3.0 3.395 0 0.0 1e-06 
0.05 3.396 0 0.0 1e-06 
3.0 3.396 0 0.0 1e-06 
0.05 3.397 0 0.0 1e-06 
3.0 3.397 0 0.0 1e-06 
0.05 3.398 0 0.0 1e-06 
3.0 3.398 0 0.0 1e-06 
0.05 3.399 0 0.0 1e-06 
3.0 3.399 0 0.0 1e-06 
0.05 3.4 0 0.0 1e-06 
3.0 3.4 0 0.0 1e-06 
0.05 3.401 0 0.0 1e-06 
3.0 3.401 0 0.0 1e-06 
0.05 3.402 0 0.0 1e-06 
3.0 3.402 0 0.0 1e-06 
0.05 3.403 0 0.0 1e-06 
3.0 3.403 0 0.0 1e-06 
0.05 3.404 0 0.0 1e-06 
3.0 3.404 0 0.0 1e-06 
0.05 3.405 0 0.0 1e-06 
3.0 3.405 0 0.0 1e-06 
0.05 3.406 0 0.0 1e-06 
3.0 3.406 0 0.0 1e-06 
0.05 3.407 0 0.0 1e-06 
3.0 3.407 0 0.0 1e-06 
0.05 3.408 0 0.0 1e-06 
3.0 3.408 0 0.0 1e-06 
0.05 3.409 0 0.0 1e-06 
3.0 3.409 0 0.0 1e-06 
0.05 3.41 0 0.0 1e-06 
3.0 3.41 0 0.0 1e-06 
0.05 3.411 0 0.0 1e-06 
3.0 3.411 0 0.0 1e-06 
0.05 3.412 0 0.0 1e-06 
3.0 3.412 0 0.0 1e-06 
0.05 3.413 0 0.0 1e-06 
3.0 3.413 0 0.0 1e-06 
0.05 3.414 0 0.0 1e-06 
3.0 3.414 0 0.0 1e-06 
0.05 3.415 0 0.0 1e-06 
3.0 3.415 0 0.0 1e-06 
0.05 3.416 0 0.0 1e-06 
3.0 3.416 0 0.0 1e-06 
0.05 3.417 0 0.0 1e-06 
3.0 3.417 0 0.0 1e-06 
0.05 3.418 0 0.0 1e-06 
3.0 3.418 0 0.0 1e-06 
0.05 3.419 0 0.0 1e-06 
3.0 3.419 0 0.0 1e-06 
0.05 3.42 0 0.0 1e-06 
3.0 3.42 0 0.0 1e-06 
0.05 3.421 0 0.0 1e-06 
3.0 3.421 0 0.0 1e-06 
0.05 3.422 0 0.0 1e-06 
3.0 3.422 0 0.0 1e-06 
0.05 3.423 0 0.0 1e-06 
3.0 3.423 0 0.0 1e-06 
0.05 3.424 0 0.0 1e-06 
3.0 3.424 0 0.0 1e-06 
0.05 3.425 0 0.0 1e-06 
3.0 3.425 0 0.0 1e-06 
0.05 3.426 0 0.0 1e-06 
3.0 3.426 0 0.0 1e-06 
0.05 3.427 0 0.0 1e-06 
3.0 3.427 0 0.0 1e-06 
0.05 3.428 0 0.0 1e-06 
3.0 3.428 0 0.0 1e-06 
0.05 3.429 0 0.0 1e-06 
3.0 3.429 0 0.0 1e-06 
0.05 3.43 0 0.0 1e-06 
3.0 3.43 0 0.0 1e-06 
0.05 3.431 0 0.0 1e-06 
3.0 3.431 0 0.0 1e-06 
0.05 3.432 0 0.0 1e-06 
3.0 3.432 0 0.0 1e-06 
0.05 3.433 0 0.0 1e-06 
3.0 3.433 0 0.0 1e-06 
0.05 3.434 0 0.0 1e-06 
3.0 3.434 0 0.0 1e-06 
0.05 3.435 0 0.0 1e-06 
3.0 3.435 0 0.0 1e-06 
0.05 3.436 0 0.0 1e-06 
3.0 3.436 0 0.0 1e-06 
0.05 3.437 0 0.0 1e-06 
3.0 3.437 0 0.0 1e-06 
0.05 3.438 0 0.0 1e-06 
3.0 3.438 0 0.0 1e-06 
0.05 3.439 0 0.0 1e-06 
3.0 3.439 0 0.0 1e-06 
0.05 3.44 0 0.0 1e-06 
3.0 3.44 0 0.0 1e-06 
0.05 3.441 0 0.0 1e-06 
3.0 3.441 0 0.0 1e-06 
0.05 3.442 0 0.0 1e-06 
3.0 3.442 0 0.0 1e-06 
0.05 3.443 0 0.0 1e-06 
3.0 3.443 0 0.0 1e-06 
0.05 3.444 0 0.0 1e-06 
3.0 3.444 0 0.0 1e-06 
0.05 3.445 0 0.0 1e-06 
3.0 3.445 0 0.0 1e-06 
0.05 3.446 0 0.0 1e-06 
3.0 3.446 0 0.0 1e-06 
0.05 3.447 0 0.0 1e-06 
3.0 3.447 0 0.0 1e-06 
0.05 3.448 0 0.0 1e-06 
3.0 3.448 0 0.0 1e-06 
0.05 3.449 0 0.0 1e-06 
3.0 3.449 0 0.0 1e-06 
0.05 3.45 0 0.0 1e-06 
3.0 3.45 0 0.0 1e-06 
0.05 3.451 0 0.0 1e-06 
3.0 3.451 0 0.0 1e-06 
0.05 3.452 0 0.0 1e-06 
3.0 3.452 0 0.0 1e-06 
0.05 3.453 0 0.0 1e-06 
3.0 3.453 0 0.0 1e-06 
0.05 3.454 0 0.0 1e-06 
3.0 3.454 0 0.0 1e-06 
0.05 3.455 0 0.0 1e-06 
3.0 3.455 0 0.0 1e-06 
0.05 3.456 0 0.0 1e-06 
3.0 3.456 0 0.0 1e-06 
0.05 3.457 0 0.0 1e-06 
3.0 3.457 0 0.0 1e-06 
0.05 3.458 0 0.0 1e-06 
3.0 3.458 0 0.0 1e-06 
0.05 3.459 0 0.0 1e-06 
3.0 3.459 0 0.0 1e-06 
0.05 3.46 0 0.0 1e-06 
3.0 3.46 0 0.0 1e-06 
0.05 3.461 0 0.0 1e-06 
3.0 3.461 0 0.0 1e-06 
0.05 3.462 0 0.0 1e-06 
3.0 3.462 0 0.0 1e-06 
0.05 3.463 0 0.0 1e-06 
3.0 3.463 0 0.0 1e-06 
0.05 3.464 0 0.0 1e-06 
3.0 3.464 0 0.0 1e-06 
0.05 3.465 0 0.0 1e-06 
3.0 3.465 0 0.0 1e-06 
0.05 3.466 0 0.0 1e-06 
3.0 3.466 0 0.0 1e-06 
0.05 3.467 0 0.0 1e-06 
3.0 3.467 0 0.0 1e-06 
0.05 3.468 0 0.0 1e-06 
3.0 3.468 0 0.0 1e-06 
0.05 3.469 0 0.0 1e-06 
3.0 3.469 0 0.0 1e-06 
0.05 3.47 0 0.0 1e-06 
3.0 3.47 0 0.0 1e-06 
0.05 3.471 0 0.0 1e-06 
3.0 3.471 0 0.0 1e-06 
0.05 3.472 0 0.0 1e-06 
3.0 3.472 0 0.0 1e-06 
0.05 3.473 0 0.0 1e-06 
3.0 3.473 0 0.0 1e-06 
0.05 3.474 0 0.0 1e-06 
3.0 3.474 0 0.0 1e-06 
0.05 3.475 0 0.0 1e-06 
3.0 3.475 0 0.0 1e-06 
0.05 3.476 0 0.0 1e-06 
3.0 3.476 0 0.0 1e-06 
0.05 3.477 0 0.0 1e-06 
3.0 3.477 0 0.0 1e-06 
0.05 3.478 0 0.0 1e-06 
3.0 3.478 0 0.0 1e-06 
0.05 3.479 0 0.0 1e-06 
3.0 3.479 0 0.0 1e-06 
0.05 3.48 0 0.0 1e-06 
3.0 3.48 0 0.0 1e-06 
0.05 3.481 0 0.0 1e-06 
3.0 3.481 0 0.0 1e-06 
0.05 3.482 0 0.0 1e-06 
3.0 3.482 0 0.0 1e-06 
0.05 3.483 0 0.0 1e-06 
3.0 3.483 0 0.0 1e-06 
0.05 3.484 0 0.0 1e-06 
3.0 3.484 0 0.0 1e-06 
0.05 3.485 0 0.0 1e-06 
3.0 3.485 0 0.0 1e-06 
0.05 3.486 0 0.0 1e-06 
3.0 3.486 0 0.0 1e-06 
0.05 3.487 0 0.0 1e-06 
3.0 3.487 0 0.0 1e-06 
0.05 3.488 0 0.0 1e-06 
3.0 3.488 0 0.0 1e-06 
0.05 3.489 0 0.0 1e-06 
3.0 3.489 0 0.0 1e-06 
0.05 3.49 0 0.0 1e-06 
3.0 3.49 0 0.0 1e-06 
0.05 3.491 0 0.0 1e-06 
3.0 3.491 0 0.0 1e-06 
0.05 3.492 0 0.0 1e-06 
3.0 3.492 0 0.0 1e-06 
0.05 3.493 0 0.0 1e-06 
3.0 3.493 0 0.0 1e-06 
0.05 3.494 0 0.0 1e-06 
3.0 3.494 0 0.0 1e-06 
0.05 3.495 0 0.0 1e-06 
3.0 3.495 0 0.0 1e-06 
0.05 3.496 0 0.0 1e-06 
3.0 3.496 0 0.0 1e-06 
0.05 3.497 0 0.0 1e-06 
3.0 3.497 0 0.0 1e-06 
0.05 3.498 0 0.0 1e-06 
3.0 3.498 0 0.0 1e-06 
0.05 3.499 0 0.0 1e-06 
3.0 3.499 0 0.0 1e-06 
0.05 3.5 0 0.0 1e-06 
3.0 3.5 0 0.0 1e-06 
0.05 3.501 0 0.0 1e-06 
3.0 3.501 0 0.0 1e-06 
0.05 3.502 0 0.0 1e-06 
3.0 3.502 0 0.0 1e-06 
0.05 3.503 0 0.0 1e-06 
3.0 3.503 0 0.0 1e-06 
0.05 3.504 0 0.0 1e-06 
3.0 3.504 0 0.0 1e-06 
0.05 3.505 0 0.0 1e-06 
3.0 3.505 0 0.0 1e-06 
0.05 3.506 0 0.0 1e-06 
3.0 3.506 0 0.0 1e-06 
0.05 3.507 0 0.0 1e-06 
3.0 3.507 0 0.0 1e-06 
0.05 3.508 0 0.0 1e-06 
3.0 3.508 0 0.0 1e-06 
0.05 3.509 0 0.0 1e-06 
3.0 3.509 0 0.0 1e-06 
0.05 3.51 0 0.0 1e-06 
3.0 3.51 0 0.0 1e-06 
0.05 3.511 0 0.0 1e-06 
3.0 3.511 0 0.0 1e-06 
0.05 3.512 0 0.0 1e-06 
3.0 3.512 0 0.0 1e-06 
0.05 3.513 0 0.0 1e-06 
3.0 3.513 0 0.0 1e-06 
0.05 3.514 0 0.0 1e-06 
3.0 3.514 0 0.0 1e-06 
0.05 3.515 0 0.0 1e-06 
3.0 3.515 0 0.0 1e-06 
0.05 3.516 0 0.0 1e-06 
3.0 3.516 0 0.0 1e-06 
0.05 3.517 0 0.0 1e-06 
3.0 3.517 0 0.0 1e-06 
0.05 3.518 0 0.0 1e-06 
3.0 3.518 0 0.0 1e-06 
0.05 3.519 0 0.0 1e-06 
3.0 3.519 0 0.0 1e-06 
0.05 3.52 0 0.0 1e-06 
3.0 3.52 0 0.0 1e-06 
0.05 3.521 0 0.0 1e-06 
3.0 3.521 0 0.0 1e-06 
0.05 3.522 0 0.0 1e-06 
3.0 3.522 0 0.0 1e-06 
0.05 3.523 0 0.0 1e-06 
3.0 3.523 0 0.0 1e-06 
0.05 3.524 0 0.0 1e-06 
3.0 3.524 0 0.0 1e-06 
0.05 3.525 0 0.0 1e-06 
3.0 3.525 0 0.0 1e-06 
0.05 3.526 0 0.0 1e-06 
3.0 3.526 0 0.0 1e-06 
0.05 3.527 0 0.0 1e-06 
3.0 3.527 0 0.0 1e-06 
0.05 3.528 0 0.0 1e-06 
3.0 3.528 0 0.0 1e-06 
0.05 3.529 0 0.0 1e-06 
3.0 3.529 0 0.0 1e-06 
0.05 3.53 0 0.0 1e-06 
3.0 3.53 0 0.0 1e-06 
0.05 3.531 0 0.0 1e-06 
3.0 3.531 0 0.0 1e-06 
0.05 3.532 0 0.0 1e-06 
3.0 3.532 0 0.0 1e-06 
0.05 3.533 0 0.0 1e-06 
3.0 3.533 0 0.0 1e-06 
0.05 3.534 0 0.0 1e-06 
3.0 3.534 0 0.0 1e-06 
0.05 3.535 0 0.0 1e-06 
3.0 3.535 0 0.0 1e-06 
0.05 3.536 0 0.0 1e-06 
3.0 3.536 0 0.0 1e-06 
0.05 3.537 0 0.0 1e-06 
3.0 3.537 0 0.0 1e-06 
0.05 3.538 0 0.0 1e-06 
3.0 3.538 0 0.0 1e-06 
0.05 3.539 0 0.0 1e-06 
3.0 3.539 0 0.0 1e-06 
0.05 3.54 0 0.0 1e-06 
3.0 3.54 0 0.0 1e-06 
0.05 3.541 0 0.0 1e-06 
3.0 3.541 0 0.0 1e-06 
0.05 3.542 0 0.0 1e-06 
3.0 3.542 0 0.0 1e-06 
0.05 3.543 0 0.0 1e-06 
3.0 3.543 0 0.0 1e-06 
0.05 3.544 0 0.0 1e-06 
3.0 3.544 0 0.0 1e-06 
0.05 3.545 0 0.0 1e-06 
3.0 3.545 0 0.0 1e-06 
0.05 3.546 0 0.0 1e-06 
3.0 3.546 0 0.0 1e-06 
0.05 3.547 0 0.0 1e-06 
3.0 3.547 0 0.0 1e-06 
0.05 3.548 0 0.0 1e-06 
3.0 3.548 0 0.0 1e-06 
0.05 3.549 0 0.0 1e-06 
3.0 3.549 0 0.0 1e-06 
0.05 3.55 0 0.0 1e-06 
3.0 3.55 0 0.0 1e-06 
0.05 3.551 0 0.0 1e-06 
3.0 3.551 0 0.0 1e-06 
0.05 3.552 0 0.0 1e-06 
3.0 3.552 0 0.0 1e-06 
0.05 3.553 0 0.0 1e-06 
3.0 3.553 0 0.0 1e-06 
0.05 3.554 0 0.0 1e-06 
3.0 3.554 0 0.0 1e-06 
0.05 3.555 0 0.0 1e-06 
3.0 3.555 0 0.0 1e-06 
0.05 3.556 0 0.0 1e-06 
3.0 3.556 0 0.0 1e-06 
0.05 3.557 0 0.0 1e-06 
3.0 3.557 0 0.0 1e-06 
0.05 3.558 0 0.0 1e-06 
3.0 3.558 0 0.0 1e-06 
0.05 3.559 0 0.0 1e-06 
3.0 3.559 0 0.0 1e-06 
0.05 3.56 0 0.0 1e-06 
3.0 3.56 0 0.0 1e-06 
0.05 3.561 0 0.0 1e-06 
3.0 3.561 0 0.0 1e-06 
0.05 3.562 0 0.0 1e-06 
3.0 3.562 0 0.0 1e-06 
0.05 3.563 0 0.0 1e-06 
3.0 3.563 0 0.0 1e-06 
0.05 3.564 0 0.0 1e-06 
3.0 3.564 0 0.0 1e-06 
0.05 3.565 0 0.0 1e-06 
3.0 3.565 0 0.0 1e-06 
0.05 3.566 0 0.0 1e-06 
3.0 3.566 0 0.0 1e-06 
0.05 3.567 0 0.0 1e-06 
3.0 3.567 0 0.0 1e-06 
0.05 3.568 0 0.0 1e-06 
3.0 3.568 0 0.0 1e-06 
0.05 3.569 0 0.0 1e-06 
3.0 3.569 0 0.0 1e-06 
0.05 3.57 0 0.0 1e-06 
3.0 3.57 0 0.0 1e-06 
0.05 3.571 0 0.0 1e-06 
3.0 3.571 0 0.0 1e-06 
0.05 3.572 0 0.0 1e-06 
3.0 3.572 0 0.0 1e-06 
0.05 3.573 0 0.0 1e-06 
3.0 3.573 0 0.0 1e-06 
0.05 3.574 0 0.0 1e-06 
3.0 3.574 0 0.0 1e-06 
0.05 3.575 0 0.0 1e-06 
3.0 3.575 0 0.0 1e-06 
0.05 3.576 0 0.0 1e-06 
3.0 3.576 0 0.0 1e-06 
0.05 3.577 0 0.0 1e-06 
3.0 3.577 0 0.0 1e-06 
0.05 3.578 0 0.0 1e-06 
3.0 3.578 0 0.0 1e-06 
0.05 3.579 0 0.0 1e-06 
3.0 3.579 0 0.0 1e-06 
0.05 3.58 0 0.0 1e-06 
3.0 3.58 0 0.0 1e-06 
0.05 3.581 0 0.0 1e-06 
3.0 3.581 0 0.0 1e-06 
0.05 3.582 0 0.0 1e-06 
3.0 3.582 0 0.0 1e-06 
0.05 3.583 0 0.0 1e-06 
3.0 3.583 0 0.0 1e-06 
0.05 3.584 0 0.0 1e-06 
3.0 3.584 0 0.0 1e-06 
0.05 3.585 0 0.0 1e-06 
3.0 3.585 0 0.0 1e-06 
0.05 3.586 0 0.0 1e-06 
3.0 3.586 0 0.0 1e-06 
0.05 3.587 0 0.0 1e-06 
3.0 3.587 0 0.0 1e-06 
0.05 3.588 0 0.0 1e-06 
3.0 3.588 0 0.0 1e-06 
0.05 3.589 0 0.0 1e-06 
3.0 3.589 0 0.0 1e-06 
0.05 3.59 0 0.0 1e-06 
3.0 3.59 0 0.0 1e-06 
0.05 3.591 0 0.0 1e-06 
3.0 3.591 0 0.0 1e-06 
0.05 3.592 0 0.0 1e-06 
3.0 3.592 0 0.0 1e-06 
0.05 3.593 0 0.0 1e-06 
3.0 3.593 0 0.0 1e-06 
0.05 3.594 0 0.0 1e-06 
3.0 3.594 0 0.0 1e-06 
0.05 3.595 0 0.0 1e-06 
3.0 3.595 0 0.0 1e-06 
0.05 3.596 0 0.0 1e-06 
3.0 3.596 0 0.0 1e-06 
0.05 3.597 0 0.0 1e-06 
3.0 3.597 0 0.0 1e-06 
0.05 3.598 0 0.0 1e-06 
3.0 3.598 0 0.0 1e-06 
0.05 3.599 0 0.0 1e-06 
3.0 3.599 0 0.0 1e-06 
0.05 3.6 0 0.0 1e-06 
3.0 3.6 0 0.0 1e-06 
0.05 3.601 0 0.0 1e-06 
3.0 3.601 0 0.0 1e-06 
0.05 3.602 0 0.0 1e-06 
3.0 3.602 0 0.0 1e-06 
0.05 3.603 0 0.0 1e-06 
3.0 3.603 0 0.0 1e-06 
0.05 3.604 0 0.0 1e-06 
3.0 3.604 0 0.0 1e-06 
0.05 3.605 0 0.0 1e-06 
3.0 3.605 0 0.0 1e-06 
0.05 3.606 0 0.0 1e-06 
3.0 3.606 0 0.0 1e-06 
0.05 3.607 0 0.0 1e-06 
3.0 3.607 0 0.0 1e-06 
0.05 3.608 0 0.0 1e-06 
3.0 3.608 0 0.0 1e-06 
0.05 3.609 0 0.0 1e-06 
3.0 3.609 0 0.0 1e-06 
0.05 3.61 0 0.0 1e-06 
3.0 3.61 0 0.0 1e-06 
0.05 3.611 0 0.0 1e-06 
3.0 3.611 0 0.0 1e-06 
0.05 3.612 0 0.0 1e-06 
3.0 3.612 0 0.0 1e-06 
0.05 3.613 0 0.0 1e-06 
3.0 3.613 0 0.0 1e-06 
0.05 3.614 0 0.0 1e-06 
3.0 3.614 0 0.0 1e-06 
0.05 3.615 0 0.0 1e-06 
3.0 3.615 0 0.0 1e-06 
0.05 3.616 0 0.0 1e-06 
3.0 3.616 0 0.0 1e-06 
0.05 3.617 0 0.0 1e-06 
3.0 3.617 0 0.0 1e-06 
0.05 3.618 0 0.0 1e-06 
3.0 3.618 0 0.0 1e-06 
0.05 3.619 0 0.0 1e-06 
3.0 3.619 0 0.0 1e-06 
0.05 3.62 0 0.0 1e-06 
3.0 3.62 0 0.0 1e-06 
0.05 3.621 0 0.0 1e-06 
3.0 3.621 0 0.0 1e-06 
0.05 3.622 0 0.0 1e-06 
3.0 3.622 0 0.0 1e-06 
0.05 3.623 0 0.0 1e-06 
3.0 3.623 0 0.0 1e-06 
0.05 3.624 0 0.0 1e-06 
3.0 3.624 0 0.0 1e-06 
0.05 3.625 0 0.0 1e-06 
3.0 3.625 0 0.0 1e-06 
0.05 3.626 0 0.0 1e-06 
3.0 3.626 0 0.0 1e-06 
0.05 3.627 0 0.0 1e-06 
3.0 3.627 0 0.0 1e-06 
0.05 3.628 0 0.0 1e-06 
3.0 3.628 0 0.0 1e-06 
0.05 3.629 0 0.0 1e-06 
3.0 3.629 0 0.0 1e-06 
0.05 3.63 0 0.0 1e-06 
3.0 3.63 0 0.0 1e-06 
0.05 3.631 0 0.0 1e-06 
3.0 3.631 0 0.0 1e-06 
0.05 3.632 0 0.0 1e-06 
3.0 3.632 0 0.0 1e-06 
0.05 3.633 0 0.0 1e-06 
3.0 3.633 0 0.0 1e-06 
0.05 3.634 0 0.0 1e-06 
3.0 3.634 0 0.0 1e-06 
0.05 3.635 0 0.0 1e-06 
3.0 3.635 0 0.0 1e-06 
0.05 3.636 0 0.0 1e-06 
3.0 3.636 0 0.0 1e-06 
0.05 3.637 0 0.0 1e-06 
3.0 3.637 0 0.0 1e-06 
0.05 3.638 0 0.0 1e-06 
3.0 3.638 0 0.0 1e-06 
0.05 3.639 0 0.0 1e-06 
3.0 3.639 0 0.0 1e-06 
0.05 3.64 0 0.0 1e-06 
3.0 3.64 0 0.0 1e-06 
0.05 3.641 0 0.0 1e-06 
3.0 3.641 0 0.0 1e-06 
0.05 3.642 0 0.0 1e-06 
3.0 3.642 0 0.0 1e-06 
0.05 3.643 0 0.0 1e-06 
3.0 3.643 0 0.0 1e-06 
0.05 3.644 0 0.0 1e-06 
3.0 3.644 0 0.0 1e-06 
0.05 3.645 0 0.0 1e-06 
3.0 3.645 0 0.0 1e-06 
0.05 3.646 0 0.0 1e-06 
3.0 3.646 0 0.0 1e-06 
0.05 3.647 0 0.0 1e-06 
3.0 3.647 0 0.0 1e-06 
0.05 3.648 0 0.0 1e-06 
3.0 3.648 0 0.0 1e-06 
0.05 3.649 0 0.0 1e-06 
3.0 3.649 0 0.0 1e-06 
0.05 3.65 0 0.0 1e-06 
3.0 3.65 0 0.0 1e-06 
0.05 3.651 0 0.0 1e-06 
3.0 3.651 0 0.0 1e-06 
0.05 3.652 0 0.0 1e-06 
3.0 3.652 0 0.0 1e-06 
0.05 3.653 0 0.0 1e-06 
3.0 3.653 0 0.0 1e-06 
0.05 3.654 0 0.0 1e-06 
3.0 3.654 0 0.0 1e-06 
0.05 3.655 0 0.0 1e-06 
3.0 3.655 0 0.0 1e-06 
0.05 3.656 0 0.0 1e-06 
3.0 3.656 0 0.0 1e-06 
0.05 3.657 0 0.0 1e-06 
3.0 3.657 0 0.0 1e-06 
0.05 3.658 0 0.0 1e-06 
3.0 3.658 0 0.0 1e-06 
0.05 3.659 0 0.0 1e-06 
3.0 3.659 0 0.0 1e-06 
0.05 3.66 0 0.0 1e-06 
3.0 3.66 0 0.0 1e-06 
0.05 3.661 0 0.0 1e-06 
3.0 3.661 0 0.0 1e-06 
0.05 3.662 0 0.0 1e-06 
3.0 3.662 0 0.0 1e-06 
0.05 3.663 0 0.0 1e-06 
3.0 3.663 0 0.0 1e-06 
0.05 3.664 0 0.0 1e-06 
3.0 3.664 0 0.0 1e-06 
0.05 3.665 0 0.0 1e-06 
3.0 3.665 0 0.0 1e-06 
0.05 3.666 0 0.0 1e-06 
3.0 3.666 0 0.0 1e-06 
0.05 3.667 0 0.0 1e-06 
3.0 3.667 0 0.0 1e-06 
0.05 3.668 0 0.0 1e-06 
3.0 3.668 0 0.0 1e-06 
0.05 3.669 0 0.0 1e-06 
3.0 3.669 0 0.0 1e-06 
0.05 3.67 0 0.0 1e-06 
3.0 3.67 0 0.0 1e-06 
0.05 3.671 0 0.0 1e-06 
3.0 3.671 0 0.0 1e-06 
0.05 3.672 0 0.0 1e-06 
3.0 3.672 0 0.0 1e-06 
0.05 3.673 0 0.0 1e-06 
3.0 3.673 0 0.0 1e-06 
0.05 3.674 0 0.0 1e-06 
3.0 3.674 0 0.0 1e-06 
0.05 3.675 0 0.0 1e-06 
3.0 3.675 0 0.0 1e-06 
0.05 3.676 0 0.0 1e-06 
3.0 3.676 0 0.0 1e-06 
0.05 3.677 0 0.0 1e-06 
3.0 3.677 0 0.0 1e-06 
0.05 3.678 0 0.0 1e-06 
3.0 3.678 0 0.0 1e-06 
0.05 3.679 0 0.0 1e-06 
3.0 3.679 0 0.0 1e-06 
0.05 3.68 0 0.0 1e-06 
3.0 3.68 0 0.0 1e-06 
0.05 3.681 0 0.0 1e-06 
3.0 3.681 0 0.0 1e-06 
0.05 3.682 0 0.0 1e-06 
3.0 3.682 0 0.0 1e-06 
0.05 3.683 0 0.0 1e-06 
3.0 3.683 0 0.0 1e-06 
0.05 3.684 0 0.0 1e-06 
3.0 3.684 0 0.0 1e-06 
0.05 3.685 0 0.0 1e-06 
3.0 3.685 0 0.0 1e-06 
0.05 3.686 0 0.0 1e-06 
3.0 3.686 0 0.0 1e-06 
0.05 3.687 0 0.0 1e-06 
3.0 3.687 0 0.0 1e-06 
0.05 3.688 0 0.0 1e-06 
3.0 3.688 0 0.0 1e-06 
0.05 3.689 0 0.0 1e-06 
3.0 3.689 0 0.0 1e-06 
0.05 3.69 0 0.0 1e-06 
3.0 3.69 0 0.0 1e-06 
0.05 3.691 0 0.0 1e-06 
3.0 3.691 0 0.0 1e-06 
0.05 3.692 0 0.0 1e-06 
3.0 3.692 0 0.0 1e-06 
0.05 3.693 0 0.0 1e-06 
3.0 3.693 0 0.0 1e-06 
0.05 3.694 0 0.0 1e-06 
3.0 3.694 0 0.0 1e-06 
0.05 3.695 0 0.0 1e-06 
3.0 3.695 0 0.0 1e-06 
0.05 3.696 0 0.0 1e-06 
3.0 3.696 0 0.0 1e-06 
0.05 3.697 0 0.0 1e-06 
3.0 3.697 0 0.0 1e-06 
0.05 3.698 0 0.0 1e-06 
3.0 3.698 0 0.0 1e-06 
0.05 3.699 0 0.0 1e-06 
3.0 3.699 0 0.0 1e-06 
0.05 3.7 0 0.0 1e-06 
3.0 3.7 0 0.0 1e-06 
0.05 3.701 0 0.0 1e-06 
3.0 3.701 0 0.0 1e-06 
0.05 3.702 0 0.0 1e-06 
3.0 3.702 0 0.0 1e-06 
0.05 3.703 0 0.0 1e-06 
3.0 3.703 0 0.0 1e-06 
0.05 3.704 0 0.0 1e-06 
3.0 3.704 0 0.0 1e-06 
0.05 3.705 0 0.0 1e-06 
3.0 3.705 0 0.0 1e-06 
0.05 3.706 0 0.0 1e-06 
3.0 3.706 0 0.0 1e-06 
0.05 3.707 0 0.0 1e-06 
3.0 3.707 0 0.0 1e-06 
0.05 3.708 0 0.0 1e-06 
3.0 3.708 0 0.0 1e-06 
0.05 3.709 0 0.0 1e-06 
3.0 3.709 0 0.0 1e-06 
0.05 3.71 0 0.0 1e-06 
3.0 3.71 0 0.0 1e-06 
0.05 3.711 0 0.0 1e-06 
3.0 3.711 0 0.0 1e-06 
0.05 3.712 0 0.0 1e-06 
3.0 3.712 0 0.0 1e-06 
0.05 3.713 0 0.0 1e-06 
3.0 3.713 0 0.0 1e-06 
0.05 3.714 0 0.0 1e-06 
3.0 3.714 0 0.0 1e-06 
0.05 3.715 0 0.0 1e-06 
3.0 3.715 0 0.0 1e-06 
0.05 3.716 0 0.0 1e-06 
3.0 3.716 0 0.0 1e-06 
0.05 3.717 0 0.0 1e-06 
3.0 3.717 0 0.0 1e-06 
0.05 3.718 0 0.0 1e-06 
3.0 3.718 0 0.0 1e-06 
0.05 3.719 0 0.0 1e-06 
3.0 3.719 0 0.0 1e-06 
0.05 3.72 0 0.0 1e-06 
3.0 3.72 0 0.0 1e-06 
0.05 3.721 0 0.0 1e-06 
3.0 3.721 0 0.0 1e-06 
0.05 3.722 0 0.0 1e-06 
3.0 3.722 0 0.0 1e-06 
0.05 3.723 0 0.0 1e-06 
3.0 3.723 0 0.0 1e-06 
0.05 3.724 0 0.0 1e-06 
3.0 3.724 0 0.0 1e-06 
0.05 3.725 0 0.0 1e-06 
3.0 3.725 0 0.0 1e-06 
0.05 3.726 0 0.0 1e-06 
3.0 3.726 0 0.0 1e-06 
0.05 3.727 0 0.0 1e-06 
3.0 3.727 0 0.0 1e-06 
0.05 3.728 0 0.0 1e-06 
3.0 3.728 0 0.0 1e-06 
0.05 3.729 0 0.0 1e-06 
3.0 3.729 0 0.0 1e-06 
0.05 3.73 0 0.0 1e-06 
3.0 3.73 0 0.0 1e-06 
0.05 3.731 0 0.0 1e-06 
3.0 3.731 0 0.0 1e-06 
0.05 3.732 0 0.0 1e-06 
3.0 3.732 0 0.0 1e-06 
0.05 3.733 0 0.0 1e-06 
3.0 3.733 0 0.0 1e-06 
0.05 3.734 0 0.0 1e-06 
3.0 3.734 0 0.0 1e-06 
0.05 3.735 0 0.0 1e-06 
3.0 3.735 0 0.0 1e-06 
0.05 3.736 0 0.0 1e-06 
3.0 3.736 0 0.0 1e-06 
0.05 3.737 0 0.0 1e-06 
3.0 3.737 0 0.0 1e-06 
0.05 3.738 0 0.0 1e-06 
3.0 3.738 0 0.0 1e-06 
0.05 3.739 0 0.0 1e-06 
3.0 3.739 0 0.0 1e-06 
0.05 3.74 0 0.0 1e-06 
3.0 3.74 0 0.0 1e-06 
0.05 3.741 0 0.0 1e-06 
3.0 3.741 0 0.0 1e-06 
0.05 3.742 0 0.0 1e-06 
3.0 3.742 0 0.0 1e-06 
0.05 3.743 0 0.0 1e-06 
3.0 3.743 0 0.0 1e-06 
0.05 3.744 0 0.0 1e-06 
3.0 3.744 0 0.0 1e-06 
0.05 3.745 0 0.0 1e-06 
3.0 3.745 0 0.0 1e-06 
0.05 3.746 0 0.0 1e-06 
3.0 3.746 0 0.0 1e-06 
0.05 3.747 0 0.0 1e-06 
3.0 3.747 0 0.0 1e-06 
0.05 3.748 0 0.0 1e-06 
3.0 3.748 0 0.0 1e-06 
0.05 3.749 0 0.0 1e-06 
3.0 3.749 0 0.0 1e-06 
0.05 3.75 0 0.0 1e-06 
3.0 3.75 0 0.0 1e-06 
0.05 3.751 0 0.0 1e-06 
3.0 3.751 0 0.0 1e-06 
0.05 3.752 0 0.0 1e-06 
3.0 3.752 0 0.0 1e-06 
0.05 3.753 0 0.0 1e-06 
3.0 3.753 0 0.0 1e-06 
0.05 3.754 0 0.0 1e-06 
3.0 3.754 0 0.0 1e-06 
0.05 3.755 0 0.0 1e-06 
3.0 3.755 0 0.0 1e-06 
0.05 3.756 0 0.0 1e-06 
3.0 3.756 0 0.0 1e-06 
0.05 3.757 0 0.0 1e-06 
3.0 3.757 0 0.0 1e-06 
0.05 3.758 0 0.0 1e-06 
3.0 3.758 0 0.0 1e-06 
0.05 3.759 0 0.0 1e-06 
3.0 3.759 0 0.0 1e-06 
0.05 3.76 0 0.0 1e-06 
3.0 3.76 0 0.0 1e-06 
0.05 3.761 0 0.0 1e-06 
3.0 3.761 0 0.0 1e-06 
0.05 3.762 0 0.0 1e-06 
3.0 3.762 0 0.0 1e-06 
0.05 3.763 0 0.0 1e-06 
3.0 3.763 0 0.0 1e-06 
0.05 3.764 0 0.0 1e-06 
3.0 3.764 0 0.0 1e-06 
0.05 3.765 0 0.0 1e-06 
3.0 3.765 0 0.0 1e-06 
0.05 3.766 0 0.0 1e-06 
3.0 3.766 0 0.0 1e-06 
0.05 3.767 0 0.0 1e-06 
3.0 3.767 0 0.0 1e-06 
0.05 3.768 0 0.0 1e-06 
3.0 3.768 0 0.0 1e-06 
0.05 3.769 0 0.0 1e-06 
3.0 3.769 0 0.0 1e-06 
0.05 3.77 0 0.0 1e-06 
3.0 3.77 0 0.0 1e-06 
0.05 3.771 0 0.0 1e-06 
3.0 3.771 0 0.0 1e-06 
0.05 3.772 0 0.0 1e-06 
3.0 3.772 0 0.0 1e-06 
0.05 3.773 0 0.0 1e-06 
3.0 3.773 0 0.0 1e-06 
0.05 3.774 0 0.0 1e-06 
3.0 3.774 0 0.0 1e-06 
0.05 3.775 0 0.0 1e-06 
3.0 3.775 0 0.0 1e-06 
0.05 3.776 0 0.0 1e-06 
3.0 3.776 0 0.0 1e-06 
0.05 3.777 0 0.0 1e-06 
3.0 3.777 0 0.0 1e-06 
0.05 3.778 0 0.0 1e-06 
3.0 3.778 0 0.0 1e-06 
0.05 3.779 0 0.0 1e-06 
3.0 3.779 0 0.0 1e-06 
0.05 3.78 0 0.0 1e-06 
3.0 3.78 0 0.0 1e-06 
0.05 3.781 0 0.0 1e-06 
3.0 3.781 0 0.0 1e-06 
0.05 3.782 0 0.0 1e-06 
3.0 3.782 0 0.0 1e-06 
0.05 3.783 0 0.0 1e-06 
3.0 3.783 0 0.0 1e-06 
0.05 3.784 0 0.0 1e-06 
3.0 3.784 0 0.0 1e-06 
0.05 3.785 0 0.0 1e-06 
3.0 3.785 0 0.0 1e-06 
0.05 3.786 0 0.0 1e-06 
3.0 3.786 0 0.0 1e-06 
0.05 3.787 0 0.0 1e-06 
3.0 3.787 0 0.0 1e-06 
0.05 3.788 0 0.0 1e-06 
3.0 3.788 0 0.0 1e-06 
0.05 3.789 0 0.0 1e-06 
3.0 3.789 0 0.0 1e-06 
0.05 3.79 0 0.0 1e-06 
3.0 3.79 0 0.0 1e-06 
0.05 3.791 0 0.0 1e-06 
3.0 3.791 0 0.0 1e-06 
0.05 3.792 0 0.0 1e-06 
3.0 3.792 0 0.0 1e-06 
0.05 3.793 0 0.0 1e-06 
3.0 3.793 0 0.0 1e-06 
0.05 3.794 0 0.0 1e-06 
3.0 3.794 0 0.0 1e-06 
0.05 3.795 0 0.0 1e-06 
3.0 3.795 0 0.0 1e-06 
0.05 3.796 0 0.0 1e-06 
3.0 3.796 0 0.0 1e-06 
0.05 3.797 0 0.0 1e-06 
3.0 3.797 0 0.0 1e-06 
0.05 3.798 0 0.0 1e-06 
3.0 3.798 0 0.0 1e-06 
0.05 3.799 0 0.0 1e-06 
3.0 3.799 0 0.0 1e-06 
0.05 3.8 0 0.0 1e-06 
3.0 3.8 0 0.0 1e-06 
0.05 3.801 0 0.0 1e-06 
3.0 3.801 0 0.0 1e-06 
0.05 3.802 0 0.0 1e-06 
3.0 3.802 0 0.0 1e-06 
0.05 3.803 0 0.0 1e-06 
3.0 3.803 0 0.0 1e-06 
0.05 3.804 0 0.0 1e-06 
3.0 3.804 0 0.0 1e-06 
0.05 3.805 0 0.0 1e-06 
3.0 3.805 0 0.0 1e-06 
0.05 3.806 0 0.0 1e-06 
3.0 3.806 0 0.0 1e-06 
0.05 3.807 0 0.0 1e-06 
3.0 3.807 0 0.0 1e-06 
0.05 3.808 0 0.0 1e-06 
3.0 3.808 0 0.0 1e-06 
0.05 3.809 0 0.0 1e-06 
3.0 3.809 0 0.0 1e-06 
0.05 3.81 0 0.0 1e-06 
3.0 3.81 0 0.0 1e-06 
0.05 3.811 0 0.0 1e-06 
3.0 3.811 0 0.0 1e-06 
0.05 3.812 0 0.0 1e-06 
3.0 3.812 0 0.0 1e-06 
0.05 3.813 0 0.0 1e-06 
3.0 3.813 0 0.0 1e-06 
0.05 3.814 0 0.0 1e-06 
3.0 3.814 0 0.0 1e-06 
0.05 3.815 0 0.0 1e-06 
3.0 3.815 0 0.0 1e-06 
0.05 3.816 0 0.0 1e-06 
3.0 3.816 0 0.0 1e-06 
0.05 3.817 0 0.0 1e-06 
3.0 3.817 0 0.0 1e-06 
0.05 3.818 0 0.0 1e-06 
3.0 3.818 0 0.0 1e-06 
0.05 3.819 0 0.0 1e-06 
3.0 3.819 0 0.0 1e-06 
0.05 3.82 0 0.0 1e-06 
3.0 3.82 0 0.0 1e-06 
0.05 3.821 0 0.0 1e-06 
3.0 3.821 0 0.0 1e-06 
0.05 3.822 0 0.0 1e-06 
3.0 3.822 0 0.0 1e-06 
0.05 3.823 0 0.0 1e-06 
3.0 3.823 0 0.0 1e-06 
0.05 3.824 0 0.0 1e-06 
3.0 3.824 0 0.0 1e-06 
0.05 3.825 0 0.0 1e-06 
3.0 3.825 0 0.0 1e-06 
0.05 3.826 0 0.0 1e-06 
3.0 3.826 0 0.0 1e-06 
0.05 3.827 0 0.0 1e-06 
3.0 3.827 0 0.0 1e-06 
0.05 3.828 0 0.0 1e-06 
3.0 3.828 0 0.0 1e-06 
0.05 3.829 0 0.0 1e-06 
3.0 3.829 0 0.0 1e-06 
0.05 3.83 0 0.0 1e-06 
3.0 3.83 0 0.0 1e-06 
0.05 3.831 0 0.0 1e-06 
3.0 3.831 0 0.0 1e-06 
0.05 3.832 0 0.0 1e-06 
3.0 3.832 0 0.0 1e-06 
0.05 3.833 0 0.0 1e-06 
3.0 3.833 0 0.0 1e-06 
0.05 3.834 0 0.0 1e-06 
3.0 3.834 0 0.0 1e-06 
0.05 3.835 0 0.0 1e-06 
3.0 3.835 0 0.0 1e-06 
0.05 3.836 0 0.0 1e-06 
3.0 3.836 0 0.0 1e-06 
0.05 3.837 0 0.0 1e-06 
3.0 3.837 0 0.0 1e-06 
0.05 3.838 0 0.0 1e-06 
3.0 3.838 0 0.0 1e-06 
0.05 3.839 0 0.0 1e-06 
3.0 3.839 0 0.0 1e-06 
0.05 3.84 0 0.0 1e-06 
3.0 3.84 0 0.0 1e-06 
0.05 3.841 0 0.0 1e-06 
3.0 3.841 0 0.0 1e-06 
0.05 3.842 0 0.0 1e-06 
3.0 3.842 0 0.0 1e-06 
0.05 3.843 0 0.0 1e-06 
3.0 3.843 0 0.0 1e-06 
0.05 3.844 0 0.0 1e-06 
3.0 3.844 0 0.0 1e-06 
0.05 3.845 0 0.0 1e-06 
3.0 3.845 0 0.0 1e-06 
0.05 3.846 0 0.0 1e-06 
3.0 3.846 0 0.0 1e-06 
0.05 3.847 0 0.0 1e-06 
3.0 3.847 0 0.0 1e-06 
0.05 3.848 0 0.0 1e-06 
3.0 3.848 0 0.0 1e-06 
0.05 3.849 0 0.0 1e-06 
3.0 3.849 0 0.0 1e-06 
0.05 3.85 0 0.0 1e-06 
3.0 3.85 0 0.0 1e-06 
0.05 3.851 0 0.0 1e-06 
3.0 3.851 0 0.0 1e-06 
0.05 3.852 0 0.0 1e-06 
3.0 3.852 0 0.0 1e-06 
0.05 3.853 0 0.0 1e-06 
3.0 3.853 0 0.0 1e-06 
0.05 3.854 0 0.0 1e-06 
3.0 3.854 0 0.0 1e-06 
0.05 3.855 0 0.0 1e-06 
3.0 3.855 0 0.0 1e-06 
0.05 3.856 0 0.0 1e-06 
3.0 3.856 0 0.0 1e-06 
0.05 3.857 0 0.0 1e-06 
3.0 3.857 0 0.0 1e-06 
0.05 3.858 0 0.0 1e-06 
3.0 3.858 0 0.0 1e-06 
0.05 3.859 0 0.0 1e-06 
3.0 3.859 0 0.0 1e-06 
0.05 3.86 0 0.0 1e-06 
3.0 3.86 0 0.0 1e-06 
0.05 3.861 0 0.0 1e-06 
3.0 3.861 0 0.0 1e-06 
0.05 3.862 0 0.0 1e-06 
3.0 3.862 0 0.0 1e-06 
0.05 3.863 0 0.0 1e-06 
3.0 3.863 0 0.0 1e-06 
0.05 3.864 0 0.0 1e-06 
3.0 3.864 0 0.0 1e-06 
0.05 3.865 0 0.0 1e-06 
3.0 3.865 0 0.0 1e-06 
0.05 3.866 0 0.0 1e-06 
3.0 3.866 0 0.0 1e-06 
0.05 3.867 0 0.0 1e-06 
3.0 3.867 0 0.0 1e-06 
0.05 3.868 0 0.0 1e-06 
3.0 3.868 0 0.0 1e-06 
0.05 3.869 0 0.0 1e-06 
3.0 3.869 0 0.0 1e-06 
0.05 3.87 0 0.0 1e-06 
3.0 3.87 0 0.0 1e-06 
0.05 3.871 0 0.0 1e-06 
3.0 3.871 0 0.0 1e-06 
0.05 3.872 0 0.0 1e-06 
3.0 3.872 0 0.0 1e-06 
0.05 3.873 0 0.0 1e-06 
3.0 3.873 0 0.0 1e-06 
0.05 3.874 0 0.0 1e-06 
3.0 3.874 0 0.0 1e-06 
0.05 3.875 0 0.0 1e-06 
3.0 3.875 0 0.0 1e-06 
0.05 3.876 0 0.0 1e-06 
3.0 3.876 0 0.0 1e-06 
0.05 3.877 0 0.0 1e-06 
3.0 3.877 0 0.0 1e-06 
0.05 3.878 0 0.0 1e-06 
3.0 3.878 0 0.0 1e-06 
0.05 3.879 0 0.0 1e-06 
3.0 3.879 0 0.0 1e-06 
0.05 3.88 0 0.0 1e-06 
3.0 3.88 0 0.0 1e-06 
0.05 3.881 0 0.0 1e-06 
3.0 3.881 0 0.0 1e-06 
0.05 3.882 0 0.0 1e-06 
3.0 3.882 0 0.0 1e-06 
0.05 3.883 0 0.0 1e-06 
3.0 3.883 0 0.0 1e-06 
0.05 3.884 0 0.0 1e-06 
3.0 3.884 0 0.0 1e-06 
0.05 3.885 0 0.0 1e-06 
3.0 3.885 0 0.0 1e-06 
0.05 3.886 0 0.0 1e-06 
3.0 3.886 0 0.0 1e-06 
0.05 3.887 0 0.0 1e-06 
3.0 3.887 0 0.0 1e-06 
0.05 3.888 0 0.0 1e-06 
3.0 3.888 0 0.0 1e-06 
0.05 3.889 0 0.0 1e-06 
3.0 3.889 0 0.0 1e-06 
0.05 3.89 0 0.0 1e-06 
3.0 3.89 0 0.0 1e-06 
0.05 3.891 0 0.0 1e-06 
3.0 3.891 0 0.0 1e-06 
0.05 3.892 0 0.0 1e-06 
3.0 3.892 0 0.0 1e-06 
0.05 3.893 0 0.0 1e-06 
3.0 3.893 0 0.0 1e-06 
0.05 3.894 0 0.0 1e-06 
3.0 3.894 0 0.0 1e-06 
0.05 3.895 0 0.0 1e-06 
3.0 3.895 0 0.0 1e-06 
0.05 3.896 0 0.0 1e-06 
3.0 3.896 0 0.0 1e-06 
0.05 3.897 0 0.0 1e-06 
3.0 3.897 0 0.0 1e-06 
0.05 3.898 0 0.0 1e-06 
3.0 3.898 0 0.0 1e-06 
0.05 3.899 0 0.0 1e-06 
3.0 3.899 0 0.0 1e-06 
0.05 3.9 0 0.0 1e-06 
3.0 3.9 0 0.0 1e-06 
0.05 3.901 0 0.0 1e-06 
3.0 3.901 0 0.0 1e-06 
0.05 3.902 0 0.0 1e-06 
3.0 3.902 0 0.0 1e-06 
0.05 3.903 0 0.0 1e-06 
3.0 3.903 0 0.0 1e-06 
0.05 3.904 0 0.0 1e-06 
3.0 3.904 0 0.0 1e-06 
0.05 3.905 0 0.0 1e-06 
3.0 3.905 0 0.0 1e-06 
0.05 3.906 0 0.0 1e-06 
3.0 3.906 0 0.0 1e-06 
0.05 3.907 0 0.0 1e-06 
3.0 3.907 0 0.0 1e-06 
0.05 3.908 0 0.0 1e-06 
3.0 3.908 0 0.0 1e-06 
0.05 3.909 0 0.0 1e-06 
3.0 3.909 0 0.0 1e-06 
0.05 3.91 0 0.0 1e-06 
3.0 3.91 0 0.0 1e-06 
0.05 3.911 0 0.0 1e-06 
3.0 3.911 0 0.0 1e-06 
0.05 3.912 0 0.0 1e-06 
3.0 3.912 0 0.0 1e-06 
0.05 3.913 0 0.0 1e-06 
3.0 3.913 0 0.0 1e-06 
0.05 3.914 0 0.0 1e-06 
3.0 3.914 0 0.0 1e-06 
0.05 3.915 0 0.0 1e-06 
3.0 3.915 0 0.0 1e-06 
0.05 3.916 0 0.0 1e-06 
3.0 3.916 0 0.0 1e-06 
0.05 3.917 0 0.0 1e-06 
3.0 3.917 0 0.0 1e-06 
0.05 3.918 0 0.0 1e-06 
3.0 3.918 0 0.0 1e-06 
0.05 3.919 0 0.0 1e-06 
3.0 3.919 0 0.0 1e-06 
0.05 3.92 0 0.0 1e-06 
3.0 3.92 0 0.0 1e-06 
0.05 3.921 0 0.0 1e-06 
3.0 3.921 0 0.0 1e-06 
0.05 3.922 0 0.0 1e-06 
3.0 3.922 0 0.0 1e-06 
0.05 3.923 0 0.0 1e-06 
3.0 3.923 0 0.0 1e-06 
0.05 3.924 0 0.0 1e-06 
3.0 3.924 0 0.0 1e-06 
0.05 3.925 0 0.0 1e-06 
3.0 3.925 0 0.0 1e-06 
0.05 3.926 0 0.0 1e-06 
3.0 3.926 0 0.0 1e-06 
0.05 3.927 0 0.0 1e-06 
3.0 3.927 0 0.0 1e-06 
0.05 3.928 0 0.0 1e-06 
3.0 3.928 0 0.0 1e-06 
0.05 3.929 0 0.0 1e-06 
3.0 3.929 0 0.0 1e-06 
0.05 3.93 0 0.0 1e-06 
3.0 3.93 0 0.0 1e-06 
0.05 3.931 0 0.0 1e-06 
3.0 3.931 0 0.0 1e-06 
0.05 3.932 0 0.0 1e-06 
3.0 3.932 0 0.0 1e-06 
0.05 3.933 0 0.0 1e-06 
3.0 3.933 0 0.0 1e-06 
0.05 3.934 0 0.0 1e-06 
3.0 3.934 0 0.0 1e-06 
0.05 3.935 0 0.0 1e-06 
3.0 3.935 0 0.0 1e-06 
0.05 3.936 0 0.0 1e-06 
3.0 3.936 0 0.0 1e-06 
0.05 3.937 0 0.0 1e-06 
3.0 3.937 0 0.0 1e-06 
0.05 3.938 0 0.0 1e-06 
3.0 3.938 0 0.0 1e-06 
0.05 3.939 0 0.0 1e-06 
3.0 3.939 0 0.0 1e-06 
0.05 3.94 0 0.0 1e-06 
3.0 3.94 0 0.0 1e-06 
0.05 3.941 0 0.0 1e-06 
3.0 3.941 0 0.0 1e-06 
0.05 3.942 0 0.0 1e-06 
3.0 3.942 0 0.0 1e-06 
0.05 3.943 0 0.0 1e-06 
3.0 3.943 0 0.0 1e-06 
0.05 3.944 0 0.0 1e-06 
3.0 3.944 0 0.0 1e-06 
0.05 3.945 0 0.0 1e-06 
3.0 3.945 0 0.0 1e-06 
0.05 3.946 0 0.0 1e-06 
3.0 3.946 0 0.0 1e-06 
0.05 3.947 0 0.0 1e-06 
3.0 3.947 0 0.0 1e-06 
0.05 3.948 0 0.0 1e-06 
3.0 3.948 0 0.0 1e-06 
0.05 3.949 0 0.0 1e-06 
3.0 3.949 0 0.0 1e-06 
0.05 3.95 0 0.0 1e-06 
3.0 3.95 0 0.0 1e-06 
0.05 3.951 0 0.0 1e-06 
3.0 3.951 0 0.0 1e-06 
0.05 3.952 0 0.0 1e-06 
3.0 3.952 0 0.0 1e-06 
0.05 3.953 0 0.0 1e-06 
3.0 3.953 0 0.0 1e-06 
0.05 3.954 0 0.0 1e-06 
3.0 3.954 0 0.0 1e-06 
0.05 3.955 0 0.0 1e-06 
3.0 3.955 0 0.0 1e-06 
0.05 3.956 0 0.0 1e-06 
3.0 3.956 0 0.0 1e-06 
0.05 3.957 0 0.0 1e-06 
3.0 3.957 0 0.0 1e-06 
0.05 3.958 0 0.0 1e-06 
3.0 3.958 0 0.0 1e-06 
0.05 3.959 0 0.0 1e-06 
3.0 3.959 0 0.0 1e-06 
0.05 3.96 0 0.0 1e-06 
3.0 3.96 0 0.0 1e-06 
0.05 3.961 0 0.0 1e-06 
3.0 3.961 0 0.0 1e-06 
0.05 3.962 0 0.0 1e-06 
3.0 3.962 0 0.0 1e-06 
0.05 3.963 0 0.0 1e-06 
3.0 3.963 0 0.0 1e-06 
0.05 3.964 0 0.0 1e-06 
3.0 3.964 0 0.0 1e-06 
0.05 3.965 0 0.0 1e-06 
3.0 3.965 0 0.0 1e-06 
0.05 3.966 0 0.0 1e-06 
3.0 3.966 0 0.0 1e-06 
0.05 3.967 0 0.0 1e-06 
3.0 3.967 0 0.0 1e-06 
0.05 3.968 0 0.0 1e-06 
3.0 3.968 0 0.0 1e-06 
0.05 3.969 0 0.0 1e-06 
3.0 3.969 0 0.0 1e-06 
0.05 3.97 0 0.0 1e-06 
3.0 3.97 0 0.0 1e-06 
0.05 3.971 0 0.0 1e-06 
3.0 3.971 0 0.0 1e-06 
0.05 3.972 0 0.0 1e-06 
3.0 3.972 0 0.0 1e-06 
0.05 3.973 0 0.0 1e-06 
3.0 3.973 0 0.0 1e-06 
0.05 3.974 0 0.0 1e-06 
3.0 3.974 0 0.0 1e-06 
0.05 3.975 0 0.0 1e-06 
3.0 3.975 0 0.0 1e-06 
0.05 3.976 0 0.0 1e-06 
3.0 3.976 0 0.0 1e-06 
0.05 3.977 0 0.0 1e-06 
3.0 3.977 0 0.0 1e-06 
0.05 3.978 0 0.0 1e-06 
3.0 3.978 0 0.0 1e-06 
0.05 3.979 0 0.0 1e-06 
3.0 3.979 0 0.0 1e-06 
0.05 3.98 0 0.0 1e-06 
3.0 3.98 0 0.0 1e-06 
0.05 3.981 0 0.0 1e-06 
3.0 3.981 0 0.0 1e-06 
0.05 3.982 0 0.0 1e-06 
3.0 3.982 0 0.0 1e-06 
0.05 3.983 0 0.0 1e-06 
3.0 3.983 0 0.0 1e-06 
0.05 3.984 0 0.0 1e-06 
3.0 3.984 0 0.0 1e-06 
0.05 3.985 0 0.0 1e-06 
3.0 3.985 0 0.0 1e-06 
0.05 3.986 0 0.0 1e-06 
3.0 3.986 0 0.0 1e-06 
0.05 3.987 0 0.0 1e-06 
3.0 3.987 0 0.0 1e-06 
0.05 3.988 0 0.0 1e-06 
3.0 3.988 0 0.0 1e-06 
0.05 3.989 0 0.0 1e-06 
3.0 3.989 0 0.0 1e-06 
0.05 3.99 0 0.0 1e-06 
3.0 3.99 0 0.0 1e-06 
0.05 3.991 0 0.0 1e-06 
3.0 3.991 0 0.0 1e-06 
0.05 3.992 0 0.0 1e-06 
3.0 3.992 0 0.0 1e-06 
0.05 3.993 0 0.0 1e-06 
3.0 3.993 0 0.0 1e-06 
0.05 3.994 0 0.0 1e-06 
3.0 3.994 0 0.0 1e-06 
0.05 3.995 0 0.0 1e-06 
3.0 3.995 0 0.0 1e-06 
0.05 3.996 0 0.0 1e-06 
3.0 3.996 0 0.0 1e-06 
0.05 3.997 0 0.0 1e-06 
3.0 3.997 0 0.0 1e-06 
0.05 3.998 0 0.0 1e-06 
3.0 3.998 0 0.0 1e-06 
0.05 3.999 0 0.0 1e-06 
3.0 3.999 0 0.0 1e-06 
0.05 4.0 0 0.0 1e-06 
3.0 4.0 0 0.0 1e-06 
0.05 4.001 0 0.0 1e-06 
3.0 4.001 0 0.0 1e-06 
0.05 4.002 0 0.0 1e-06 
3.0 4.002 0 0.0 1e-06 
0.05 4.003 0 0.0 1e-06 
3.0 4.003 0 0.0 1e-06 
0.05 4.004 0 0.0 1e-06 
3.0 4.004 0 0.0 1e-06 
0.05 4.005 0 0.0 1e-06 
3.0 4.005 0 0.0 1e-06 
0.05 4.006 0 0.0 1e-06 
3.0 4.006 0 0.0 1e-06 
0.05 4.007 0 0.0 1e-06 
3.0 4.007 0 0.0 1e-06 
0.05 4.008 0 0.0 1e-06 
3.0 4.008 0 0.0 1e-06 
0.05 4.009 0 0.0 1e-06 
3.0 4.009 0 0.0 1e-06 
0.05 4.01 0 0.0 1e-06 
3.0 4.01 0 0.0 1e-06 
0.05 4.011 0 0.0 1e-06 
3.0 4.011 0 0.0 1e-06 
0.05 4.012 0 0.0 1e-06 
3.0 4.012 0 0.0 1e-06 
0.05 4.013 0 0.0 1e-06 
3.0 4.013 0 0.0 1e-06 
0.05 4.014 0 0.0 1e-06 
3.0 4.014 0 0.0 1e-06 
0.05 4.015 0 0.0 1e-06 
3.0 4.015 0 0.0 1e-06 
0.05 4.016 0 0.0 1e-06 
3.0 4.016 0 0.0 1e-06 
0.05 4.017 0 0.0 1e-06 
3.0 4.017 0 0.0 1e-06 
0.05 4.018 0 0.0 1e-06 
3.0 4.018 0 0.0 1e-06 
0.05 4.019 0 0.0 1e-06 
3.0 4.019 0 0.0 1e-06 
0.05 4.02 0 0.0 1e-06 
3.0 4.02 0 0.0 1e-06 
0.05 4.021 0 0.0 1e-06 
3.0 4.021 0 0.0 1e-06 
0.05 4.022 0 0.0 1e-06 
3.0 4.022 0 0.0 1e-06 
0.05 4.023 0 0.0 1e-06 
3.0 4.023 0 0.0 1e-06 
0.05 4.024 0 0.0 1e-06 
3.0 4.024 0 0.0 1e-06 
0.05 4.025 0 0.0 1e-06 
3.0 4.025 0 0.0 1e-06 
0.05 4.026 0 0.0 1e-06 
3.0 4.026 0 0.0 1e-06 
0.05 4.027 0 0.0 1e-06 
3.0 4.027 0 0.0 1e-06 
0.05 4.028 0 0.0 1e-06 
3.0 4.028 0 0.0 1e-06 
0.05 4.029 0 0.0 1e-06 
3.0 4.029 0 0.0 1e-06 
0.05 4.03 0 0.0 1e-06 
3.0 4.03 0 0.0 1e-06 
0.05 4.031 0 0.0 1e-06 
3.0 4.031 0 0.0 1e-06 
0.05 4.032 0 0.0 1e-06 
3.0 4.032 0 0.0 1e-06 
0.05 4.033 0 0.0 1e-06 
3.0 4.033 0 0.0 1e-06 
0.05 4.034 0 0.0 1e-06 
3.0 4.034 0 0.0 1e-06 
0.05 4.035 0 0.0 1e-06 
3.0 4.035 0 0.0 1e-06 
0.05 4.036 0 0.0 1e-06 
3.0 4.036 0 0.0 1e-06 
0.05 4.037 0 0.0 1e-06 
3.0 4.037 0 0.0 1e-06 
0.05 4.038 0 0.0 1e-06 
3.0 4.038 0 0.0 1e-06 
0.05 4.039 0 0.0 1e-06 
3.0 4.039 0 0.0 1e-06 
0.05 4.04 0 0.0 1e-06 
3.0 4.04 0 0.0 1e-06 
0.05 4.041 0 0.0 1e-06 
3.0 4.041 0 0.0 1e-06 
0.05 4.042 0 0.0 1e-06 
3.0 4.042 0 0.0 1e-06 
0.05 4.043 0 0.0 1e-06 
3.0 4.043 0 0.0 1e-06 
0.05 4.044 0 0.0 1e-06 
3.0 4.044 0 0.0 1e-06 
0.05 4.045 0 0.0 1e-06 
3.0 4.045 0 0.0 1e-06 
0.05 4.046 0 0.0 1e-06 
3.0 4.046 0 0.0 1e-06 
0.05 4.047 0 0.0 1e-06 
3.0 4.047 0 0.0 1e-06 
0.05 4.048 0 0.0 1e-06 
3.0 4.048 0 0.0 1e-06 
0.05 4.049 0 0.0 1e-06 
3.0 4.049 0 0.0 1e-06 
0.05 4.05 0 0.0 1e-06 
3.0 4.05 0 0.0 1e-06 
0.05 4.051 0 0.0 1e-06 
3.0 4.051 0 0.0 1e-06 
0.05 4.052 0 0.0 1e-06 
3.0 4.052 0 0.0 1e-06 
0.05 4.053 0 0.0 1e-06 
3.0 4.053 0 0.0 1e-06 
0.05 4.054 0 0.0 1e-06 
3.0 4.054 0 0.0 1e-06 
0.05 4.055 0 0.0 1e-06 
3.0 4.055 0 0.0 1e-06 
0.05 4.056 0 0.0 1e-06 
3.0 4.056 0 0.0 1e-06 
0.05 4.057 0 0.0 1e-06 
3.0 4.057 0 0.0 1e-06 
0.05 4.058 0 0.0 1e-06 
3.0 4.058 0 0.0 1e-06 
0.05 4.059 0 0.0 1e-06 
3.0 4.059 0 0.0 1e-06 
0.05 4.06 0 0.0 1e-06 
3.0 4.06 0 0.0 1e-06 
0.05 4.061 0 0.0 1e-06 
3.0 4.061 0 0.0 1e-06 
0.05 4.062 0 0.0 1e-06 
3.0 4.062 0 0.0 1e-06 
0.05 4.063 0 0.0 1e-06 
3.0 4.063 0 0.0 1e-06 
0.05 4.064 0 0.0 1e-06 
3.0 4.064 0 0.0 1e-06 
0.05 4.065 0 0.0 1e-06 
3.0 4.065 0 0.0 1e-06 
0.05 4.066 0 0.0 1e-06 
3.0 4.066 0 0.0 1e-06 
0.05 4.067 0 0.0 1e-06 
3.0 4.067 0 0.0 1e-06 
0.05 4.068 0 0.0 1e-06 
3.0 4.068 0 0.0 1e-06 
0.05 4.069 0 0.0 1e-06 
3.0 4.069 0 0.0 1e-06 
0.05 4.07 0 0.0 1e-06 
3.0 4.07 0 0.0 1e-06 
0.05 4.071 0 0.0 1e-06 
3.0 4.071 0 0.0 1e-06 
0.05 4.072 0 0.0 1e-06 
3.0 4.072 0 0.0 1e-06 
0.05 4.073 0 0.0 1e-06 
3.0 4.073 0 0.0 1e-06 
0.05 4.074 0 0.0 1e-06 
3.0 4.074 0 0.0 1e-06 
0.05 4.075 0 0.0 1e-06 
3.0 4.075 0 0.0 1e-06 
0.05 4.076 0 0.0 1e-06 
3.0 4.076 0 0.0 1e-06 
0.05 4.077 0 0.0 1e-06 
3.0 4.077 0 0.0 1e-06 
0.05 4.078 0 0.0 1e-06 
3.0 4.078 0 0.0 1e-06 
0.05 4.079 0 0.0 1e-06 
3.0 4.079 0 0.0 1e-06 
0.05 4.08 0 0.0 1e-06 
3.0 4.08 0 0.0 1e-06 
0.05 4.081 0 0.0 1e-06 
3.0 4.081 0 0.0 1e-06 
0.05 4.082 0 0.0 1e-06 
3.0 4.082 0 0.0 1e-06 
0.05 4.083 0 0.0 1e-06 
3.0 4.083 0 0.0 1e-06 
0.05 4.084 0 0.0 1e-06 
3.0 4.084 0 0.0 1e-06 
0.05 4.085 0 0.0 1e-06 
3.0 4.085 0 0.0 1e-06 
0.05 4.086 0 0.0 1e-06 
3.0 4.086 0 0.0 1e-06 
0.05 4.087 0 0.0 1e-06 
3.0 4.087 0 0.0 1e-06 
0.05 4.088 0 0.0 1e-06 
3.0 4.088 0 0.0 1e-06 
0.05 4.089 0 0.0 1e-06 
3.0 4.089 0 0.0 1e-06 
0.05 4.09 0 0.0 1e-06 
3.0 4.09 0 0.0 1e-06 
0.05 4.091 0 0.0 1e-06 
3.0 4.091 0 0.0 1e-06 
0.05 4.092 0 0.0 1e-06 
3.0 4.092 0 0.0 1e-06 
0.05 4.093 0 0.0 1e-06 
3.0 4.093 0 0.0 1e-06 
0.05 4.094 0 0.0 1e-06 
3.0 4.094 0 0.0 1e-06 
0.05 4.095 0 0.0 1e-06 
3.0 4.095 0 0.0 1e-06 
0.05 4.096 0 0.0 1e-06 
3.0 4.096 0 0.0 1e-06 
0.05 4.097 0 0.0 1e-06 
3.0 4.097 0 0.0 1e-06 
0.05 4.098 0 0.0 1e-06 
3.0 4.098 0 0.0 1e-06 
0.05 4.099 0 0.0 1e-06 
3.0 4.099 0 0.0 1e-06 
0.05 4.1 0 0.0 1e-06 
3.0 4.1 0 0.0 1e-06 
0.05 4.101 0 0.0 1e-06 
3.0 4.101 0 0.0 1e-06 
0.05 4.102 0 0.0 1e-06 
3.0 4.102 0 0.0 1e-06 
0.05 4.103 0 0.0 1e-06 
3.0 4.103 0 0.0 1e-06 
0.05 4.104 0 0.0 1e-06 
3.0 4.104 0 0.0 1e-06 
0.05 4.105 0 0.0 1e-06 
3.0 4.105 0 0.0 1e-06 
0.05 4.106 0 0.0 1e-06 
3.0 4.106 0 0.0 1e-06 
0.05 4.107 0 0.0 1e-06 
3.0 4.107 0 0.0 1e-06 
0.05 4.108 0 0.0 1e-06 
3.0 4.108 0 0.0 1e-06 
0.05 4.109 0 0.0 1e-06 
3.0 4.109 0 0.0 1e-06 
0.05 4.11 0 0.0 1e-06 
3.0 4.11 0 0.0 1e-06 
0.05 4.111 0 0.0 1e-06 
3.0 4.111 0 0.0 1e-06 
0.05 4.112 0 0.0 1e-06 
3.0 4.112 0 0.0 1e-06 
0.05 4.113 0 0.0 1e-06 
3.0 4.113 0 0.0 1e-06 
0.05 4.114 0 0.0 1e-06 
3.0 4.114 0 0.0 1e-06 
0.05 4.115 0 0.0 1e-06 
3.0 4.115 0 0.0 1e-06 
0.05 4.116 0 0.0 1e-06 
3.0 4.116 0 0.0 1e-06 
0.05 4.117 0 0.0 1e-06 
3.0 4.117 0 0.0 1e-06 
0.05 4.118 0 0.0 1e-06 
3.0 4.118 0 0.0 1e-06 
0.05 4.119 0 0.0 1e-06 
3.0 4.119 0 0.0 1e-06 
0.05 4.12 0 0.0 1e-06 
3.0 4.12 0 0.0 1e-06 
0.05 4.121 0 0.0 1e-06 
3.0 4.121 0 0.0 1e-06 
0.05 4.122 0 0.0 1e-06 
3.0 4.122 0 0.0 1e-06 
0.05 4.123 0 0.0 1e-06 
3.0 4.123 0 0.0 1e-06 
0.05 4.124 0 0.0 1e-06 
3.0 4.124 0 0.0 1e-06 
0.05 4.125 0 0.0 1e-06 
3.0 4.125 0 0.0 1e-06 
0.05 4.126 0 0.0 1e-06 
3.0 4.126 0 0.0 1e-06 
0.05 4.127 0 0.0 1e-06 
3.0 4.127 0 0.0 1e-06 
0.05 4.128 0 0.0 1e-06 
3.0 4.128 0 0.0 1e-06 
0.05 4.129 0 0.0 1e-06 
3.0 4.129 0 0.0 1e-06 
0.05 4.13 0 0.0 1e-06 
3.0 4.13 0 0.0 1e-06 
0.05 4.131 0 0.0 1e-06 
3.0 4.131 0 0.0 1e-06 
0.05 4.132 0 0.0 1e-06 
3.0 4.132 0 0.0 1e-06 
0.05 4.133 0 0.0 1e-06 
3.0 4.133 0 0.0 1e-06 
0.05 4.134 0 0.0 1e-06 
3.0 4.134 0 0.0 1e-06 
0.05 4.135 0 0.0 1e-06 
3.0 4.135 0 0.0 1e-06 
0.05 4.136 0 0.0 1e-06 
3.0 4.136 0 0.0 1e-06 
0.05 4.137 0 0.0 1e-06 
3.0 4.137 0 0.0 1e-06 
0.05 4.138 0 0.0 1e-06 
3.0 4.138 0 0.0 1e-06 
0.05 4.139 0 0.0 1e-06 
3.0 4.139 0 0.0 1e-06 
0.05 4.14 0 0.0 1e-06 
3.0 4.14 0 0.0 1e-06 
0.05 4.141 0 0.0 1e-06 
3.0 4.141 0 0.0 1e-06 
0.05 4.142 0 0.0 1e-06 
3.0 4.142 0 0.0 1e-06 
0.05 4.143 0 0.0 1e-06 
3.0 4.143 0 0.0 1e-06 
0.05 4.144 0 0.0 1e-06 
3.0 4.144 0 0.0 1e-06 
0.05 4.145 0 0.0 1e-06 
3.0 4.145 0 0.0 1e-06 
0.05 4.146 0 0.0 1e-06 
3.0 4.146 0 0.0 1e-06 
0.05 4.147 0 0.0 1e-06 
3.0 4.147 0 0.0 1e-06 
0.05 4.148 0 0.0 1e-06 
3.0 4.148 0 0.0 1e-06 
0.05 4.149 0 0.0 1e-06 
3.0 4.149 0 0.0 1e-06 
0.05 4.15 0 0.0 1e-06 
3.0 4.15 0 0.0 1e-06 
0.05 4.151 0 0.0 1e-06 
3.0 4.151 0 0.0 1e-06 
0.05 4.152 0 0.0 1e-06 
3.0 4.152 0 0.0 1e-06 
0.05 4.153 0 0.0 1e-06 
3.0 4.153 0 0.0 1e-06 
0.05 4.154 0 0.0 1e-06 
3.0 4.154 0 0.0 1e-06 
0.05 4.155 0 0.0 1e-06 
3.0 4.155 0 0.0 1e-06 
0.05 4.156 0 0.0 1e-06 
3.0 4.156 0 0.0 1e-06 
0.05 4.157 0 0.0 1e-06 
3.0 4.157 0 0.0 1e-06 
0.05 4.158 0 0.0 1e-06 
3.0 4.158 0 0.0 1e-06 
0.05 4.159 0 0.0 1e-06 
3.0 4.159 0 0.0 1e-06 
0.05 4.16 0 0.0 1e-06 
3.0 4.16 0 0.0 1e-06 
0.05 4.161 0 0.0 1e-06 
3.0 4.161 0 0.0 1e-06 
0.05 4.162 0 0.0 1e-06 
3.0 4.162 0 0.0 1e-06 
0.05 4.163 0 0.0 1e-06 
3.0 4.163 0 0.0 1e-06 
0.05 4.164 0 0.0 1e-06 
3.0 4.164 0 0.0 1e-06 
0.05 4.165 0 0.0 1e-06 
3.0 4.165 0 0.0 1e-06 
0.05 4.166 0 0.0 1e-06 
3.0 4.166 0 0.0 1e-06 
0.05 4.167 0 0.0 1e-06 
3.0 4.167 0 0.0 1e-06 
0.05 4.168 0 0.0 1e-06 
3.0 4.168 0 0.0 1e-06 
0.05 4.169 0 0.0 1e-06 
3.0 4.169 0 0.0 1e-06 
0.05 4.17 0 0.0 1e-06 
3.0 4.17 0 0.0 1e-06 
0.05 4.171 0 0.0 1e-06 
3.0 4.171 0 0.0 1e-06 
0.05 4.172 0 0.0 1e-06 
3.0 4.172 0 0.0 1e-06 
0.05 4.173 0 0.0 1e-06 
3.0 4.173 0 0.0 1e-06 
0.05 4.174 0 0.0 1e-06 
3.0 4.174 0 0.0 1e-06 
0.05 4.175 0 0.0 1e-06 
3.0 4.175 0 0.0 1e-06 
0.05 4.176 0 0.0 1e-06 
3.0 4.176 0 0.0 1e-06 
0.05 4.177 0 0.0 1e-06 
3.0 4.177 0 0.0 1e-06 
0.05 4.178 0 0.0 1e-06 
3.0 4.178 0 0.0 1e-06 
0.05 4.179 0 0.0 1e-06 
3.0 4.179 0 0.0 1e-06 
0.05 4.18 0 0.0 1e-06 
3.0 4.18 0 0.0 1e-06 
0.05 4.181 0 0.0 1e-06 
3.0 4.181 0 0.0 1e-06 
0.05 4.182 0 0.0 1e-06 
3.0 4.182 0 0.0 1e-06 
0.05 4.183 0 0.0 1e-06 
3.0 4.183 0 0.0 1e-06 
0.05 4.184 0 0.0 1e-06 
3.0 4.184 0 0.0 1e-06 
0.05 4.185 0 0.0 1e-06 
3.0 4.185 0 0.0 1e-06 
0.05 4.186 0 0.0 1e-06 
3.0 4.186 0 0.0 1e-06 
0.05 4.187 0 0.0 1e-06 
3.0 4.187 0 0.0 1e-06 
0.05 4.188 0 0.0 1e-06 
3.0 4.188 0 0.0 1e-06 
0.05 4.189 0 0.0 1e-06 
3.0 4.189 0 0.0 1e-06 
0.05 4.19 0 0.0 1e-06 
3.0 4.19 0 0.0 1e-06 
0.05 4.191 0 0.0 1e-06 
3.0 4.191 0 0.0 1e-06 
0.05 4.192 0 0.0 1e-06 
3.0 4.192 0 0.0 1e-06 
0.05 4.193 0 0.0 1e-06 
3.0 4.193 0 0.0 1e-06 
0.05 4.194 0 0.0 1e-06 
3.0 4.194 0 0.0 1e-06 
0.05 4.195 0 0.0 1e-06 
3.0 4.195 0 0.0 1e-06 
0.05 4.196 0 0.0 1e-06 
3.0 4.196 0 0.0 1e-06 
0.05 4.197 0 0.0 1e-06 
3.0 4.197 0 0.0 1e-06 
0.05 4.198 0 0.0 1e-06 
3.0 4.198 0 0.0 1e-06 
0.05 4.199 0 0.0 1e-06 
3.0 4.199 0 0.0 1e-06 
0.05 4.2 0 0.0 1e-06 
3.0 4.2 0 0.0 1e-06 
0.05 4.201 0 0.0 1e-06 
3.0 4.201 0 0.0 1e-06 
0.05 4.202 0 0.0 1e-06 
3.0 4.202 0 0.0 1e-06 
0.05 4.203 0 0.0 1e-06 
3.0 4.203 0 0.0 1e-06 
0.05 4.204 0 0.0 1e-06 
3.0 4.204 0 0.0 1e-06 
0.05 4.205 0 0.0 1e-06 
3.0 4.205 0 0.0 1e-06 
0.05 4.206 0 0.0 1e-06 
3.0 4.206 0 0.0 1e-06 
0.05 4.207 0 0.0 1e-06 
3.0 4.207 0 0.0 1e-06 
0.05 4.208 0 0.0 1e-06 
3.0 4.208 0 0.0 1e-06 
0.05 4.209 0 0.0 1e-06 
3.0 4.209 0 0.0 1e-06 
0.05 4.21 0 0.0 1e-06 
3.0 4.21 0 0.0 1e-06 
0.05 4.211 0 0.0 1e-06 
3.0 4.211 0 0.0 1e-06 
0.05 4.212 0 0.0 1e-06 
3.0 4.212 0 0.0 1e-06 
0.05 4.213 0 0.0 1e-06 
3.0 4.213 0 0.0 1e-06 
0.05 4.214 0 0.0 1e-06 
3.0 4.214 0 0.0 1e-06 
0.05 4.215 0 0.0 1e-06 
3.0 4.215 0 0.0 1e-06 
0.05 4.216 0 0.0 1e-06 
3.0 4.216 0 0.0 1e-06 
0.05 4.217 0 0.0 1e-06 
3.0 4.217 0 0.0 1e-06 
0.05 4.218 0 0.0 1e-06 
3.0 4.218 0 0.0 1e-06 
0.05 4.219 0 0.0 1e-06 
3.0 4.219 0 0.0 1e-06 
0.05 4.22 0 0.0 1e-06 
3.0 4.22 0 0.0 1e-06 
0.05 4.221 0 0.0 1e-06 
3.0 4.221 0 0.0 1e-06 
0.05 4.222 0 0.0 1e-06 
3.0 4.222 0 0.0 1e-06 
0.05 4.223 0 0.0 1e-06 
3.0 4.223 0 0.0 1e-06 
0.05 4.224 0 0.0 1e-06 
3.0 4.224 0 0.0 1e-06 
0.05 4.225 0 0.0 1e-06 
3.0 4.225 0 0.0 1e-06 
0.05 4.226 0 0.0 1e-06 
3.0 4.226 0 0.0 1e-06 
0.05 4.227 0 0.0 1e-06 
3.0 4.227 0 0.0 1e-06 
0.05 4.228 0 0.0 1e-06 
3.0 4.228 0 0.0 1e-06 
0.05 4.229 0 0.0 1e-06 
3.0 4.229 0 0.0 1e-06 
0.05 4.23 0 0.0 1e-06 
3.0 4.23 0 0.0 1e-06 
0.05 4.231 0 0.0 1e-06 
3.0 4.231 0 0.0 1e-06 
0.05 4.232 0 0.0 1e-06 
3.0 4.232 0 0.0 1e-06 
0.05 4.233 0 0.0 1e-06 
3.0 4.233 0 0.0 1e-06 
0.05 4.234 0 0.0 1e-06 
3.0 4.234 0 0.0 1e-06 
0.05 4.235 0 0.0 1e-06 
3.0 4.235 0 0.0 1e-06 
0.05 4.236 0 0.0 1e-06 
3.0 4.236 0 0.0 1e-06 
0.05 4.237 0 0.0 1e-06 
3.0 4.237 0 0.0 1e-06 
0.05 4.238 0 0.0 1e-06 
3.0 4.238 0 0.0 1e-06 
0.05 4.239 0 0.0 1e-06 
3.0 4.239 0 0.0 1e-06 
0.05 4.24 0 0.0 1e-06 
3.0 4.24 0 0.0 1e-06 
0.05 4.241 0 0.0 1e-06 
3.0 4.241 0 0.0 1e-06 
0.05 4.242 0 0.0 1e-06 
3.0 4.242 0 0.0 1e-06 
0.05 4.243 0 0.0 1e-06 
3.0 4.243 0 0.0 1e-06 
0.05 4.244 0 0.0 1e-06 
3.0 4.244 0 0.0 1e-06 
0.05 4.245 0 0.0 1e-06 
3.0 4.245 0 0.0 1e-06 
0.05 4.246 0 0.0 1e-06 
3.0 4.246 0 0.0 1e-06 
0.05 4.247 0 0.0 1e-06 
3.0 4.247 0 0.0 1e-06 
0.05 4.248 0 0.0 1e-06 
3.0 4.248 0 0.0 1e-06 
0.05 4.249 0 0.0 1e-06 
3.0 4.249 0 0.0 1e-06 
0.05 4.25 0 0.0 1e-06 
3.0 4.25 0 0.0 1e-06 
0.05 4.251 0 0.0 1e-06 
3.0 4.251 0 0.0 1e-06 
0.05 4.252 0 0.0 1e-06 
3.0 4.252 0 0.0 1e-06 
0.05 4.253 0 0.0 1e-06 
3.0 4.253 0 0.0 1e-06 
0.05 4.254 0 0.0 1e-06 
3.0 4.254 0 0.0 1e-06 
0.05 4.255 0 0.0 1e-06 
3.0 4.255 0 0.0 1e-06 
0.05 4.256 0 0.0 1e-06 
3.0 4.256 0 0.0 1e-06 
0.05 4.257 0 0.0 1e-06 
3.0 4.257 0 0.0 1e-06 
0.05 4.258 0 0.0 1e-06 
3.0 4.258 0 0.0 1e-06 
0.05 4.259 0 0.0 1e-06 
3.0 4.259 0 0.0 1e-06 
0.05 4.26 0 0.0 1e-06 
3.0 4.26 0 0.0 1e-06 
0.05 4.261 0 0.0 1e-06 
3.0 4.261 0 0.0 1e-06 
0.05 4.262 0 0.0 1e-06 
3.0 4.262 0 0.0 1e-06 
0.05 4.263 0 0.0 1e-06 
3.0 4.263 0 0.0 1e-06 
0.05 4.264 0 0.0 1e-06 
3.0 4.264 0 0.0 1e-06 
0.05 4.265 0 0.0 1e-06 
3.0 4.265 0 0.0 1e-06 
0.05 4.266 0 0.0 1e-06 
3.0 4.266 0 0.0 1e-06 
0.05 4.267 0 0.0 1e-06 
3.0 4.267 0 0.0 1e-06 
0.05 4.268 0 0.0 1e-06 
3.0 4.268 0 0.0 1e-06 
0.05 4.269 0 0.0 1e-06 
3.0 4.269 0 0.0 1e-06 
0.05 4.27 0 0.0 1e-06 
3.0 4.27 0 0.0 1e-06 
0.05 4.271 0 0.0 1e-06 
3.0 4.271 0 0.0 1e-06 
0.05 4.272 0 0.0 1e-06 
3.0 4.272 0 0.0 1e-06 
0.05 4.273 0 0.0 1e-06 
3.0 4.273 0 0.0 1e-06 
0.05 4.274 0 0.0 1e-06 
3.0 4.274 0 0.0 1e-06 
0.05 4.275 0 0.0 1e-06 
3.0 4.275 0 0.0 1e-06 
0.05 4.276 0 0.0 1e-06 
3.0 4.276 0 0.0 1e-06 
0.05 4.277 0 0.0 1e-06 
3.0 4.277 0 0.0 1e-06 
0.05 4.278 0 0.0 1e-06 
3.0 4.278 0 0.0 1e-06 
0.05 4.279 0 0.0 1e-06 
3.0 4.279 0 0.0 1e-06 
0.05 4.28 0 0.0 1e-06 
3.0 4.28 0 0.0 1e-06 
0.05 4.281 0 0.0 1e-06 
3.0 4.281 0 0.0 1e-06 
0.05 4.282 0 0.0 1e-06 
3.0 4.282 0 0.0 1e-06 
0.05 4.283 0 0.0 1e-06 
3.0 4.283 0 0.0 1e-06 
0.05 4.284 0 0.0 1e-06 
3.0 4.284 0 0.0 1e-06 
0.05 4.285 0 0.0 1e-06 
3.0 4.285 0 0.0 1e-06 
0.05 4.286 0 0.0 1e-06 
3.0 4.286 0 0.0 1e-06 
0.05 4.287 0 0.0 1e-06 
3.0 4.287 0 0.0 1e-06 
0.05 4.288 0 0.0 1e-06 
3.0 4.288 0 0.0 1e-06 
0.05 4.289 0 0.0 1e-06 
3.0 4.289 0 0.0 1e-06 
0.05 4.29 0 0.0 1e-06 
3.0 4.29 0 0.0 1e-06 
0.05 4.291 0 0.0 1e-06 
3.0 4.291 0 0.0 1e-06 
0.05 4.292 0 0.0 1e-06 
3.0 4.292 0 0.0 1e-06 
0.05 4.293 0 0.0 1e-06 
3.0 4.293 0 0.0 1e-06 
0.05 4.294 0 0.0 1e-06 
3.0 4.294 0 0.0 1e-06 
0.05 4.295 0 0.0 1e-06 
3.0 4.295 0 0.0 1e-06 
0.05 4.296 0 0.0 1e-06 
3.0 4.296 0 0.0 1e-06 
0.05 4.297 0 0.0 1e-06 
3.0 4.297 0 0.0 1e-06 
0.05 4.298 0 0.0 1e-06 
3.0 4.298 0 0.0 1e-06 
0.05 4.299 0 0.0 1e-06 
3.0 4.299 0 0.0 1e-06 
0.05 4.3 0 0.0 1e-06 
3.0 4.3 0 0.0 1e-06 
0.05 4.301 0 0.0 1e-06 
3.0 4.301 0 0.0 1e-06 
0.05 4.302 0 0.0 1e-06 
3.0 4.302 0 0.0 1e-06 
0.05 4.303 0 0.0 1e-06 
3.0 4.303 0 0.0 1e-06 
0.05 4.304 0 0.0 1e-06 
3.0 4.304 0 0.0 1e-06 
0.05 4.305 0 0.0 1e-06 
3.0 4.305 0 0.0 1e-06 
0.05 4.306 0 0.0 1e-06 
3.0 4.306 0 0.0 1e-06 
0.05 4.307 0 0.0 1e-06 
3.0 4.307 0 0.0 1e-06 
0.05 4.308 0 0.0 1e-06 
3.0 4.308 0 0.0 1e-06 
0.05 4.309 0 0.0 1e-06 
3.0 4.309 0 0.0 1e-06 
0.05 4.31 0 0.0 1e-06 
3.0 4.31 0 0.0 1e-06 
0.05 4.311 0 0.0 1e-06 
3.0 4.311 0 0.0 1e-06 
0.05 4.312 0 0.0 1e-06 
3.0 4.312 0 0.0 1e-06 
0.05 4.313 0 0.0 1e-06 
3.0 4.313 0 0.0 1e-06 
0.05 4.314 0 0.0 1e-06 
3.0 4.314 0 0.0 1e-06 
0.05 4.315 0 0.0 1e-06 
3.0 4.315 0 0.0 1e-06 
0.05 4.316 0 0.0 1e-06 
3.0 4.316 0 0.0 1e-06 
0.05 4.317 0 0.0 1e-06 
3.0 4.317 0 0.0 1e-06 
0.05 4.318 0 0.0 1e-06 
3.0 4.318 0 0.0 1e-06 
0.05 4.319 0 0.0 1e-06 
3.0 4.319 0 0.0 1e-06 
0.05 4.32 0 0.0 1e-06 
3.0 4.32 0 0.0 1e-06 
0.05 4.321 0 0.0 1e-06 
3.0 4.321 0 0.0 1e-06 
0.05 4.322 0 0.0 1e-06 
3.0 4.322 0 0.0 1e-06 
0.05 4.323 0 0.0 1e-06 
3.0 4.323 0 0.0 1e-06 
0.05 4.324 0 0.0 1e-06 
3.0 4.324 0 0.0 1e-06 
0.05 4.325 0 0.0 1e-06 
3.0 4.325 0 0.0 1e-06 
0.05 4.326 0 0.0 1e-06 
3.0 4.326 0 0.0 1e-06 
0.05 4.327 0 0.0 1e-06 
3.0 4.327 0 0.0 1e-06 
0.05 4.328 0 0.0 1e-06 
3.0 4.328 0 0.0 1e-06 
0.05 4.329 0 0.0 1e-06 
3.0 4.329 0 0.0 1e-06 
0.05 4.33 0 0.0 1e-06 
3.0 4.33 0 0.0 1e-06 
0.05 4.331 0 0.0 1e-06 
3.0 4.331 0 0.0 1e-06 
0.05 4.332 0 0.0 1e-06 
3.0 4.332 0 0.0 1e-06 
0.05 4.333 0 0.0 1e-06 
3.0 4.333 0 0.0 1e-06 
0.05 4.334 0 0.0 1e-06 
3.0 4.334 0 0.0 1e-06 
0.05 4.335 0 0.0 1e-06 
3.0 4.335 0 0.0 1e-06 
0.05 4.336 0 0.0 1e-06 
3.0 4.336 0 0.0 1e-06 
0.05 4.337 0 0.0 1e-06 
3.0 4.337 0 0.0 1e-06 
0.05 4.338 0 0.0 1e-06 
3.0 4.338 0 0.0 1e-06 
0.05 4.339 0 0.0 1e-06 
3.0 4.339 0 0.0 1e-06 
0.05 4.34 0 0.0 1e-06 
3.0 4.34 0 0.0 1e-06 
0.05 4.341 0 0.0 1e-06 
3.0 4.341 0 0.0 1e-06 
0.05 4.342 0 0.0 1e-06 
3.0 4.342 0 0.0 1e-06 
0.05 4.343 0 0.0 1e-06 
3.0 4.343 0 0.0 1e-06 
0.05 4.344 0 0.0 1e-06 
3.0 4.344 0 0.0 1e-06 
0.05 4.345 0 0.0 1e-06 
3.0 4.345 0 0.0 1e-06 
0.05 4.346 0 0.0 1e-06 
3.0 4.346 0 0.0 1e-06 
0.05 4.347 0 0.0 1e-06 
3.0 4.347 0 0.0 1e-06 
0.05 4.348 0 0.0 1e-06 
3.0 4.348 0 0.0 1e-06 
0.05 4.349 0 0.0 1e-06 
3.0 4.349 0 0.0 1e-06 
0.05 4.35 0 0.0 1e-06 
3.0 4.35 0 0.0 1e-06 
0.05 4.351 0 0.0 1e-06 
3.0 4.351 0 0.0 1e-06 
0.05 4.352 0 0.0 1e-06 
3.0 4.352 0 0.0 1e-06 
0.05 4.353 0 0.0 1e-06 
3.0 4.353 0 0.0 1e-06 
0.05 4.354 0 0.0 1e-06 
3.0 4.354 0 0.0 1e-06 
0.05 4.355 0 0.0 1e-06 
3.0 4.355 0 0.0 1e-06 
0.05 4.356 0 0.0 1e-06 
3.0 4.356 0 0.0 1e-06 
0.05 4.357 0 0.0 1e-06 
3.0 4.357 0 0.0 1e-06 
0.05 4.358 0 0.0 1e-06 
3.0 4.358 0 0.0 1e-06 
0.05 4.359 0 0.0 1e-06 
3.0 4.359 0 0.0 1e-06 
0.05 4.36 0 0.0 1e-06 
3.0 4.36 0 0.0 1e-06 
0.05 4.361 0 0.0 1e-06 
3.0 4.361 0 0.0 1e-06 
0.05 4.362 0 0.0 1e-06 
3.0 4.362 0 0.0 1e-06 
0.05 4.363 0 0.0 1e-06 
3.0 4.363 0 0.0 1e-06 
0.05 4.364 0 0.0 1e-06 
3.0 4.364 0 0.0 1e-06 
0.05 4.365 0 0.0 1e-06 
3.0 4.365 0 0.0 1e-06 
0.05 4.366 0 0.0 1e-06 
3.0 4.366 0 0.0 1e-06 
0.05 4.367 0 0.0 1e-06 
3.0 4.367 0 0.0 1e-06 
0.05 4.368 0 0.0 1e-06 
3.0 4.368 0 0.0 1e-06 
0.05 4.369 0 0.0 1e-06 
3.0 4.369 0 0.0 1e-06 
0.05 4.37 0 0.0 1e-06 
3.0 4.37 0 0.0 1e-06 
0.05 4.371 0 0.0 1e-06 
3.0 4.371 0 0.0 1e-06 
0.05 4.372 0 0.0 1e-06 
3.0 4.372 0 0.0 1e-06 
0.05 4.373 0 0.0 1e-06 
3.0 4.373 0 0.0 1e-06 
0.05 4.374 0 0.0 1e-06 
3.0 4.374 0 0.0 1e-06 
0.05 4.375 0 0.0 1e-06 
3.0 4.375 0 0.0 1e-06 
0.05 4.376 0 0.0 1e-06 
3.0 4.376 0 0.0 1e-06 
0.05 4.377 0 0.0 1e-06 
3.0 4.377 0 0.0 1e-06 
0.05 4.378 0 0.0 1e-06 
3.0 4.378 0 0.0 1e-06 
0.05 4.379 0 0.0 1e-06 
3.0 4.379 0 0.0 1e-06 
0.05 4.38 0 0.0 1e-06 
3.0 4.38 0 0.0 1e-06 
0.05 4.381 0 0.0 1e-06 
3.0 4.381 0 0.0 1e-06 
0.05 4.382 0 0.0 1e-06 
3.0 4.382 0 0.0 1e-06 
0.05 4.383 0 0.0 1e-06 
3.0 4.383 0 0.0 1e-06 
0.05 4.384 0 0.0 1e-06 
3.0 4.384 0 0.0 1e-06 
0.05 4.385 0 0.0 1e-06 
3.0 4.385 0 0.0 1e-06 
0.05 4.386 0 0.0 1e-06 
3.0 4.386 0 0.0 1e-06 
0.05 4.387 0 0.0 1e-06 
3.0 4.387 0 0.0 1e-06 
0.05 4.388 0 0.0 1e-06 
3.0 4.388 0 0.0 1e-06 
0.05 4.389 0 0.0 1e-06 
3.0 4.389 0 0.0 1e-06 
0.05 4.39 0 0.0 1e-06 
3.0 4.39 0 0.0 1e-06 
0.05 4.391 0 0.0 1e-06 
3.0 4.391 0 0.0 1e-06 
0.05 4.392 0 0.0 1e-06 
3.0 4.392 0 0.0 1e-06 
0.05 4.393 0 0.0 1e-06 
3.0 4.393 0 0.0 1e-06 
0.05 4.394 0 0.0 1e-06 
3.0 4.394 0 0.0 1e-06 
0.05 4.395 0 0.0 1e-06 
3.0 4.395 0 0.0 1e-06 
0.05 4.396 0 0.0 1e-06 
3.0 4.396 0 0.0 1e-06 
0.05 4.397 0 0.0 1e-06 
3.0 4.397 0 0.0 1e-06 
0.05 4.398 0 0.0 1e-06 
3.0 4.398 0 0.0 1e-06 
0.05 4.399 0 0.0 1e-06 
3.0 4.399 0 0.0 1e-06 
0.05 4.4 0 0.0 1e-06 
3.0 4.4 0 0.0 1e-06 
0.05 4.401 0 0.0 1e-06 
3.0 4.401 0 0.0 1e-06 
0.05 4.402 0 0.0 1e-06 
3.0 4.402 0 0.0 1e-06 
0.05 4.403 0 0.0 1e-06 
3.0 4.403 0 0.0 1e-06 
0.05 4.404 0 0.0 1e-06 
3.0 4.404 0 0.0 1e-06 
0.05 4.405 0 0.0 1e-06 
3.0 4.405 0 0.0 1e-06 
0.05 4.406 0 0.0 1e-06 
3.0 4.406 0 0.0 1e-06 
0.05 4.407 0 0.0 1e-06 
3.0 4.407 0 0.0 1e-06 
0.05 4.408 0 0.0 1e-06 
3.0 4.408 0 0.0 1e-06 
0.05 4.409 0 0.0 1e-06 
3.0 4.409 0 0.0 1e-06 
0.05 4.41 0 0.0 1e-06 
3.0 4.41 0 0.0 1e-06 
0.05 4.411 0 0.0 1e-06 
3.0 4.411 0 0.0 1e-06 
0.05 4.412 0 0.0 1e-06 
3.0 4.412 0 0.0 1e-06 
0.05 4.413 0 0.0 1e-06 
3.0 4.413 0 0.0 1e-06 
0.05 4.414 0 0.0 1e-06 
3.0 4.414 0 0.0 1e-06 
0.05 4.415 0 0.0 1e-06 
3.0 4.415 0 0.0 1e-06 
0.05 4.416 0 0.0 1e-06 
3.0 4.416 0 0.0 1e-06 
0.05 4.417 0 0.0 1e-06 
3.0 4.417 0 0.0 1e-06 
0.05 4.418 0 0.0 1e-06 
3.0 4.418 0 0.0 1e-06 
0.05 4.419 0 0.0 1e-06 
3.0 4.419 0 0.0 1e-06 
0.05 4.42 0 0.0 1e-06 
3.0 4.42 0 0.0 1e-06 
0.05 4.421 0 0.0 1e-06 
3.0 4.421 0 0.0 1e-06 
0.05 4.422 0 0.0 1e-06 
3.0 4.422 0 0.0 1e-06 
0.05 4.423 0 0.0 1e-06 
3.0 4.423 0 0.0 1e-06 
0.05 4.424 0 0.0 1e-06 
3.0 4.424 0 0.0 1e-06 
0.05 4.425 0 0.0 1e-06 
3.0 4.425 0 0.0 1e-06 
0.05 4.426 0 0.0 1e-06 
3.0 4.426 0 0.0 1e-06 
0.05 4.427 0 0.0 1e-06 
3.0 4.427 0 0.0 1e-06 
0.05 4.428 0 0.0 1e-06 
3.0 4.428 0 0.0 1e-06 
0.05 4.429 0 0.0 1e-06 
3.0 4.429 0 0.0 1e-06 
0.05 4.43 0 0.0 1e-06 
3.0 4.43 0 0.0 1e-06 
0.05 4.431 0 0.0 1e-06 
3.0 4.431 0 0.0 1e-06 
0.05 4.432 0 0.0 1e-06 
3.0 4.432 0 0.0 1e-06 
0.05 4.433 0 0.0 1e-06 
3.0 4.433 0 0.0 1e-06 
0.05 4.434 0 0.0 1e-06 
3.0 4.434 0 0.0 1e-06 
0.05 4.435 0 0.0 1e-06 
3.0 4.435 0 0.0 1e-06 
0.05 4.436 0 0.0 1e-06 
3.0 4.436 0 0.0 1e-06 
0.05 4.437 0 0.0 1e-06 
3.0 4.437 0 0.0 1e-06 
0.05 4.438 0 0.0 1e-06 
3.0 4.438 0 0.0 1e-06 
0.05 4.439 0 0.0 1e-06 
3.0 4.439 0 0.0 1e-06 
0.05 4.44 0 0.0 1e-06 
3.0 4.44 0 0.0 1e-06 
0.05 4.441 0 0.0 1e-06 
3.0 4.441 0 0.0 1e-06 
0.05 4.442 0 0.0 1e-06 
3.0 4.442 0 0.0 1e-06 
0.05 4.443 0 0.0 1e-06 
3.0 4.443 0 0.0 1e-06 
0.05 4.444 0 0.0 1e-06 
3.0 4.444 0 0.0 1e-06 
0.05 4.445 0 0.0 1e-06 
3.0 4.445 0 0.0 1e-06 
0.05 4.446 0 0.0 1e-06 
3.0 4.446 0 0.0 1e-06 
0.05 4.447 0 0.0 1e-06 
3.0 4.447 0 0.0 1e-06 
0.05 4.448 0 0.0 1e-06 
3.0 4.448 0 0.0 1e-06 
0.05 4.449 0 0.0 1e-06 
3.0 4.449 0 0.0 1e-06 
0.05 4.45 0 0.0 1e-06 
3.0 4.45 0 0.0 1e-06 
0.05 4.451 0 0.0 1e-06 
3.0 4.451 0 0.0 1e-06 
0.05 4.452 0 0.0 1e-06 
3.0 4.452 0 0.0 1e-06 
0.05 4.453 0 0.0 1e-06 
3.0 4.453 0 0.0 1e-06 
0.05 4.454 0 0.0 1e-06 
3.0 4.454 0 0.0 1e-06 
0.05 4.455 0 0.0 1e-06 
3.0 4.455 0 0.0 1e-06 
0.05 4.456 0 0.0 1e-06 
3.0 4.456 0 0.0 1e-06 
0.05 4.457 0 0.0 1e-06 
3.0 4.457 0 0.0 1e-06 
0.05 4.458 0 0.0 1e-06 
3.0 4.458 0 0.0 1e-06 
0.05 4.459 0 0.0 1e-06 
3.0 4.459 0 0.0 1e-06 
0.05 4.46 0 0.0 1e-06 
3.0 4.46 0 0.0 1e-06 
0.05 4.461 0 0.0 1e-06 
3.0 4.461 0 0.0 1e-06 
0.05 4.462 0 0.0 1e-06 
3.0 4.462 0 0.0 1e-06 
0.05 4.463 0 0.0 1e-06 
3.0 4.463 0 0.0 1e-06 
0.05 4.464 0 0.0 1e-06 
3.0 4.464 0 0.0 1e-06 
0.05 4.465 0 0.0 1e-06 
3.0 4.465 0 0.0 1e-06 
0.05 4.466 0 0.0 1e-06 
3.0 4.466 0 0.0 1e-06 
0.05 4.467 0 0.0 1e-06 
3.0 4.467 0 0.0 1e-06 
0.05 4.468 0 0.0 1e-06 
3.0 4.468 0 0.0 1e-06 
0.05 4.469 0 0.0 1e-06 
3.0 4.469 0 0.0 1e-06 
0.05 4.47 0 0.0 1e-06 
3.0 4.47 0 0.0 1e-06 
0.05 4.471 0 0.0 1e-06 
3.0 4.471 0 0.0 1e-06 
0.05 4.472 0 0.0 1e-06 
3.0 4.472 0 0.0 1e-06 
0.05 4.473 0 0.0 1e-06 
3.0 4.473 0 0.0 1e-06 
0.05 4.474 0 0.0 1e-06 
3.0 4.474 0 0.0 1e-06 
0.05 4.475 0 0.0 1e-06 
3.0 4.475 0 0.0 1e-06 
0.05 4.476 0 0.0 1e-06 
3.0 4.476 0 0.0 1e-06 
0.05 4.477 0 0.0 1e-06 
3.0 4.477 0 0.0 1e-06 
0.05 4.478 0 0.0 1e-06 
3.0 4.478 0 0.0 1e-06 
0.05 4.479 0 0.0 1e-06 
3.0 4.479 0 0.0 1e-06 
0.05 4.48 0 0.0 1e-06 
3.0 4.48 0 0.0 1e-06 
0.05 4.481 0 0.0 1e-06 
3.0 4.481 0 0.0 1e-06 
0.05 4.482 0 0.0 1e-06 
3.0 4.482 0 0.0 1e-06 
0.05 4.483 0 0.0 1e-06 
3.0 4.483 0 0.0 1e-06 
0.05 4.484 0 0.0 1e-06 
3.0 4.484 0 0.0 1e-06 
0.05 4.485 0 0.0 1e-06 
3.0 4.485 0 0.0 1e-06 
0.05 4.486 0 0.0 1e-06 
3.0 4.486 0 0.0 1e-06 
0.05 4.487 0 0.0 1e-06 
3.0 4.487 0 0.0 1e-06 
0.05 4.488 0 0.0 1e-06 
3.0 4.488 0 0.0 1e-06 
0.05 4.489 0 0.0 1e-06 
3.0 4.489 0 0.0 1e-06 
0.05 4.49 0 0.0 1e-06 
3.0 4.49 0 0.0 1e-06 
0.05 4.491 0 0.0 1e-06 
3.0 4.491 0 0.0 1e-06 
0.05 4.492 0 0.0 1e-06 
3.0 4.492 0 0.0 1e-06 
0.05 4.493 0 0.0 1e-06 
3.0 4.493 0 0.0 1e-06 
0.05 4.494 0 0.0 1e-06 
3.0 4.494 0 0.0 1e-06 
0.05 4.495 0 0.0 1e-06 
3.0 4.495 0 0.0 1e-06 
0.05 4.496 0 0.0 1e-06 
3.0 4.496 0 0.0 1e-06 
0.05 4.497 0 0.0 1e-06 
3.0 4.497 0 0.0 1e-06 
0.05 4.498 0 0.0 1e-06 
3.0 4.498 0 0.0 1e-06 
0.05 4.499 0 0.0 1e-06 
3.0 4.499 0 0.0 1e-06 
0.05 4.5 0 0.0 1e-06 
3.0 4.5 0 0.0 1e-06 
0.05 4.501 0 0.0 1e-06 
3.0 4.501 0 0.0 1e-06 
0.05 4.502 0 0.0 1e-06 
3.0 4.502 0 0.0 1e-06 
0.05 4.503 0 0.0 1e-06 
3.0 4.503 0 0.0 1e-06 
0.05 4.504 0 0.0 1e-06 
3.0 4.504 0 0.0 1e-06 
0.05 4.505 0 0.0 1e-06 
3.0 4.505 0 0.0 1e-06 
0.05 4.506 0 0.0 1e-06 
3.0 4.506 0 0.0 1e-06 
0.05 4.507 0 0.0 1e-06 
3.0 4.507 0 0.0 1e-06 
0.05 4.508 0 0.0 1e-06 
3.0 4.508 0 0.0 1e-06 
0.05 4.509 0 0.0 1e-06 
3.0 4.509 0 0.0 1e-06 
0.05 4.51 0 0.0 1e-06 
3.0 4.51 0 0.0 1e-06 
0.05 4.511 0 0.0 1e-06 
3.0 4.511 0 0.0 1e-06 
0.05 4.512 0 0.0 1e-06 
3.0 4.512 0 0.0 1e-06 
0.05 4.513 0 0.0 1e-06 
3.0 4.513 0 0.0 1e-06 
0.05 4.514 0 0.0 1e-06 
3.0 4.514 0 0.0 1e-06 
0.05 4.515 0 0.0 1e-06 
3.0 4.515 0 0.0 1e-06 
0.05 4.516 0 0.0 1e-06 
3.0 4.516 0 0.0 1e-06 
0.05 4.517 0 0.0 1e-06 
3.0 4.517 0 0.0 1e-06 
0.05 4.518 0 0.0 1e-06 
3.0 4.518 0 0.0 1e-06 
0.05 4.519 0 0.0 1e-06 
3.0 4.519 0 0.0 1e-06 
0.05 4.52 0 0.0 1e-06 
3.0 4.52 0 0.0 1e-06 
0.05 4.521 0 0.0 1e-06 
3.0 4.521 0 0.0 1e-06 
0.05 4.522 0 0.0 1e-06 
3.0 4.522 0 0.0 1e-06 
0.05 4.523 0 0.0 1e-06 
3.0 4.523 0 0.0 1e-06 
0.05 4.524 0 0.0 1e-06 
3.0 4.524 0 0.0 1e-06 
0.05 4.525 0 0.0 1e-06 
3.0 4.525 0 0.0 1e-06 
0.05 4.526 0 0.0 1e-06 
3.0 4.526 0 0.0 1e-06 
0.05 4.527 0 0.0 1e-06 
3.0 4.527 0 0.0 1e-06 
0.05 4.528 0 0.0 1e-06 
3.0 4.528 0 0.0 1e-06 
0.05 4.529 0 0.0 1e-06 
3.0 4.529 0 0.0 1e-06 
0.05 4.53 0 0.0 1e-06 
3.0 4.53 0 0.0 1e-06 
0.05 4.531 0 0.0 1e-06 
3.0 4.531 0 0.0 1e-06 
0.05 4.532 0 0.0 1e-06 
3.0 4.532 0 0.0 1e-06 
0.05 4.533 0 0.0 1e-06 
3.0 4.533 0 0.0 1e-06 
0.05 4.534 0 0.0 1e-06 
3.0 4.534 0 0.0 1e-06 
0.05 4.535 0 0.0 1e-06 
3.0 4.535 0 0.0 1e-06 
0.05 4.536 0 0.0 1e-06 
3.0 4.536 0 0.0 1e-06 
0.05 4.537 0 0.0 1e-06 
3.0 4.537 0 0.0 1e-06 
0.05 4.538 0 0.0 1e-06 
3.0 4.538 0 0.0 1e-06 
0.05 4.539 0 0.0 1e-06 
3.0 4.539 0 0.0 1e-06 
0.05 4.54 0 0.0 1e-06 
3.0 4.54 0 0.0 1e-06 
0.05 4.541 0 0.0 1e-06 
3.0 4.541 0 0.0 1e-06 
0.05 4.542 0 0.0 1e-06 
3.0 4.542 0 0.0 1e-06 
0.05 4.543 0 0.0 1e-06 
3.0 4.543 0 0.0 1e-06 
0.05 4.544 0 0.0 1e-06 
3.0 4.544 0 0.0 1e-06 
0.05 4.545 0 0.0 1e-06 
3.0 4.545 0 0.0 1e-06 
0.05 4.546 0 0.0 1e-06 
3.0 4.546 0 0.0 1e-06 
0.05 4.547 0 0.0 1e-06 
3.0 4.547 0 0.0 1e-06 
0.05 4.548 0 0.0 1e-06 
3.0 4.548 0 0.0 1e-06 
0.05 4.549 0 0.0 1e-06 
3.0 4.549 0 0.0 1e-06 
0.05 4.55 0 0.0 1e-06 
3.0 4.55 0 0.0 1e-06 
0.05 4.551 0 0.0 1e-06 
3.0 4.551 0 0.0 1e-06 
0.05 4.552 0 0.0 1e-06 
3.0 4.552 0 0.0 1e-06 
0.05 4.553 0 0.0 1e-06 
3.0 4.553 0 0.0 1e-06 
0.05 4.554 0 0.0 1e-06 
3.0 4.554 0 0.0 1e-06 
0.05 4.555 0 0.0 1e-06 
3.0 4.555 0 0.0 1e-06 
0.05 4.556 0 0.0 1e-06 
3.0 4.556 0 0.0 1e-06 
0.05 4.557 0 0.0 1e-06 
3.0 4.557 0 0.0 1e-06 
0.05 4.558 0 0.0 1e-06 
3.0 4.558 0 0.0 1e-06 
0.05 4.559 0 0.0 1e-06 
3.0 4.559 0 0.0 1e-06 
0.05 4.56 0 0.0 1e-06 
3.0 4.56 0 0.0 1e-06 
0.05 4.561 0 0.0 1e-06 
3.0 4.561 0 0.0 1e-06 
0.05 4.562 0 0.0 1e-06 
3.0 4.562 0 0.0 1e-06 
0.05 4.563 0 0.0 1e-06 
3.0 4.563 0 0.0 1e-06 
0.05 4.564 0 0.0 1e-06 
3.0 4.564 0 0.0 1e-06 
0.05 4.565 0 0.0 1e-06 
3.0 4.565 0 0.0 1e-06 
0.05 4.566 0 0.0 1e-06 
3.0 4.566 0 0.0 1e-06 
0.05 4.567 0 0.0 1e-06 
3.0 4.567 0 0.0 1e-06 
0.05 4.568 0 0.0 1e-06 
3.0 4.568 0 0.0 1e-06 
0.05 4.569 0 0.0 1e-06 
3.0 4.569 0 0.0 1e-06 
0.05 4.57 0 0.0 1e-06 
3.0 4.57 0 0.0 1e-06 
0.05 4.571 0 0.0 1e-06 
3.0 4.571 0 0.0 1e-06 
0.05 4.572 0 0.0 1e-06 
3.0 4.572 0 0.0 1e-06 
0.05 4.573 0 0.0 1e-06 
3.0 4.573 0 0.0 1e-06 
0.05 4.574 0 0.0 1e-06 
3.0 4.574 0 0.0 1e-06 
0.05 4.575 0 0.0 1e-06 
3.0 4.575 0 0.0 1e-06 
0.05 4.576 0 0.0 1e-06 
3.0 4.576 0 0.0 1e-06 
0.05 4.577 0 0.0 1e-06 
3.0 4.577 0 0.0 1e-06 
0.05 4.578 0 0.0 1e-06 
3.0 4.578 0 0.0 1e-06 
0.05 4.579 0 0.0 1e-06 
3.0 4.579 0 0.0 1e-06 
0.05 4.58 0 0.0 1e-06 
3.0 4.58 0 0.0 1e-06 
0.05 4.581 0 0.0 1e-06 
3.0 4.581 0 0.0 1e-06 
0.05 4.582 0 0.0 1e-06 
3.0 4.582 0 0.0 1e-06 
0.05 4.583 0 0.0 1e-06 
3.0 4.583 0 0.0 1e-06 
0.05 4.584 0 0.0 1e-06 
3.0 4.584 0 0.0 1e-06 
0.05 4.585 0 0.0 1e-06 
3.0 4.585 0 0.0 1e-06 
0.05 4.586 0 0.0 1e-06 
3.0 4.586 0 0.0 1e-06 
0.05 4.587 0 0.0 1e-06 
3.0 4.587 0 0.0 1e-06 
0.05 4.588 0 0.0 1e-06 
3.0 4.588 0 0.0 1e-06 
0.05 4.589 0 0.0 1e-06 
3.0 4.589 0 0.0 1e-06 
0.05 4.59 0 0.0 1e-06 
3.0 4.59 0 0.0 1e-06 
0.05 4.591 0 0.0 1e-06 
3.0 4.591 0 0.0 1e-06 
0.05 4.592 0 0.0 1e-06 
3.0 4.592 0 0.0 1e-06 
0.05 4.593 0 0.0 1e-06 
3.0 4.593 0 0.0 1e-06 
0.05 4.594 0 0.0 1e-06 
3.0 4.594 0 0.0 1e-06 
0.05 4.595 0 0.0 1e-06 
3.0 4.595 0 0.0 1e-06 
0.05 4.596 0 0.0 1e-06 
3.0 4.596 0 0.0 1e-06 
0.05 4.597 0 0.0 1e-06 
3.0 4.597 0 0.0 1e-06 
0.05 4.598 0 0.0 1e-06 
3.0 4.598 0 0.0 1e-06 
0.05 4.599 0 0.0 1e-06 
3.0 4.599 0 0.0 1e-06 
0.05 4.6 0 0.0 1e-06 
3.0 4.6 0 0.0 1e-06 
0.05 4.601 0 0.0 1e-06 
3.0 4.601 0 0.0 1e-06 
0.05 4.602 0 0.0 1e-06 
3.0 4.602 0 0.0 1e-06 
0.05 4.603 0 0.0 1e-06 
3.0 4.603 0 0.0 1e-06 
0.05 4.604 0 0.0 1e-06 
3.0 4.604 0 0.0 1e-06 
0.05 4.605 0 0.0 1e-06 
3.0 4.605 0 0.0 1e-06 
0.05 4.606 0 0.0 1e-06 
3.0 4.606 0 0.0 1e-06 
0.05 4.607 0 0.0 1e-06 
3.0 4.607 0 0.0 1e-06 
0.05 4.608 0 0.0 1e-06 
3.0 4.608 0 0.0 1e-06 
0.05 4.609 0 0.0 1e-06 
3.0 4.609 0 0.0 1e-06 
0.05 4.61 0 0.0 1e-06 
3.0 4.61 0 0.0 1e-06 
0.05 4.611 0 0.0 1e-06 
3.0 4.611 0 0.0 1e-06 
0.05 4.612 0 0.0 1e-06 
3.0 4.612 0 0.0 1e-06 
0.05 4.613 0 0.0 1e-06 
3.0 4.613 0 0.0 1e-06 
0.05 4.614 0 0.0 1e-06 
3.0 4.614 0 0.0 1e-06 
0.05 4.615 0 0.0 1e-06 
3.0 4.615 0 0.0 1e-06 
0.05 4.616 0 0.0 1e-06 
3.0 4.616 0 0.0 1e-06 
0.05 4.617 0 0.0 1e-06 
3.0 4.617 0 0.0 1e-06 
0.05 4.618 0 0.0 1e-06 
3.0 4.618 0 0.0 1e-06 
0.05 4.619 0 0.0 1e-06 
3.0 4.619 0 0.0 1e-06 
0.05 4.62 0 0.0 1e-06 
3.0 4.62 0 0.0 1e-06 
0.05 4.621 0 0.0 1e-06 
3.0 4.621 0 0.0 1e-06 
0.05 4.622 0 0.0 1e-06 
3.0 4.622 0 0.0 1e-06 
0.05 4.623 0 0.0 1e-06 
3.0 4.623 0 0.0 1e-06 
0.05 4.624 0 0.0 1e-06 
3.0 4.624 0 0.0 1e-06 
0.05 4.625 0 0.0 1e-06 
3.0 4.625 0 0.0 1e-06 
0.05 4.626 0 0.0 1e-06 
3.0 4.626 0 0.0 1e-06 
0.05 4.627 0 0.0 1e-06 
3.0 4.627 0 0.0 1e-06 
0.05 4.628 0 0.0 1e-06 
3.0 4.628 0 0.0 1e-06 
0.05 4.629 0 0.0 1e-06 
3.0 4.629 0 0.0 1e-06 
0.05 4.63 0 0.0 1e-06 
3.0 4.63 0 0.0 1e-06 
0.05 4.631 0 0.0 1e-06 
3.0 4.631 0 0.0 1e-06 
0.05 4.632 0 0.0 1e-06 
3.0 4.632 0 0.0 1e-06 
0.05 4.633 0 0.0 1e-06 
3.0 4.633 0 0.0 1e-06 
0.05 4.634 0 0.0 1e-06 
3.0 4.634 0 0.0 1e-06 
0.05 4.635 0 0.0 1e-06 
3.0 4.635 0 0.0 1e-06 
0.05 4.636 0 0.0 1e-06 
3.0 4.636 0 0.0 1e-06 
0.05 4.637 0 0.0 1e-06 
3.0 4.637 0 0.0 1e-06 
0.05 4.638 0 0.0 1e-06 
3.0 4.638 0 0.0 1e-06 
0.05 4.639 0 0.0 1e-06 
3.0 4.639 0 0.0 1e-06 
0.05 4.64 0 0.0 1e-06 
3.0 4.64 0 0.0 1e-06 
0.05 4.641 0 0.0 1e-06 
3.0 4.641 0 0.0 1e-06 
0.05 4.642 0 0.0 1e-06 
3.0 4.642 0 0.0 1e-06 
0.05 4.643 0 0.0 1e-06 
3.0 4.643 0 0.0 1e-06 
0.05 4.644 0 0.0 1e-06 
3.0 4.644 0 0.0 1e-06 
0.05 4.645 0 0.0 1e-06 
3.0 4.645 0 0.0 1e-06 
0.05 4.646 0 0.0 1e-06 
3.0 4.646 0 0.0 1e-06 
0.05 4.647 0 0.0 1e-06 
3.0 4.647 0 0.0 1e-06 
0.05 4.648 0 0.0 1e-06 
3.0 4.648 0 0.0 1e-06 
0.05 4.649 0 0.0 1e-06 
3.0 4.649 0 0.0 1e-06 
0.05 4.65 0 0.0 1e-06 
3.0 4.65 0 0.0 1e-06 
0.05 4.651 0 0.0 1e-06 
3.0 4.651 0 0.0 1e-06 
0.05 4.652 0 0.0 1e-06 
3.0 4.652 0 0.0 1e-06 
0.05 4.653 0 0.0 1e-06 
3.0 4.653 0 0.0 1e-06 
0.05 4.654 0 0.0 1e-06 
3.0 4.654 0 0.0 1e-06 
0.05 4.655 0 0.0 1e-06 
3.0 4.655 0 0.0 1e-06 
0.05 4.656 0 0.0 1e-06 
3.0 4.656 0 0.0 1e-06 
0.05 4.657 0 0.0 1e-06 
3.0 4.657 0 0.0 1e-06 
0.05 4.658 0 0.0 1e-06 
3.0 4.658 0 0.0 1e-06 
0.05 4.659 0 0.0 1e-06 
3.0 4.659 0 0.0 1e-06 
0.05 4.66 0 0.0 1e-06 
3.0 4.66 0 0.0 1e-06 
0.05 4.661 0 0.0 1e-06 
3.0 4.661 0 0.0 1e-06 
0.05 4.662 0 0.0 1e-06 
3.0 4.662 0 0.0 1e-06 
0.05 4.663 0 0.0 1e-06 
3.0 4.663 0 0.0 1e-06 
0.05 4.664 0 0.0 1e-06 
3.0 4.664 0 0.0 1e-06 
0.05 4.665 0 0.0 1e-06 
3.0 4.665 0 0.0 1e-06 
0.05 4.666 0 0.0 1e-06 
3.0 4.666 0 0.0 1e-06 
0.05 4.667 0 0.0 1e-06 
3.0 4.667 0 0.0 1e-06 
0.05 4.668 0 0.0 1e-06 
3.0 4.668 0 0.0 1e-06 
0.05 4.669 0 0.0 1e-06 
3.0 4.669 0 0.0 1e-06 
0.05 4.67 0 0.0 1e-06 
3.0 4.67 0 0.0 1e-06 
0.05 4.671 0 0.0 1e-06 
3.0 4.671 0 0.0 1e-06 
0.05 4.672 0 0.0 1e-06 
3.0 4.672 0 0.0 1e-06 
0.05 4.673 0 0.0 1e-06 
3.0 4.673 0 0.0 1e-06 
0.05 4.674 0 0.0 1e-06 
3.0 4.674 0 0.0 1e-06 
0.05 4.675 0 0.0 1e-06 
3.0 4.675 0 0.0 1e-06 
0.05 4.676 0 0.0 1e-06 
3.0 4.676 0 0.0 1e-06 
0.05 4.677 0 0.0 1e-06 
3.0 4.677 0 0.0 1e-06 
0.05 4.678 0 0.0 1e-06 
3.0 4.678 0 0.0 1e-06 
0.05 4.679 0 0.0 1e-06 
3.0 4.679 0 0.0 1e-06 
0.05 4.68 0 0.0 1e-06 
3.0 4.68 0 0.0 1e-06 
0.05 4.681 0 0.0 1e-06 
3.0 4.681 0 0.0 1e-06 
0.05 4.682 0 0.0 1e-06 
3.0 4.682 0 0.0 1e-06 
0.05 4.683 0 0.0 1e-06 
3.0 4.683 0 0.0 1e-06 
0.05 4.684 0 0.0 1e-06 
3.0 4.684 0 0.0 1e-06 
0.05 4.685 0 0.0 1e-06 
3.0 4.685 0 0.0 1e-06 
0.05 4.686 0 0.0 1e-06 
3.0 4.686 0 0.0 1e-06 
0.05 4.687 0 0.0 1e-06 
3.0 4.687 0 0.0 1e-06 
0.05 4.688 0 0.0 1e-06 
3.0 4.688 0 0.0 1e-06 
0.05 4.689 0 0.0 1e-06 
3.0 4.689 0 0.0 1e-06 
0.05 4.69 0 0.0 1e-06 
3.0 4.69 0 0.0 1e-06 
0.05 4.691 0 0.0 1e-06 
3.0 4.691 0 0.0 1e-06 
0.05 4.692 0 0.0 1e-06 
3.0 4.692 0 0.0 1e-06 
0.05 4.693 0 0.0 1e-06 
3.0 4.693 0 0.0 1e-06 
0.05 4.694 0 0.0 1e-06 
3.0 4.694 0 0.0 1e-06 
0.05 4.695 0 0.0 1e-06 
3.0 4.695 0 0.0 1e-06 
0.05 4.696 0 0.0 1e-06 
3.0 4.696 0 0.0 1e-06 
0.05 4.697 0 0.0 1e-06 
3.0 4.697 0 0.0 1e-06 
0.05 4.698 0 0.0 1e-06 
3.0 4.698 0 0.0 1e-06 
0.05 4.699 0 0.0 1e-06 
3.0 4.699 0 0.0 1e-06 
0.05 4.7 0 0.0 1e-06 
3.0 4.7 0 0.0 1e-06 
0.05 4.701 0 0.0 1e-06 
3.0 4.701 0 0.0 1e-06 
0.05 4.702 0 0.0 1e-06 
3.0 4.702 0 0.0 1e-06 
0.05 4.703 0 0.0 1e-06 
3.0 4.703 0 0.0 1e-06 
0.05 4.704 0 0.0 1e-06 
3.0 4.704 0 0.0 1e-06 
0.05 4.705 0 0.0 1e-06 
3.0 4.705 0 0.0 1e-06 
0.05 4.706 0 0.0 1e-06 
3.0 4.706 0 0.0 1e-06 
0.05 4.707 0 0.0 1e-06 
3.0 4.707 0 0.0 1e-06 
0.05 4.708 0 0.0 1e-06 
3.0 4.708 0 0.0 1e-06 
0.05 4.709 0 0.0 1e-06 
3.0 4.709 0 0.0 1e-06 
0.05 4.71 0 0.0 1e-06 
3.0 4.71 0 0.0 1e-06 
0.05 4.711 0 0.0 1e-06 
3.0 4.711 0 0.0 1e-06 
0.05 4.712 0 0.0 1e-06 
3.0 4.712 0 0.0 1e-06 
0.05 4.713 0 0.0 1e-06 
3.0 4.713 0 0.0 1e-06 
0.05 4.714 0 0.0 1e-06 
3.0 4.714 0 0.0 1e-06 
0.05 4.715 0 0.0 1e-06 
3.0 4.715 0 0.0 1e-06 
0.05 4.716 0 0.0 1e-06 
3.0 4.716 0 0.0 1e-06 
0.05 4.717 0 0.0 1e-06 
3.0 4.717 0 0.0 1e-06 
0.05 4.718 0 0.0 1e-06 
3.0 4.718 0 0.0 1e-06 
0.05 4.719 0 0.0 1e-06 
3.0 4.719 0 0.0 1e-06 
0.05 4.72 0 0.0 1e-06 
3.0 4.72 0 0.0 1e-06 
0.05 4.721 0 0.0 1e-06 
3.0 4.721 0 0.0 1e-06 
0.05 4.722 0 0.0 1e-06 
3.0 4.722 0 0.0 1e-06 
0.05 4.723 0 0.0 1e-06 
3.0 4.723 0 0.0 1e-06 
0.05 4.724 0 0.0 1e-06 
3.0 4.724 0 0.0 1e-06 
0.05 4.725 0 0.0 1e-06 
3.0 4.725 0 0.0 1e-06 
0.05 4.726 0 0.0 1e-06 
3.0 4.726 0 0.0 1e-06 
0.05 4.727 0 0.0 1e-06 
3.0 4.727 0 0.0 1e-06 
0.05 4.728 0 0.0 1e-06 
3.0 4.728 0 0.0 1e-06 
0.05 4.729 0 0.0 1e-06 
3.0 4.729 0 0.0 1e-06 
0.05 4.73 0 0.0 1e-06 
3.0 4.73 0 0.0 1e-06 
0.05 4.731 0 0.0 1e-06 
3.0 4.731 0 0.0 1e-06 
0.05 4.732 0 0.0 1e-06 
3.0 4.732 0 0.0 1e-06 
0.05 4.733 0 0.0 1e-06 
3.0 4.733 0 0.0 1e-06 
0.05 4.734 0 0.0 1e-06 
3.0 4.734 0 0.0 1e-06 
0.05 4.735 0 0.0 1e-06 
3.0 4.735 0 0.0 1e-06 
0.05 4.736 0 0.0 1e-06 
3.0 4.736 0 0.0 1e-06 
0.05 4.737 0 0.0 1e-06 
3.0 4.737 0 0.0 1e-06 
0.05 4.738 0 0.0 1e-06 
3.0 4.738 0 0.0 1e-06 
0.05 4.739 0 0.0 1e-06 
3.0 4.739 0 0.0 1e-06 
0.05 4.74 0 0.0 1e-06 
3.0 4.74 0 0.0 1e-06 
0.05 4.741 0 0.0 1e-06 
3.0 4.741 0 0.0 1e-06 
0.05 4.742 0 0.0 1e-06 
3.0 4.742 0 0.0 1e-06 
0.05 4.743 0 0.0 1e-06 
3.0 4.743 0 0.0 1e-06 
0.05 4.744 0 0.0 1e-06 
3.0 4.744 0 0.0 1e-06 
0.05 4.745 0 0.0 1e-06 
3.0 4.745 0 0.0 1e-06 
0.05 4.746 0 0.0 1e-06 
3.0 4.746 0 0.0 1e-06 
0.05 4.747 0 0.0 1e-06 
3.0 4.747 0 0.0 1e-06 
0.05 4.748 0 0.0 1e-06 
3.0 4.748 0 0.0 1e-06 
0.05 4.749 0 0.0 1e-06 
3.0 4.749 0 0.0 1e-06 
0.05 4.75 0 0.0 1e-06 
3.0 4.75 0 0.0 1e-06 
0.05 4.751 0 0.0 1e-06 
3.0 4.751 0 0.0 1e-06 
0.05 4.752 0 0.0 1e-06 
3.0 4.752 0 0.0 1e-06 
0.05 4.753 0 0.0 1e-06 
3.0 4.753 0 0.0 1e-06 
0.05 4.754 0 0.0 1e-06 
3.0 4.754 0 0.0 1e-06 
0.05 4.755 0 0.0 1e-06 
3.0 4.755 0 0.0 1e-06 
0.05 4.756 0 0.0 1e-06 
3.0 4.756 0 0.0 1e-06 
0.05 4.757 0 0.0 1e-06 
3.0 4.757 0 0.0 1e-06 
0.05 4.758 0 0.0 1e-06 
3.0 4.758 0 0.0 1e-06 
0.05 4.759 0 0.0 1e-06 
3.0 4.759 0 0.0 1e-06 
0.05 4.76 0 0.0 1e-06 
3.0 4.76 0 0.0 1e-06 
0.05 4.761 0 0.0 1e-06 
3.0 4.761 0 0.0 1e-06 
0.05 4.762 0 0.0 1e-06 
3.0 4.762 0 0.0 1e-06 
0.05 4.763 0 0.0 1e-06 
3.0 4.763 0 0.0 1e-06 
0.05 4.764 0 0.0 1e-06 
3.0 4.764 0 0.0 1e-06 
0.05 4.765 0 0.0 1e-06 
3.0 4.765 0 0.0 1e-06 
0.05 4.766 0 0.0 1e-06 
3.0 4.766 0 0.0 1e-06 
0.05 4.767 0 0.0 1e-06 
3.0 4.767 0 0.0 1e-06 
0.05 4.768 0 0.0 1e-06 
3.0 4.768 0 0.0 1e-06 
0.05 4.769 0 0.0 1e-06 
3.0 4.769 0 0.0 1e-06 
0.05 4.77 0 0.0 1e-06 
3.0 4.77 0 0.0 1e-06 
0.05 4.771 0 0.0 1e-06 
3.0 4.771 0 0.0 1e-06 
0.05 4.772 0 0.0 1e-06 
3.0 4.772 0 0.0 1e-06 
0.05 4.773 0 0.0 1e-06 
3.0 4.773 0 0.0 1e-06 
0.05 4.774 0 0.0 1e-06 
3.0 4.774 0 0.0 1e-06 
0.05 4.775 0 0.0 1e-06 
3.0 4.775 0 0.0 1e-06 
0.05 4.776 0 0.0 1e-06 
3.0 4.776 0 0.0 1e-06 
0.05 4.777 0 0.0 1e-06 
3.0 4.777 0 0.0 1e-06 
0.05 4.778 0 0.0 1e-06 
3.0 4.778 0 0.0 1e-06 
0.05 4.779 0 0.0 1e-06 
3.0 4.779 0 0.0 1e-06 
0.05 4.78 0 0.0 1e-06 
3.0 4.78 0 0.0 1e-06 
0.05 4.781 0 0.0 1e-06 
3.0 4.781 0 0.0 1e-06 
0.05 4.782 0 0.0 1e-06 
3.0 4.782 0 0.0 1e-06 
0.05 4.783 0 0.0 1e-06 
3.0 4.783 0 0.0 1e-06 
0.05 4.784 0 0.0 1e-06 
3.0 4.784 0 0.0 1e-06 
0.05 4.785 0 0.0 1e-06 
3.0 4.785 0 0.0 1e-06 
0.05 4.786 0 0.0 1e-06 
3.0 4.786 0 0.0 1e-06 
0.05 4.787 0 0.0 1e-06 
3.0 4.787 0 0.0 1e-06 
0.05 4.788 0 0.0 1e-06 
3.0 4.788 0 0.0 1e-06 
0.05 4.789 0 0.0 1e-06 
3.0 4.789 0 0.0 1e-06 
0.05 4.79 0 0.0 1e-06 
3.0 4.79 0 0.0 1e-06 
0.05 4.791 0 0.0 1e-06 
3.0 4.791 0 0.0 1e-06 
0.05 4.792 0 0.0 1e-06 
3.0 4.792 0 0.0 1e-06 
0.05 4.793 0 0.0 1e-06 
3.0 4.793 0 0.0 1e-06 
0.05 4.794 0 0.0 1e-06 
3.0 4.794 0 0.0 1e-06 
0.05 4.795 0 0.0 1e-06 
3.0 4.795 0 0.0 1e-06 
0.05 4.796 0 0.0 1e-06 
3.0 4.796 0 0.0 1e-06 
0.05 4.797 0 0.0 1e-06 
3.0 4.797 0 0.0 1e-06 
0.05 4.798 0 0.0 1e-06 
3.0 4.798 0 0.0 1e-06 
0.05 4.799 0 0.0 1e-06 
3.0 4.799 0 0.0 1e-06 
0.05 4.8 0 0.0 1e-06 
3.0 4.8 0 0.0 1e-06 
0.05 4.801 0 0.0 1e-06 
3.0 4.801 0 0.0 1e-06 
0.05 4.802 0 0.0 1e-06 
3.0 4.802 0 0.0 1e-06 
0.05 4.803 0 0.0 1e-06 
3.0 4.803 0 0.0 1e-06 
0.05 4.804 0 0.0 1e-06 
3.0 4.804 0 0.0 1e-06 
0.05 4.805 0 0.0 1e-06 
3.0 4.805 0 0.0 1e-06 
0.05 4.806 0 0.0 1e-06 
3.0 4.806 0 0.0 1e-06 
0.05 4.807 0 0.0 1e-06 
3.0 4.807 0 0.0 1e-06 
0.05 4.808 0 0.0 1e-06 
3.0 4.808 0 0.0 1e-06 
0.05 4.809 0 0.0 1e-06 
3.0 4.809 0 0.0 1e-06 
0.05 4.81 0 0.0 1e-06 
3.0 4.81 0 0.0 1e-06 
0.05 4.811 0 0.0 1e-06 
3.0 4.811 0 0.0 1e-06 
0.05 4.812 0 0.0 1e-06 
3.0 4.812 0 0.0 1e-06 
0.05 4.813 0 0.0 1e-06 
3.0 4.813 0 0.0 1e-06 
0.05 4.814 0 0.0 1e-06 
3.0 4.814 0 0.0 1e-06 
0.05 4.815 0 0.0 1e-06 
3.0 4.815 0 0.0 1e-06 
0.05 4.816 0 0.0 1e-06 
3.0 4.816 0 0.0 1e-06 
0.05 4.817 0 0.0 1e-06 
3.0 4.817 0 0.0 1e-06 
0.05 4.818 0 0.0 1e-06 
3.0 4.818 0 0.0 1e-06 
0.05 4.819 0 0.0 1e-06 
3.0 4.819 0 0.0 1e-06 
0.05 4.82 0 0.0 1e-06 
3.0 4.82 0 0.0 1e-06 
0.05 4.821 0 0.0 1e-06 
3.0 4.821 0 0.0 1e-06 
0.05 4.822 0 0.0 1e-06 
3.0 4.822 0 0.0 1e-06 
0.05 4.823 0 0.0 1e-06 
3.0 4.823 0 0.0 1e-06 
0.05 4.824 0 0.0 1e-06 
3.0 4.824 0 0.0 1e-06 
0.05 4.825 0 0.0 1e-06 
3.0 4.825 0 0.0 1e-06 
0.05 4.826 0 0.0 1e-06 
3.0 4.826 0 0.0 1e-06 
0.05 4.827 0 0.0 1e-06 
3.0 4.827 0 0.0 1e-06 
0.05 4.828 0 0.0 1e-06 
3.0 4.828 0 0.0 1e-06 
0.05 4.829 0 0.0 1e-06 
3.0 4.829 0 0.0 1e-06 
0.05 4.83 0 0.0 1e-06 
3.0 4.83 0 0.0 1e-06 
0.05 4.831 0 0.0 1e-06 
3.0 4.831 0 0.0 1e-06 
0.05 4.832 0 0.0 1e-06 
3.0 4.832 0 0.0 1e-06 
0.05 4.833 0 0.0 1e-06 
3.0 4.833 0 0.0 1e-06 
0.05 4.834 0 0.0 1e-06 
3.0 4.834 0 0.0 1e-06 
0.05 4.835 0 0.0 1e-06 
3.0 4.835 0 0.0 1e-06 
0.05 4.836 0 0.0 1e-06 
3.0 4.836 0 0.0 1e-06 
0.05 4.837 0 0.0 1e-06 
3.0 4.837 0 0.0 1e-06 
0.05 4.838 0 0.0 1e-06 
3.0 4.838 0 0.0 1e-06 
0.05 4.839 0 0.0 1e-06 
3.0 4.839 0 0.0 1e-06 
0.05 4.84 0 0.0 1e-06 
3.0 4.84 0 0.0 1e-06 
0.05 4.841 0 0.0 1e-06 
3.0 4.841 0 0.0 1e-06 
0.05 4.842 0 0.0 1e-06 
3.0 4.842 0 0.0 1e-06 
0.05 4.843 0 0.0 1e-06 
3.0 4.843 0 0.0 1e-06 
0.05 4.844 0 0.0 1e-06 
3.0 4.844 0 0.0 1e-06 
0.05 4.845 0 0.0 1e-06 
3.0 4.845 0 0.0 1e-06 
0.05 4.846 0 0.0 1e-06 
3.0 4.846 0 0.0 1e-06 
0.05 4.847 0 0.0 1e-06 
3.0 4.847 0 0.0 1e-06 
0.05 4.848 0 0.0 1e-06 
3.0 4.848 0 0.0 1e-06 
0.05 4.849 0 0.0 1e-06 
3.0 4.849 0 0.0 1e-06 
0.05 4.85 0 0.0 1e-06 
3.0 4.85 0 0.0 1e-06 
0.05 4.851 0 0.0 1e-06 
3.0 4.851 0 0.0 1e-06 
0.05 4.852 0 0.0 1e-06 
3.0 4.852 0 0.0 1e-06 
0.05 4.853 0 0.0 1e-06 
3.0 4.853 0 0.0 1e-06 
0.05 4.854 0 0.0 1e-06 
3.0 4.854 0 0.0 1e-06 
0.05 4.855 0 0.0 1e-06 
3.0 4.855 0 0.0 1e-06 
0.05 4.856 0 0.0 1e-06 
3.0 4.856 0 0.0 1e-06 
0.05 4.857 0 0.0 1e-06 
3.0 4.857 0 0.0 1e-06 
0.05 4.858 0 0.0 1e-06 
3.0 4.858 0 0.0 1e-06 
0.05 4.859 0 0.0 1e-06 
3.0 4.859 0 0.0 1e-06 
0.05 4.86 0 0.0 1e-06 
3.0 4.86 0 0.0 1e-06 
0.05 4.861 0 0.0 1e-06 
3.0 4.861 0 0.0 1e-06 
0.05 4.862 0 0.0 1e-06 
3.0 4.862 0 0.0 1e-06 
0.05 4.863 0 0.0 1e-06 
3.0 4.863 0 0.0 1e-06 
0.05 4.864 0 0.0 1e-06 
3.0 4.864 0 0.0 1e-06 
0.05 4.865 0 0.0 1e-06 
3.0 4.865 0 0.0 1e-06 
0.05 4.866 0 0.0 1e-06 
3.0 4.866 0 0.0 1e-06 
0.05 4.867 0 0.0 1e-06 
3.0 4.867 0 0.0 1e-06 
0.05 4.868 0 0.0 1e-06 
3.0 4.868 0 0.0 1e-06 
0.05 4.869 0 0.0 1e-06 
3.0 4.869 0 0.0 1e-06 
0.05 4.87 0 0.0 1e-06 
3.0 4.87 0 0.0 1e-06 
0.05 4.871 0 0.0 1e-06 
3.0 4.871 0 0.0 1e-06 
0.05 4.872 0 0.0 1e-06 
3.0 4.872 0 0.0 1e-06 
0.05 4.873 0 0.0 1e-06 
3.0 4.873 0 0.0 1e-06 
0.05 4.874 0 0.0 1e-06 
3.0 4.874 0 0.0 1e-06 
0.05 4.875 0 0.0 1e-06 
3.0 4.875 0 0.0 1e-06 
0.05 4.876 0 0.0 1e-06 
3.0 4.876 0 0.0 1e-06 
0.05 4.877 0 0.0 1e-06 
3.0 4.877 0 0.0 1e-06 
0.05 4.878 0 0.0 1e-06 
3.0 4.878 0 0.0 1e-06 
0.05 4.879 0 0.0 1e-06 
3.0 4.879 0 0.0 1e-06 
0.05 4.88 0 0.0 1e-06 
3.0 4.88 0 0.0 1e-06 
0.05 4.881 0 0.0 1e-06 
3.0 4.881 0 0.0 1e-06 
0.05 4.882 0 0.0 1e-06 
3.0 4.882 0 0.0 1e-06 
0.05 4.883 0 0.0 1e-06 
3.0 4.883 0 0.0 1e-06 
0.05 4.884 0 0.0 1e-06 
3.0 4.884 0 0.0 1e-06 
0.05 4.885 0 0.0 1e-06 
3.0 4.885 0 0.0 1e-06 
0.05 4.886 0 0.0 1e-06 
3.0 4.886 0 0.0 1e-06 
0.05 4.887 0 0.0 1e-06 
3.0 4.887 0 0.0 1e-06 
0.05 4.888 0 0.0 1e-06 
3.0 4.888 0 0.0 1e-06 
0.05 4.889 0 0.0 1e-06 
3.0 4.889 0 0.0 1e-06 
0.05 4.89 0 0.0 1e-06 
3.0 4.89 0 0.0 1e-06 
0.05 4.891 0 0.0 1e-06 
3.0 4.891 0 0.0 1e-06 
0.05 4.892 0 0.0 1e-06 
3.0 4.892 0 0.0 1e-06 
0.05 4.893 0 0.0 1e-06 
3.0 4.893 0 0.0 1e-06 
0.05 4.894 0 0.0 1e-06 
3.0 4.894 0 0.0 1e-06 
0.05 4.895 0 0.0 1e-06 
3.0 4.895 0 0.0 1e-06 
0.05 4.896 0 0.0 1e-06 
3.0 4.896 0 0.0 1e-06 
0.05 4.897 0 0.0 1e-06 
3.0 4.897 0 0.0 1e-06 
0.05 4.898 0 0.0 1e-06 
3.0 4.898 0 0.0 1e-06 
0.05 4.899 0 0.0 1e-06 
3.0 4.899 0 0.0 1e-06 
0.05 4.9 0 0.0 1e-06 
3.0 4.9 0 0.0 1e-06 
0.05 4.901 0 0.0 1e-06 
3.0 4.901 0 0.0 1e-06 
0.05 4.902 0 0.0 1e-06 
3.0 4.902 0 0.0 1e-06 
0.05 4.903 0 0.0 1e-06 
3.0 4.903 0 0.0 1e-06 
0.05 4.904 0 0.0 1e-06 
3.0 4.904 0 0.0 1e-06 
0.05 4.905 0 0.0 1e-06 
3.0 4.905 0 0.0 1e-06 
0.05 4.906 0 0.0 1e-06 
3.0 4.906 0 0.0 1e-06 
0.05 4.907 0 0.0 1e-06 
3.0 4.907 0 0.0 1e-06 
0.05 4.908 0 0.0 1e-06 
3.0 4.908 0 0.0 1e-06 
0.05 4.909 0 0.0 1e-06 
3.0 4.909 0 0.0 1e-06 
0.05 4.91 0 0.0 1e-06 
3.0 4.91 0 0.0 1e-06 
0.05 4.911 0 0.0 1e-06 
3.0 4.911 0 0.0 1e-06 
0.05 4.912 0 0.0 1e-06 
3.0 4.912 0 0.0 1e-06 
0.05 4.913 0 0.0 1e-06 
3.0 4.913 0 0.0 1e-06 
0.05 4.914 0 0.0 1e-06 
3.0 4.914 0 0.0 1e-06 
0.05 4.915 0 0.0 1e-06 
3.0 4.915 0 0.0 1e-06 
0.05 4.916 0 0.0 1e-06 
3.0 4.916 0 0.0 1e-06 
0.05 4.917 0 0.0 1e-06 
3.0 4.917 0 0.0 1e-06 
0.05 4.918 0 0.0 1e-06 
3.0 4.918 0 0.0 1e-06 
0.05 4.919 0 0.0 1e-06 
3.0 4.919 0 0.0 1e-06 
0.05 4.92 0 0.0 1e-06 
3.0 4.92 0 0.0 1e-06 
0.05 4.921 0 0.0 1e-06 
3.0 4.921 0 0.0 1e-06 
0.05 4.922 0 0.0 1e-06 
3.0 4.922 0 0.0 1e-06 
0.05 4.923 0 0.0 1e-06 
3.0 4.923 0 0.0 1e-06 
0.05 4.924 0 0.0 1e-06 
3.0 4.924 0 0.0 1e-06 
0.05 4.925 0 0.0 1e-06 
3.0 4.925 0 0.0 1e-06 
0.05 4.926 0 0.0 1e-06 
3.0 4.926 0 0.0 1e-06 
0.05 4.927 0 0.0 1e-06 
3.0 4.927 0 0.0 1e-06 
0.05 4.928 0 0.0 1e-06 
3.0 4.928 0 0.0 1e-06 
0.05 4.929 0 0.0 1e-06 
3.0 4.929 0 0.0 1e-06 
0.05 4.93 0 0.0 1e-06 
3.0 4.93 0 0.0 1e-06 
0.05 4.931 0 0.0 1e-06 
3.0 4.931 0 0.0 1e-06 
0.05 4.932 0 0.0 1e-06 
3.0 4.932 0 0.0 1e-06 
0.05 4.933 0 0.0 1e-06 
3.0 4.933 0 0.0 1e-06 
0.05 4.934 0 0.0 1e-06 
3.0 4.934 0 0.0 1e-06 
0.05 4.935 0 0.0 1e-06 
3.0 4.935 0 0.0 1e-06 
0.05 4.936 0 0.0 1e-06 
3.0 4.936 0 0.0 1e-06 
0.05 4.937 0 0.0 1e-06 
3.0 4.937 0 0.0 1e-06 
0.05 4.938 0 0.0 1e-06 
3.0 4.938 0 0.0 1e-06 
0.05 4.939 0 0.0 1e-06 
3.0 4.939 0 0.0 1e-06 
0.05 4.94 0 0.0 1e-06 
3.0 4.94 0 0.0 1e-06 
0.05 4.941 0 0.0 1e-06 
3.0 4.941 0 0.0 1e-06 
0.05 4.942 0 0.0 1e-06 
3.0 4.942 0 0.0 1e-06 
0.05 4.943 0 0.0 1e-06 
3.0 4.943 0 0.0 1e-06 
0.05 4.944 0 0.0 1e-06 
3.0 4.944 0 0.0 1e-06 
0.05 4.945 0 0.0 1e-06 
3.0 4.945 0 0.0 1e-06 
0.05 4.946 0 0.0 1e-06 
3.0 4.946 0 0.0 1e-06 
0.05 4.947 0 0.0 1e-06 
3.0 4.947 0 0.0 1e-06 
0.05 4.948 0 0.0 1e-06 
3.0 4.948 0 0.0 1e-06 
0.05 4.949 0 0.0 1e-06 
3.0 4.949 0 0.0 1e-06 
0.05 4.95 0 0.0 1e-06 
3.0 4.95 0 0.0 1e-06 
0.05 4.951 0 0.0 1e-06 
3.0 4.951 0 0.0 1e-06 
0.05 4.952 0 0.0 1e-06 
3.0 4.952 0 0.0 1e-06 
0.05 4.953 0 0.0 1e-06 
3.0 4.953 0 0.0 1e-06 
0.05 4.954 0 0.0 1e-06 
3.0 4.954 0 0.0 1e-06 
0.05 4.955 0 0.0 1e-06 
3.0 4.955 0 0.0 1e-06 
0.05 4.956 0 0.0 1e-06 
3.0 4.956 0 0.0 1e-06 
0.05 4.957 0 0.0 1e-06 
3.0 4.957 0 0.0 1e-06 
0.05 4.958 0 0.0 1e-06 
3.0 4.958 0 0.0 1e-06 
0.05 4.959 0 0.0 1e-06 
3.0 4.959 0 0.0 1e-06 
0.05 4.96 0 0.0 1e-06 
3.0 4.96 0 0.0 1e-06 
0.05 4.961 0 0.0 1e-06 
3.0 4.961 0 0.0 1e-06 
0.05 4.962 0 0.0 1e-06 
3.0 4.962 0 0.0 1e-06 
0.05 4.963 0 0.0 1e-06 
3.0 4.963 0 0.0 1e-06 
0.05 4.964 0 0.0 1e-06 
3.0 4.964 0 0.0 1e-06 
0.05 4.965 0 0.0 1e-06 
3.0 4.965 0 0.0 1e-06 
0.05 4.966 0 0.0 1e-06 
3.0 4.966 0 0.0 1e-06 
0.05 4.967 0 0.0 1e-06 
3.0 4.967 0 0.0 1e-06 
0.05 4.968 0 0.0 1e-06 
3.0 4.968 0 0.0 1e-06 
0.05 4.969 0 0.0 1e-06 
3.0 4.969 0 0.0 1e-06 
0.05 4.97 0 0.0 1e-06 
3.0 4.97 0 0.0 1e-06 
0.05 4.971 0 0.0 1e-06 
3.0 4.971 0 0.0 1e-06 
0.05 4.972 0 0.0 1e-06 
3.0 4.972 0 0.0 1e-06 
0.05 4.973 0 0.0 1e-06 
3.0 4.973 0 0.0 1e-06 
0.05 4.974 0 0.0 1e-06 
3.0 4.974 0 0.0 1e-06 
0.05 4.975 0 0.0 1e-06 
3.0 4.975 0 0.0 1e-06 
0.05 4.976 0 0.0 1e-06 
3.0 4.976 0 0.0 1e-06 
0.05 4.977 0 0.0 1e-06 
3.0 4.977 0 0.0 1e-06 
0.05 4.978 0 0.0 1e-06 
3.0 4.978 0 0.0 1e-06 
0.05 4.979 0 0.0 1e-06 
3.0 4.979 0 0.0 1e-06 
0.05 4.98 0 0.0 1e-06 
3.0 4.98 0 0.0 1e-06 
0.05 4.981 0 0.0 1e-06 
3.0 4.981 0 0.0 1e-06 
0.05 4.982 0 0.0 1e-06 
3.0 4.982 0 0.0 1e-06 
0.05 4.983 0 0.0 1e-06 
3.0 4.983 0 0.0 1e-06 
0.05 4.984 0 0.0 1e-06 
3.0 4.984 0 0.0 1e-06 
0.05 4.985 0 0.0 1e-06 
3.0 4.985 0 0.0 1e-06 
0.05 4.986 0 0.0 1e-06 
3.0 4.986 0 0.0 1e-06 
0.05 4.987 0 0.0 1e-06 
3.0 4.987 0 0.0 1e-06 
0.05 4.988 0 0.0 1e-06 
3.0 4.988 0 0.0 1e-06 
0.05 4.989 0 0.0 1e-06 
3.0 4.989 0 0.0 1e-06 
0.05 4.99 0 0.0 1e-06 
3.0 4.99 0 0.0 1e-06 
0.05 4.991 0 0.0 1e-06 
3.0 4.991 0 0.0 1e-06 
0.05 4.992 0 0.0 1e-06 
3.0 4.992 0 0.0 1e-06 
0.05 4.993 0 0.0 1e-06 
3.0 4.993 0 0.0 1e-06 
0.05 4.994 0 0.0 1e-06 
3.0 4.994 0 0.0 1e-06 
0.05 4.995 0 0.0 1e-06 
3.0 4.995 0 0.0 1e-06 
0.05 4.996 0 0.0 1e-06 
3.0 4.996 0 0.0 1e-06 
0.05 4.997 0 0.0 1e-06 
3.0 4.997 0 0.0 1e-06 
0.05 4.998 0 0.0 1e-06 
3.0 4.998 0 0.0 1e-06 
0.05 4.999 0 0.0 1e-06 
3.0 4.999 0 0.0 1e-06 
0.05 0.0 0 3.0 1e-06 
3.0 0.0 0 3.0 1e-06 
0.05 0.001 0 3.0 1e-06 
3.0 0.001 0 3.0 1e-06 
0.05 0.002 0 3.0 1e-06 
3.0 0.002 0 3.0 1e-06 
0.05 0.003 0 3.0 1e-06 
3.0 0.003 0 3.0 1e-06 
0.05 0.004 0 3.0 1e-06 
3.0 0.004 0 3.0 1e-06 
0.05 0.005 0 3.0 1e-06 
3.0 0.005 0 3.0 1e-06 
0.05 0.006 0 3.0 1e-06 
3.0 0.006 0 3.0 1e-06 
0.05 0.007 0 3.0 1e-06 
3.0 0.007 0 3.0 1e-06 
0.05 0.008 0 3.0 1e-06 
3.0 0.008 0 3.0 1e-06 
0.05 0.009 0 3.0 1e-06 
3.0 0.009 0 3.0 1e-06 
0.05 0.01 0 3.0 1e-06 
3.0 0.01 0 3.0 1e-06 
0.05 0.011 0 3.0 1e-06 
3.0 0.011 0 3.0 1e-06 
0.05 0.012 0 3.0 1e-06 
3.0 0.012 0 3.0 1e-06 
0.05 0.013 0 3.0 1e-06 
3.0 0.013 0 3.0 1e-06 
0.05 0.014 0 3.0 1e-06 
3.0 0.014 0 3.0 1e-06 
0.05 0.015 0 3.0 1e-06 
3.0 0.015 0 3.0 1e-06 
0.05 0.016 0 3.0 1e-06 
3.0 0.016 0 3.0 1e-06 
0.05 0.017 0 3.0 1e-06 
3.0 0.017 0 3.0 1e-06 
0.05 0.018 0 3.0 1e-06 
3.0 0.018 0 3.0 1e-06 
0.05 0.019 0 3.0 1e-06 
3.0 0.019 0 3.0 1e-06 
0.05 0.02 0 3.0 1e-06 
3.0 0.02 0 3.0 1e-06 
0.05 0.021 0 3.0 1e-06 
3.0 0.021 0 3.0 1e-06 
0.05 0.022 0 3.0 1e-06 
3.0 0.022 0 3.0 1e-06 
0.05 0.023 0 3.0 1e-06 
3.0 0.023 0 3.0 1e-06 
0.05 0.024 0 3.0 1e-06 
3.0 0.024 0 3.0 1e-06 
0.05 0.025 0 3.0 1e-06 
3.0 0.025 0 3.0 1e-06 
0.05 0.026 0 3.0 1e-06 
3.0 0.026 0 3.0 1e-06 
0.05 0.027 0 3.0 1e-06 
3.0 0.027 0 3.0 1e-06 
0.05 0.028 0 3.0 1e-06 
3.0 0.028 0 3.0 1e-06 
0.05 0.029 0 3.0 1e-06 
3.0 0.029 0 3.0 1e-06 
0.05 0.03 0 3.0 1e-06 
3.0 0.03 0 3.0 1e-06 
0.05 0.031 0 3.0 1e-06 
3.0 0.031 0 3.0 1e-06 
0.05 0.032 0 3.0 1e-06 
3.0 0.032 0 3.0 1e-06 
0.05 0.033 0 3.0 1e-06 
3.0 0.033 0 3.0 1e-06 
0.05 0.034 0 3.0 1e-06 
3.0 0.034 0 3.0 1e-06 
0.05 0.035 0 3.0 1e-06 
3.0 0.035 0 3.0 1e-06 
0.05 0.036 0 3.0 1e-06 
3.0 0.036 0 3.0 1e-06 
0.05 0.037 0 3.0 1e-06 
3.0 0.037 0 3.0 1e-06 
0.05 0.038 0 3.0 1e-06 
3.0 0.038 0 3.0 1e-06 
0.05 0.039 0 3.0 1e-06 
3.0 0.039 0 3.0 1e-06 
0.05 0.04 0 3.0 1e-06 
3.0 0.04 0 3.0 1e-06 
0.05 0.041 0 3.0 1e-06 
3.0 0.041 0 3.0 1e-06 
0.05 0.042 0 3.0 1e-06 
3.0 0.042 0 3.0 1e-06 
0.05 0.043 0 3.0 1e-06 
3.0 0.043 0 3.0 1e-06 
0.05 0.044 0 3.0 1e-06 
3.0 0.044 0 3.0 1e-06 
0.05 0.045 0 3.0 1e-06 
3.0 0.045 0 3.0 1e-06 
0.05 0.046 0 3.0 1e-06 
3.0 0.046 0 3.0 1e-06 
0.05 0.047 0 3.0 1e-06 
3.0 0.047 0 3.0 1e-06 
0.05 0.048 0 3.0 1e-06 
3.0 0.048 0 3.0 1e-06 
0.05 0.049 0 3.0 1e-06 
3.0 0.049 0 3.0 1e-06 
0.05 0.05 0 3.0 1e-06 
3.0 0.05 0 3.0 1e-06 
0.05 0.051 0 3.0 1e-06 
3.0 0.051 0 3.0 1e-06 
0.05 0.052 0 3.0 1e-06 
3.0 0.052 0 3.0 1e-06 
0.05 0.053 0 3.0 1e-06 
3.0 0.053 0 3.0 1e-06 
0.05 0.054 0 3.0 1e-06 
3.0 0.054 0 3.0 1e-06 
0.05 0.055 0 3.0 1e-06 
3.0 0.055 0 3.0 1e-06 
0.05 0.056 0 3.0 1e-06 
3.0 0.056 0 3.0 1e-06 
0.05 0.057 0 3.0 1e-06 
3.0 0.057 0 3.0 1e-06 
0.05 0.058 0 3.0 1e-06 
3.0 0.058 0 3.0 1e-06 
0.05 0.059 0 3.0 1e-06 
3.0 0.059 0 3.0 1e-06 
0.05 0.06 0 3.0 1e-06 
3.0 0.06 0 3.0 1e-06 
0.05 0.061 0 3.0 1e-06 
3.0 0.061 0 3.0 1e-06 
0.05 0.062 0 3.0 1e-06 
3.0 0.062 0 3.0 1e-06 
0.05 0.063 0 3.0 1e-06 
3.0 0.063 0 3.0 1e-06 
0.05 0.064 0 3.0 1e-06 
3.0 0.064 0 3.0 1e-06 
0.05 0.065 0 3.0 1e-06 
3.0 0.065 0 3.0 1e-06 
0.05 0.066 0 3.0 1e-06 
3.0 0.066 0 3.0 1e-06 
0.05 0.067 0 3.0 1e-06 
3.0 0.067 0 3.0 1e-06 
0.05 0.068 0 3.0 1e-06 
3.0 0.068 0 3.0 1e-06 
0.05 0.069 0 3.0 1e-06 
3.0 0.069 0 3.0 1e-06 
0.05 0.07 0 3.0 1e-06 
3.0 0.07 0 3.0 1e-06 
0.05 0.071 0 3.0 1e-06 
3.0 0.071 0 3.0 1e-06 
0.05 0.072 0 3.0 1e-06 
3.0 0.072 0 3.0 1e-06 
0.05 0.073 0 3.0 1e-06 
3.0 0.073 0 3.0 1e-06 
0.05 0.074 0 3.0 1e-06 
3.0 0.074 0 3.0 1e-06 
0.05 0.075 0 3.0 1e-06 
3.0 0.075 0 3.0 1e-06 
0.05 0.076 0 3.0 1e-06 
3.0 0.076 0 3.0 1e-06 
0.05 0.077 0 3.0 1e-06 
3.0 0.077 0 3.0 1e-06 
0.05 0.078 0 3.0 1e-06 
3.0 0.078 0 3.0 1e-06 
0.05 0.079 0 3.0 1e-06 
3.0 0.079 0 3.0 1e-06 
0.05 0.08 0 3.0 1e-06 
3.0 0.08 0 3.0 1e-06 
0.05 0.081 0 3.0 1e-06 
3.0 0.081 0 3.0 1e-06 
0.05 0.082 0 3.0 1e-06 
3.0 0.082 0 3.0 1e-06 
0.05 0.083 0 3.0 1e-06 
3.0 0.083 0 3.0 1e-06 
0.05 0.084 0 3.0 1e-06 
3.0 0.084 0 3.0 1e-06 
0.05 0.085 0 3.0 1e-06 
3.0 0.085 0 3.0 1e-06 
0.05 0.086 0 3.0 1e-06 
3.0 0.086 0 3.0 1e-06 
0.05 0.087 0 3.0 1e-06 
3.0 0.087 0 3.0 1e-06 
0.05 0.088 0 3.0 1e-06 
3.0 0.088 0 3.0 1e-06 
0.05 0.089 0 3.0 1e-06 
3.0 0.089 0 3.0 1e-06 
0.05 0.09 0 3.0 1e-06 
3.0 0.09 0 3.0 1e-06 
0.05 0.091 0 3.0 1e-06 
3.0 0.091 0 3.0 1e-06 
0.05 0.092 0 3.0 1e-06 
3.0 0.092 0 3.0 1e-06 
0.05 0.093 0 3.0 1e-06 
3.0 0.093 0 3.0 1e-06 
0.05 0.094 0 3.0 1e-06 
3.0 0.094 0 3.0 1e-06 
0.05 0.095 0 3.0 1e-06 
3.0 0.095 0 3.0 1e-06 
0.05 0.096 0 3.0 1e-06 
3.0 0.096 0 3.0 1e-06 
0.05 0.097 0 3.0 1e-06 
3.0 0.097 0 3.0 1e-06 
0.05 0.098 0 3.0 1e-06 
3.0 0.098 0 3.0 1e-06 
0.05 0.099 0 3.0 1e-06 
3.0 0.099 0 3.0 1e-06 
0.05 0.1 0 3.0 1e-06 
3.0 0.1 0 3.0 1e-06 
0.05 0.101 0 3.0 1e-06 
3.0 0.101 0 3.0 1e-06 
0.05 0.102 0 3.0 1e-06 
3.0 0.102 0 3.0 1e-06 
0.05 0.103 0 3.0 1e-06 
3.0 0.103 0 3.0 1e-06 
0.05 0.104 0 3.0 1e-06 
3.0 0.104 0 3.0 1e-06 
0.05 0.105 0 3.0 1e-06 
3.0 0.105 0 3.0 1e-06 
0.05 0.106 0 3.0 1e-06 
3.0 0.106 0 3.0 1e-06 
0.05 0.107 0 3.0 1e-06 
3.0 0.107 0 3.0 1e-06 
0.05 0.108 0 3.0 1e-06 
3.0 0.108 0 3.0 1e-06 
0.05 0.109 0 3.0 1e-06 
3.0 0.109 0 3.0 1e-06 
0.05 0.11 0 3.0 1e-06 
3.0 0.11 0 3.0 1e-06 
0.05 0.111 0 3.0 1e-06 
3.0 0.111 0 3.0 1e-06 
0.05 0.112 0 3.0 1e-06 
3.0 0.112 0 3.0 1e-06 
0.05 0.113 0 3.0 1e-06 
3.0 0.113 0 3.0 1e-06 
0.05 0.114 0 3.0 1e-06 
3.0 0.114 0 3.0 1e-06 
0.05 0.115 0 3.0 1e-06 
3.0 0.115 0 3.0 1e-06 
0.05 0.116 0 3.0 1e-06 
3.0 0.116 0 3.0 1e-06 
0.05 0.117 0 3.0 1e-06 
3.0 0.117 0 3.0 1e-06 
0.05 0.118 0 3.0 1e-06 
3.0 0.118 0 3.0 1e-06 
0.05 0.119 0 3.0 1e-06 
3.0 0.119 0 3.0 1e-06 
0.05 0.12 0 3.0 1e-06 
3.0 0.12 0 3.0 1e-06 
0.05 0.121 0 3.0 1e-06 
3.0 0.121 0 3.0 1e-06 
0.05 0.122 0 3.0 1e-06 
3.0 0.122 0 3.0 1e-06 
0.05 0.123 0 3.0 1e-06 
3.0 0.123 0 3.0 1e-06 
0.05 0.124 0 3.0 1e-06 
3.0 0.124 0 3.0 1e-06 
0.05 0.125 0 3.0 1e-06 
3.0 0.125 0 3.0 1e-06 
0.05 0.126 0 3.0 1e-06 
3.0 0.126 0 3.0 1e-06 
0.05 0.127 0 3.0 1e-06 
3.0 0.127 0 3.0 1e-06 
0.05 0.128 0 3.0 1e-06 
3.0 0.128 0 3.0 1e-06 
0.05 0.129 0 3.0 1e-06 
3.0 0.129 0 3.0 1e-06 
0.05 0.13 0 3.0 1e-06 
3.0 0.13 0 3.0 1e-06 
0.05 0.131 0 3.0 1e-06 
3.0 0.131 0 3.0 1e-06 
0.05 0.132 0 3.0 1e-06 
3.0 0.132 0 3.0 1e-06 
0.05 0.133 0 3.0 1e-06 
3.0 0.133 0 3.0 1e-06 
0.05 0.134 0 3.0 1e-06 
3.0 0.134 0 3.0 1e-06 
0.05 0.135 0 3.0 1e-06 
3.0 0.135 0 3.0 1e-06 
0.05 0.136 0 3.0 1e-06 
3.0 0.136 0 3.0 1e-06 
0.05 0.137 0 3.0 1e-06 
3.0 0.137 0 3.0 1e-06 
0.05 0.138 0 3.0 1e-06 
3.0 0.138 0 3.0 1e-06 
0.05 0.139 0 3.0 1e-06 
3.0 0.139 0 3.0 1e-06 
0.05 0.14 0 3.0 1e-06 
3.0 0.14 0 3.0 1e-06 
0.05 0.141 0 3.0 1e-06 
3.0 0.141 0 3.0 1e-06 
0.05 0.142 0 3.0 1e-06 
3.0 0.142 0 3.0 1e-06 
0.05 0.143 0 3.0 1e-06 
3.0 0.143 0 3.0 1e-06 
0.05 0.144 0 3.0 1e-06 
3.0 0.144 0 3.0 1e-06 
0.05 0.145 0 3.0 1e-06 
3.0 0.145 0 3.0 1e-06 
0.05 0.146 0 3.0 1e-06 
3.0 0.146 0 3.0 1e-06 
0.05 0.147 0 3.0 1e-06 
3.0 0.147 0 3.0 1e-06 
0.05 0.148 0 3.0 1e-06 
3.0 0.148 0 3.0 1e-06 
0.05 0.149 0 3.0 1e-06 
3.0 0.149 0 3.0 1e-06 
0.05 0.15 0 3.0 1e-06 
3.0 0.15 0 3.0 1e-06 
0.05 0.151 0 3.0 1e-06 
3.0 0.151 0 3.0 1e-06 
0.05 0.152 0 3.0 1e-06 
3.0 0.152 0 3.0 1e-06 
0.05 0.153 0 3.0 1e-06 
3.0 0.153 0 3.0 1e-06 
0.05 0.154 0 3.0 1e-06 
3.0 0.154 0 3.0 1e-06 
0.05 0.155 0 3.0 1e-06 
3.0 0.155 0 3.0 1e-06 
0.05 0.156 0 3.0 1e-06 
3.0 0.156 0 3.0 1e-06 
0.05 0.157 0 3.0 1e-06 
3.0 0.157 0 3.0 1e-06 
0.05 0.158 0 3.0 1e-06 
3.0 0.158 0 3.0 1e-06 
0.05 0.159 0 3.0 1e-06 
3.0 0.159 0 3.0 1e-06 
0.05 0.16 0 3.0 1e-06 
3.0 0.16 0 3.0 1e-06 
0.05 0.161 0 3.0 1e-06 
3.0 0.161 0 3.0 1e-06 
0.05 0.162 0 3.0 1e-06 
3.0 0.162 0 3.0 1e-06 
0.05 0.163 0 3.0 1e-06 
3.0 0.163 0 3.0 1e-06 
0.05 0.164 0 3.0 1e-06 
3.0 0.164 0 3.0 1e-06 
0.05 0.165 0 3.0 1e-06 
3.0 0.165 0 3.0 1e-06 
0.05 0.166 0 3.0 1e-06 
3.0 0.166 0 3.0 1e-06 
0.05 0.167 0 3.0 1e-06 
3.0 0.167 0 3.0 1e-06 
0.05 0.168 0 3.0 1e-06 
3.0 0.168 0 3.0 1e-06 
0.05 0.169 0 3.0 1e-06 
3.0 0.169 0 3.0 1e-06 
0.05 0.17 0 3.0 1e-06 
3.0 0.17 0 3.0 1e-06 
0.05 0.171 0 3.0 1e-06 
3.0 0.171 0 3.0 1e-06 
0.05 0.172 0 3.0 1e-06 
3.0 0.172 0 3.0 1e-06 
0.05 0.173 0 3.0 1e-06 
3.0 0.173 0 3.0 1e-06 
0.05 0.174 0 3.0 1e-06 
3.0 0.174 0 3.0 1e-06 
0.05 0.175 0 3.0 1e-06 
3.0 0.175 0 3.0 1e-06 
0.05 0.176 0 3.0 1e-06 
3.0 0.176 0 3.0 1e-06 
0.05 0.177 0 3.0 1e-06 
3.0 0.177 0 3.0 1e-06 
0.05 0.178 0 3.0 1e-06 
3.0 0.178 0 3.0 1e-06 
0.05 0.179 0 3.0 1e-06 
3.0 0.179 0 3.0 1e-06 
0.05 0.18 0 3.0 1e-06 
3.0 0.18 0 3.0 1e-06 
0.05 0.181 0 3.0 1e-06 
3.0 0.181 0 3.0 1e-06 
0.05 0.182 0 3.0 1e-06 
3.0 0.182 0 3.0 1e-06 
0.05 0.183 0 3.0 1e-06 
3.0 0.183 0 3.0 1e-06 
0.05 0.184 0 3.0 1e-06 
3.0 0.184 0 3.0 1e-06 
0.05 0.185 0 3.0 1e-06 
3.0 0.185 0 3.0 1e-06 
0.05 0.186 0 3.0 1e-06 
3.0 0.186 0 3.0 1e-06 
0.05 0.187 0 3.0 1e-06 
3.0 0.187 0 3.0 1e-06 
0.05 0.188 0 3.0 1e-06 
3.0 0.188 0 3.0 1e-06 
0.05 0.189 0 3.0 1e-06 
3.0 0.189 0 3.0 1e-06 
0.05 0.19 0 3.0 1e-06 
3.0 0.19 0 3.0 1e-06 
0.05 0.191 0 3.0 1e-06 
3.0 0.191 0 3.0 1e-06 
0.05 0.192 0 3.0 1e-06 
3.0 0.192 0 3.0 1e-06 
0.05 0.193 0 3.0 1e-06 
3.0 0.193 0 3.0 1e-06 
0.05 0.194 0 3.0 1e-06 
3.0 0.194 0 3.0 1e-06 
0.05 0.195 0 3.0 1e-06 
3.0 0.195 0 3.0 1e-06 
0.05 0.196 0 3.0 1e-06 
3.0 0.196 0 3.0 1e-06 
0.05 0.197 0 3.0 1e-06 
3.0 0.197 0 3.0 1e-06 
0.05 0.198 0 3.0 1e-06 
3.0 0.198 0 3.0 1e-06 
0.05 0.199 0 3.0 1e-06 
3.0 0.199 0 3.0 1e-06 
0.05 0.2 0 3.0 1e-06 
3.0 0.2 0 3.0 1e-06 
0.05 0.201 0 3.0 1e-06 
3.0 0.201 0 3.0 1e-06 
0.05 0.202 0 3.0 1e-06 
3.0 0.202 0 3.0 1e-06 
0.05 0.203 0 3.0 1e-06 
3.0 0.203 0 3.0 1e-06 
0.05 0.204 0 3.0 1e-06 
3.0 0.204 0 3.0 1e-06 
0.05 0.205 0 3.0 1e-06 
3.0 0.205 0 3.0 1e-06 
0.05 0.206 0 3.0 1e-06 
3.0 0.206 0 3.0 1e-06 
0.05 0.207 0 3.0 1e-06 
3.0 0.207 0 3.0 1e-06 
0.05 0.208 0 3.0 1e-06 
3.0 0.208 0 3.0 1e-06 
0.05 0.209 0 3.0 1e-06 
3.0 0.209 0 3.0 1e-06 
0.05 0.21 0 3.0 1e-06 
3.0 0.21 0 3.0 1e-06 
0.05 0.211 0 3.0 1e-06 
3.0 0.211 0 3.0 1e-06 
0.05 0.212 0 3.0 1e-06 
3.0 0.212 0 3.0 1e-06 
0.05 0.213 0 3.0 1e-06 
3.0 0.213 0 3.0 1e-06 
0.05 0.214 0 3.0 1e-06 
3.0 0.214 0 3.0 1e-06 
0.05 0.215 0 3.0 1e-06 
3.0 0.215 0 3.0 1e-06 
0.05 0.216 0 3.0 1e-06 
3.0 0.216 0 3.0 1e-06 
0.05 0.217 0 3.0 1e-06 
3.0 0.217 0 3.0 1e-06 
0.05 0.218 0 3.0 1e-06 
3.0 0.218 0 3.0 1e-06 
0.05 0.219 0 3.0 1e-06 
3.0 0.219 0 3.0 1e-06 
0.05 0.22 0 3.0 1e-06 
3.0 0.22 0 3.0 1e-06 
0.05 0.221 0 3.0 1e-06 
3.0 0.221 0 3.0 1e-06 
0.05 0.222 0 3.0 1e-06 
3.0 0.222 0 3.0 1e-06 
0.05 0.223 0 3.0 1e-06 
3.0 0.223 0 3.0 1e-06 
0.05 0.224 0 3.0 1e-06 
3.0 0.224 0 3.0 1e-06 
0.05 0.225 0 3.0 1e-06 
3.0 0.225 0 3.0 1e-06 
0.05 0.226 0 3.0 1e-06 
3.0 0.226 0 3.0 1e-06 
0.05 0.227 0 3.0 1e-06 
3.0 0.227 0 3.0 1e-06 
0.05 0.228 0 3.0 1e-06 
3.0 0.228 0 3.0 1e-06 
0.05 0.229 0 3.0 1e-06 
3.0 0.229 0 3.0 1e-06 
0.05 0.23 0 3.0 1e-06 
3.0 0.23 0 3.0 1e-06 
0.05 0.231 0 3.0 1e-06 
3.0 0.231 0 3.0 1e-06 
0.05 0.232 0 3.0 1e-06 
3.0 0.232 0 3.0 1e-06 
0.05 0.233 0 3.0 1e-06 
3.0 0.233 0 3.0 1e-06 
0.05 0.234 0 3.0 1e-06 
3.0 0.234 0 3.0 1e-06 
0.05 0.235 0 3.0 1e-06 
3.0 0.235 0 3.0 1e-06 
0.05 0.236 0 3.0 1e-06 
3.0 0.236 0 3.0 1e-06 
0.05 0.237 0 3.0 1e-06 
3.0 0.237 0 3.0 1e-06 
0.05 0.238 0 3.0 1e-06 
3.0 0.238 0 3.0 1e-06 
0.05 0.239 0 3.0 1e-06 
3.0 0.239 0 3.0 1e-06 
0.05 0.24 0 3.0 1e-06 
3.0 0.24 0 3.0 1e-06 
0.05 0.241 0 3.0 1e-06 
3.0 0.241 0 3.0 1e-06 
0.05 0.242 0 3.0 1e-06 
3.0 0.242 0 3.0 1e-06 
0.05 0.243 0 3.0 1e-06 
3.0 0.243 0 3.0 1e-06 
0.05 0.244 0 3.0 1e-06 
3.0 0.244 0 3.0 1e-06 
0.05 0.245 0 3.0 1e-06 
3.0 0.245 0 3.0 1e-06 
0.05 0.246 0 3.0 1e-06 
3.0 0.246 0 3.0 1e-06 
0.05 0.247 0 3.0 1e-06 
3.0 0.247 0 3.0 1e-06 
0.05 0.248 0 3.0 1e-06 
3.0 0.248 0 3.0 1e-06 
0.05 0.249 0 3.0 1e-06 
3.0 0.249 0 3.0 1e-06 
0.05 0.25 0 3.0 1e-06 
3.0 0.25 0 3.0 1e-06 
0.05 0.251 0 3.0 1e-06 
3.0 0.251 0 3.0 1e-06 
0.05 0.252 0 3.0 1e-06 
3.0 0.252 0 3.0 1e-06 
0.05 0.253 0 3.0 1e-06 
3.0 0.253 0 3.0 1e-06 
0.05 0.254 0 3.0 1e-06 
3.0 0.254 0 3.0 1e-06 
0.05 0.255 0 3.0 1e-06 
3.0 0.255 0 3.0 1e-06 
0.05 0.256 0 3.0 1e-06 
3.0 0.256 0 3.0 1e-06 
0.05 0.257 0 3.0 1e-06 
3.0 0.257 0 3.0 1e-06 
0.05 0.258 0 3.0 1e-06 
3.0 0.258 0 3.0 1e-06 
0.05 0.259 0 3.0 1e-06 
3.0 0.259 0 3.0 1e-06 
0.05 0.26 0 3.0 1e-06 
3.0 0.26 0 3.0 1e-06 
0.05 0.261 0 3.0 1e-06 
3.0 0.261 0 3.0 1e-06 
0.05 0.262 0 3.0 1e-06 
3.0 0.262 0 3.0 1e-06 
0.05 0.263 0 3.0 1e-06 
3.0 0.263 0 3.0 1e-06 
0.05 0.264 0 3.0 1e-06 
3.0 0.264 0 3.0 1e-06 
0.05 0.265 0 3.0 1e-06 
3.0 0.265 0 3.0 1e-06 
0.05 0.266 0 3.0 1e-06 
3.0 0.266 0 3.0 1e-06 
0.05 0.267 0 3.0 1e-06 
3.0 0.267 0 3.0 1e-06 
0.05 0.268 0 3.0 1e-06 
3.0 0.268 0 3.0 1e-06 
0.05 0.269 0 3.0 1e-06 
3.0 0.269 0 3.0 1e-06 
0.05 0.27 0 3.0 1e-06 
3.0 0.27 0 3.0 1e-06 
0.05 0.271 0 3.0 1e-06 
3.0 0.271 0 3.0 1e-06 
0.05 0.272 0 3.0 1e-06 
3.0 0.272 0 3.0 1e-06 
0.05 0.273 0 3.0 1e-06 
3.0 0.273 0 3.0 1e-06 
0.05 0.274 0 3.0 1e-06 
3.0 0.274 0 3.0 1e-06 
0.05 0.275 0 3.0 1e-06 
3.0 0.275 0 3.0 1e-06 
0.05 0.276 0 3.0 1e-06 
3.0 0.276 0 3.0 1e-06 
0.05 0.277 0 3.0 1e-06 
3.0 0.277 0 3.0 1e-06 
0.05 0.278 0 3.0 1e-06 
3.0 0.278 0 3.0 1e-06 
0.05 0.279 0 3.0 1e-06 
3.0 0.279 0 3.0 1e-06 
0.05 0.28 0 3.0 1e-06 
3.0 0.28 0 3.0 1e-06 
0.05 0.281 0 3.0 1e-06 
3.0 0.281 0 3.0 1e-06 
0.05 0.282 0 3.0 1e-06 
3.0 0.282 0 3.0 1e-06 
0.05 0.283 0 3.0 1e-06 
3.0 0.283 0 3.0 1e-06 
0.05 0.284 0 3.0 1e-06 
3.0 0.284 0 3.0 1e-06 
0.05 0.285 0 3.0 1e-06 
3.0 0.285 0 3.0 1e-06 
0.05 0.286 0 3.0 1e-06 
3.0 0.286 0 3.0 1e-06 
0.05 0.287 0 3.0 1e-06 
3.0 0.287 0 3.0 1e-06 
0.05 0.288 0 3.0 1e-06 
3.0 0.288 0 3.0 1e-06 
0.05 0.289 0 3.0 1e-06 
3.0 0.289 0 3.0 1e-06 
0.05 0.29 0 3.0 1e-06 
3.0 0.29 0 3.0 1e-06 
0.05 0.291 0 3.0 1e-06 
3.0 0.291 0 3.0 1e-06 
0.05 0.292 0 3.0 1e-06 
3.0 0.292 0 3.0 1e-06 
0.05 0.293 0 3.0 1e-06 
3.0 0.293 0 3.0 1e-06 
0.05 0.294 0 3.0 1e-06 
3.0 0.294 0 3.0 1e-06 
0.05 0.295 0 3.0 1e-06 
3.0 0.295 0 3.0 1e-06 
0.05 0.296 0 3.0 1e-06 
3.0 0.296 0 3.0 1e-06 
0.05 0.297 0 3.0 1e-06 
3.0 0.297 0 3.0 1e-06 
0.05 0.298 0 3.0 1e-06 
3.0 0.298 0 3.0 1e-06 
0.05 0.299 0 3.0 1e-06 
3.0 0.299 0 3.0 1e-06 
0.05 0.3 0 3.0 1e-06 
3.0 0.3 0 3.0 1e-06 
0.05 0.301 0 3.0 1e-06 
3.0 0.301 0 3.0 1e-06 
0.05 0.302 0 3.0 1e-06 
3.0 0.302 0 3.0 1e-06 
0.05 0.303 0 3.0 1e-06 
3.0 0.303 0 3.0 1e-06 
0.05 0.304 0 3.0 1e-06 
3.0 0.304 0 3.0 1e-06 
0.05 0.305 0 3.0 1e-06 
3.0 0.305 0 3.0 1e-06 
0.05 0.306 0 3.0 1e-06 
3.0 0.306 0 3.0 1e-06 
0.05 0.307 0 3.0 1e-06 
3.0 0.307 0 3.0 1e-06 
0.05 0.308 0 3.0 1e-06 
3.0 0.308 0 3.0 1e-06 
0.05 0.309 0 3.0 1e-06 
3.0 0.309 0 3.0 1e-06 
0.05 0.31 0 3.0 1e-06 
3.0 0.31 0 3.0 1e-06 
0.05 0.311 0 3.0 1e-06 
3.0 0.311 0 3.0 1e-06 
0.05 0.312 0 3.0 1e-06 
3.0 0.312 0 3.0 1e-06 
0.05 0.313 0 3.0 1e-06 
3.0 0.313 0 3.0 1e-06 
0.05 0.314 0 3.0 1e-06 
3.0 0.314 0 3.0 1e-06 
0.05 0.315 0 3.0 1e-06 
3.0 0.315 0 3.0 1e-06 
0.05 0.316 0 3.0 1e-06 
3.0 0.316 0 3.0 1e-06 
0.05 0.317 0 3.0 1e-06 
3.0 0.317 0 3.0 1e-06 
0.05 0.318 0 3.0 1e-06 
3.0 0.318 0 3.0 1e-06 
0.05 0.319 0 3.0 1e-06 
3.0 0.319 0 3.0 1e-06 
0.05 0.32 0 3.0 1e-06 
3.0 0.32 0 3.0 1e-06 
0.05 0.321 0 3.0 1e-06 
3.0 0.321 0 3.0 1e-06 
0.05 0.322 0 3.0 1e-06 
3.0 0.322 0 3.0 1e-06 
0.05 0.323 0 3.0 1e-06 
3.0 0.323 0 3.0 1e-06 
0.05 0.324 0 3.0 1e-06 
3.0 0.324 0 3.0 1e-06 
0.05 0.325 0 3.0 1e-06 
3.0 0.325 0 3.0 1e-06 
0.05 0.326 0 3.0 1e-06 
3.0 0.326 0 3.0 1e-06 
0.05 0.327 0 3.0 1e-06 
3.0 0.327 0 3.0 1e-06 
0.05 0.328 0 3.0 1e-06 
3.0 0.328 0 3.0 1e-06 
0.05 0.329 0 3.0 1e-06 
3.0 0.329 0 3.0 1e-06 
0.05 0.33 0 3.0 1e-06 
3.0 0.33 0 3.0 1e-06 
0.05 0.331 0 3.0 1e-06 
3.0 0.331 0 3.0 1e-06 
0.05 0.332 0 3.0 1e-06 
3.0 0.332 0 3.0 1e-06 
0.05 0.333 0 3.0 1e-06 
3.0 0.333 0 3.0 1e-06 
0.05 0.334 0 3.0 1e-06 
3.0 0.334 0 3.0 1e-06 
0.05 0.335 0 3.0 1e-06 
3.0 0.335 0 3.0 1e-06 
0.05 0.336 0 3.0 1e-06 
3.0 0.336 0 3.0 1e-06 
0.05 0.337 0 3.0 1e-06 
3.0 0.337 0 3.0 1e-06 
0.05 0.338 0 3.0 1e-06 
3.0 0.338 0 3.0 1e-06 
0.05 0.339 0 3.0 1e-06 
3.0 0.339 0 3.0 1e-06 
0.05 0.34 0 3.0 1e-06 
3.0 0.34 0 3.0 1e-06 
0.05 0.341 0 3.0 1e-06 
3.0 0.341 0 3.0 1e-06 
0.05 0.342 0 3.0 1e-06 
3.0 0.342 0 3.0 1e-06 
0.05 0.343 0 3.0 1e-06 
3.0 0.343 0 3.0 1e-06 
0.05 0.344 0 3.0 1e-06 
3.0 0.344 0 3.0 1e-06 
0.05 0.345 0 3.0 1e-06 
3.0 0.345 0 3.0 1e-06 
0.05 0.346 0 3.0 1e-06 
3.0 0.346 0 3.0 1e-06 
0.05 0.347 0 3.0 1e-06 
3.0 0.347 0 3.0 1e-06 
0.05 0.348 0 3.0 1e-06 
3.0 0.348 0 3.0 1e-06 
0.05 0.349 0 3.0 1e-06 
3.0 0.349 0 3.0 1e-06 
0.05 0.35 0 3.0 1e-06 
3.0 0.35 0 3.0 1e-06 
0.05 0.351 0 3.0 1e-06 
3.0 0.351 0 3.0 1e-06 
0.05 0.352 0 3.0 1e-06 
3.0 0.352 0 3.0 1e-06 
0.05 0.353 0 3.0 1e-06 
3.0 0.353 0 3.0 1e-06 
0.05 0.354 0 3.0 1e-06 
3.0 0.354 0 3.0 1e-06 
0.05 0.355 0 3.0 1e-06 
3.0 0.355 0 3.0 1e-06 
0.05 0.356 0 3.0 1e-06 
3.0 0.356 0 3.0 1e-06 
0.05 0.357 0 3.0 1e-06 
3.0 0.357 0 3.0 1e-06 
0.05 0.358 0 3.0 1e-06 
3.0 0.358 0 3.0 1e-06 
0.05 0.359 0 3.0 1e-06 
3.0 0.359 0 3.0 1e-06 
0.05 0.36 0 3.0 1e-06 
3.0 0.36 0 3.0 1e-06 
0.05 0.361 0 3.0 1e-06 
3.0 0.361 0 3.0 1e-06 
0.05 0.362 0 3.0 1e-06 
3.0 0.362 0 3.0 1e-06 
0.05 0.363 0 3.0 1e-06 
3.0 0.363 0 3.0 1e-06 
0.05 0.364 0 3.0 1e-06 
3.0 0.364 0 3.0 1e-06 
0.05 0.365 0 3.0 1e-06 
3.0 0.365 0 3.0 1e-06 
0.05 0.366 0 3.0 1e-06 
3.0 0.366 0 3.0 1e-06 
0.05 0.367 0 3.0 1e-06 
3.0 0.367 0 3.0 1e-06 
0.05 0.368 0 3.0 1e-06 
3.0 0.368 0 3.0 1e-06 
0.05 0.369 0 3.0 1e-06 
3.0 0.369 0 3.0 1e-06 
0.05 0.37 0 3.0 1e-06 
3.0 0.37 0 3.0 1e-06 
0.05 0.371 0 3.0 1e-06 
3.0 0.371 0 3.0 1e-06 
0.05 0.372 0 3.0 1e-06 
3.0 0.372 0 3.0 1e-06 
0.05 0.373 0 3.0 1e-06 
3.0 0.373 0 3.0 1e-06 
0.05 0.374 0 3.0 1e-06 
3.0 0.374 0 3.0 1e-06 
0.05 0.375 0 3.0 1e-06 
3.0 0.375 0 3.0 1e-06 
0.05 0.376 0 3.0 1e-06 
3.0 0.376 0 3.0 1e-06 
0.05 0.377 0 3.0 1e-06 
3.0 0.377 0 3.0 1e-06 
0.05 0.378 0 3.0 1e-06 
3.0 0.378 0 3.0 1e-06 
0.05 0.379 0 3.0 1e-06 
3.0 0.379 0 3.0 1e-06 
0.05 0.38 0 3.0 1e-06 
3.0 0.38 0 3.0 1e-06 
0.05 0.381 0 3.0 1e-06 
3.0 0.381 0 3.0 1e-06 
0.05 0.382 0 3.0 1e-06 
3.0 0.382 0 3.0 1e-06 
0.05 0.383 0 3.0 1e-06 
3.0 0.383 0 3.0 1e-06 
0.05 0.384 0 3.0 1e-06 
3.0 0.384 0 3.0 1e-06 
0.05 0.385 0 3.0 1e-06 
3.0 0.385 0 3.0 1e-06 
0.05 0.386 0 3.0 1e-06 
3.0 0.386 0 3.0 1e-06 
0.05 0.387 0 3.0 1e-06 
3.0 0.387 0 3.0 1e-06 
0.05 0.388 0 3.0 1e-06 
3.0 0.388 0 3.0 1e-06 
0.05 0.389 0 3.0 1e-06 
3.0 0.389 0 3.0 1e-06 
0.05 0.39 0 3.0 1e-06 
3.0 0.39 0 3.0 1e-06 
0.05 0.391 0 3.0 1e-06 
3.0 0.391 0 3.0 1e-06 
0.05 0.392 0 3.0 1e-06 
3.0 0.392 0 3.0 1e-06 
0.05 0.393 0 3.0 1e-06 
3.0 0.393 0 3.0 1e-06 
0.05 0.394 0 3.0 1e-06 
3.0 0.394 0 3.0 1e-06 
0.05 0.395 0 3.0 1e-06 
3.0 0.395 0 3.0 1e-06 
0.05 0.396 0 3.0 1e-06 
3.0 0.396 0 3.0 1e-06 
0.05 0.397 0 3.0 1e-06 
3.0 0.397 0 3.0 1e-06 
0.05 0.398 0 3.0 1e-06 
3.0 0.398 0 3.0 1e-06 
0.05 0.399 0 3.0 1e-06 
3.0 0.399 0 3.0 1e-06 
0.05 0.4 0 3.0 1e-06 
3.0 0.4 0 3.0 1e-06 
0.05 0.401 0 3.0 1e-06 
3.0 0.401 0 3.0 1e-06 
0.05 0.402 0 3.0 1e-06 
3.0 0.402 0 3.0 1e-06 
0.05 0.403 0 3.0 1e-06 
3.0 0.403 0 3.0 1e-06 
0.05 0.404 0 3.0 1e-06 
3.0 0.404 0 3.0 1e-06 
0.05 0.405 0 3.0 1e-06 
3.0 0.405 0 3.0 1e-06 
0.05 0.406 0 3.0 1e-06 
3.0 0.406 0 3.0 1e-06 
0.05 0.407 0 3.0 1e-06 
3.0 0.407 0 3.0 1e-06 
0.05 0.408 0 3.0 1e-06 
3.0 0.408 0 3.0 1e-06 
0.05 0.409 0 3.0 1e-06 
3.0 0.409 0 3.0 1e-06 
0.05 0.41 0 3.0 1e-06 
3.0 0.41 0 3.0 1e-06 
0.05 0.411 0 3.0 1e-06 
3.0 0.411 0 3.0 1e-06 
0.05 0.412 0 3.0 1e-06 
3.0 0.412 0 3.0 1e-06 
0.05 0.413 0 3.0 1e-06 
3.0 0.413 0 3.0 1e-06 
0.05 0.414 0 3.0 1e-06 
3.0 0.414 0 3.0 1e-06 
0.05 0.415 0 3.0 1e-06 
3.0 0.415 0 3.0 1e-06 
0.05 0.416 0 3.0 1e-06 
3.0 0.416 0 3.0 1e-06 
0.05 0.417 0 3.0 1e-06 
3.0 0.417 0 3.0 1e-06 
0.05 0.418 0 3.0 1e-06 
3.0 0.418 0 3.0 1e-06 
0.05 0.419 0 3.0 1e-06 
3.0 0.419 0 3.0 1e-06 
0.05 0.42 0 3.0 1e-06 
3.0 0.42 0 3.0 1e-06 
0.05 0.421 0 3.0 1e-06 
3.0 0.421 0 3.0 1e-06 
0.05 0.422 0 3.0 1e-06 
3.0 0.422 0 3.0 1e-06 
0.05 0.423 0 3.0 1e-06 
3.0 0.423 0 3.0 1e-06 
0.05 0.424 0 3.0 1e-06 
3.0 0.424 0 3.0 1e-06 
0.05 0.425 0 3.0 1e-06 
3.0 0.425 0 3.0 1e-06 
0.05 0.426 0 3.0 1e-06 
3.0 0.426 0 3.0 1e-06 
0.05 0.427 0 3.0 1e-06 
3.0 0.427 0 3.0 1e-06 
0.05 0.428 0 3.0 1e-06 
3.0 0.428 0 3.0 1e-06 
0.05 0.429 0 3.0 1e-06 
3.0 0.429 0 3.0 1e-06 
0.05 0.43 0 3.0 1e-06 
3.0 0.43 0 3.0 1e-06 
0.05 0.431 0 3.0 1e-06 
3.0 0.431 0 3.0 1e-06 
0.05 0.432 0 3.0 1e-06 
3.0 0.432 0 3.0 1e-06 
0.05 0.433 0 3.0 1e-06 
3.0 0.433 0 3.0 1e-06 
0.05 0.434 0 3.0 1e-06 
3.0 0.434 0 3.0 1e-06 
0.05 0.435 0 3.0 1e-06 
3.0 0.435 0 3.0 1e-06 
0.05 0.436 0 3.0 1e-06 
3.0 0.436 0 3.0 1e-06 
0.05 0.437 0 3.0 1e-06 
3.0 0.437 0 3.0 1e-06 
0.05 0.438 0 3.0 1e-06 
3.0 0.438 0 3.0 1e-06 
0.05 0.439 0 3.0 1e-06 
3.0 0.439 0 3.0 1e-06 
0.05 0.44 0 3.0 1e-06 
3.0 0.44 0 3.0 1e-06 
0.05 0.441 0 3.0 1e-06 
3.0 0.441 0 3.0 1e-06 
0.05 0.442 0 3.0 1e-06 
3.0 0.442 0 3.0 1e-06 
0.05 0.443 0 3.0 1e-06 
3.0 0.443 0 3.0 1e-06 
0.05 0.444 0 3.0 1e-06 
3.0 0.444 0 3.0 1e-06 
0.05 0.445 0 3.0 1e-06 
3.0 0.445 0 3.0 1e-06 
0.05 0.446 0 3.0 1e-06 
3.0 0.446 0 3.0 1e-06 
0.05 0.447 0 3.0 1e-06 
3.0 0.447 0 3.0 1e-06 
0.05 0.448 0 3.0 1e-06 
3.0 0.448 0 3.0 1e-06 
0.05 0.449 0 3.0 1e-06 
3.0 0.449 0 3.0 1e-06 
0.05 0.45 0 3.0 1e-06 
3.0 0.45 0 3.0 1e-06 
0.05 0.451 0 3.0 1e-06 
3.0 0.451 0 3.0 1e-06 
0.05 0.452 0 3.0 1e-06 
3.0 0.452 0 3.0 1e-06 
0.05 0.453 0 3.0 1e-06 
3.0 0.453 0 3.0 1e-06 
0.05 0.454 0 3.0 1e-06 
3.0 0.454 0 3.0 1e-06 
0.05 0.455 0 3.0 1e-06 
3.0 0.455 0 3.0 1e-06 
0.05 0.456 0 3.0 1e-06 
3.0 0.456 0 3.0 1e-06 
0.05 0.457 0 3.0 1e-06 
3.0 0.457 0 3.0 1e-06 
0.05 0.458 0 3.0 1e-06 
3.0 0.458 0 3.0 1e-06 
0.05 0.459 0 3.0 1e-06 
3.0 0.459 0 3.0 1e-06 
0.05 0.46 0 3.0 1e-06 
3.0 0.46 0 3.0 1e-06 
0.05 0.461 0 3.0 1e-06 
3.0 0.461 0 3.0 1e-06 
0.05 0.462 0 3.0 1e-06 
3.0 0.462 0 3.0 1e-06 
0.05 0.463 0 3.0 1e-06 
3.0 0.463 0 3.0 1e-06 
0.05 0.464 0 3.0 1e-06 
3.0 0.464 0 3.0 1e-06 
0.05 0.465 0 3.0 1e-06 
3.0 0.465 0 3.0 1e-06 
0.05 0.466 0 3.0 1e-06 
3.0 0.466 0 3.0 1e-06 
0.05 0.467 0 3.0 1e-06 
3.0 0.467 0 3.0 1e-06 
0.05 0.468 0 3.0 1e-06 
3.0 0.468 0 3.0 1e-06 
0.05 0.469 0 3.0 1e-06 
3.0 0.469 0 3.0 1e-06 
0.05 0.47 0 3.0 1e-06 
3.0 0.47 0 3.0 1e-06 
0.05 0.471 0 3.0 1e-06 
3.0 0.471 0 3.0 1e-06 
0.05 0.472 0 3.0 1e-06 
3.0 0.472 0 3.0 1e-06 
0.05 0.473 0 3.0 1e-06 
3.0 0.473 0 3.0 1e-06 
0.05 0.474 0 3.0 1e-06 
3.0 0.474 0 3.0 1e-06 
0.05 0.475 0 3.0 1e-06 
3.0 0.475 0 3.0 1e-06 
0.05 0.476 0 3.0 1e-06 
3.0 0.476 0 3.0 1e-06 
0.05 0.477 0 3.0 1e-06 
3.0 0.477 0 3.0 1e-06 
0.05 0.478 0 3.0 1e-06 
3.0 0.478 0 3.0 1e-06 
0.05 0.479 0 3.0 1e-06 
3.0 0.479 0 3.0 1e-06 
0.05 0.48 0 3.0 1e-06 
3.0 0.48 0 3.0 1e-06 
0.05 0.481 0 3.0 1e-06 
3.0 0.481 0 3.0 1e-06 
0.05 0.482 0 3.0 1e-06 
3.0 0.482 0 3.0 1e-06 
0.05 0.483 0 3.0 1e-06 
3.0 0.483 0 3.0 1e-06 
0.05 0.484 0 3.0 1e-06 
3.0 0.484 0 3.0 1e-06 
0.05 0.485 0 3.0 1e-06 
3.0 0.485 0 3.0 1e-06 
0.05 0.486 0 3.0 1e-06 
3.0 0.486 0 3.0 1e-06 
0.05 0.487 0 3.0 1e-06 
3.0 0.487 0 3.0 1e-06 
0.05 0.488 0 3.0 1e-06 
3.0 0.488 0 3.0 1e-06 
0.05 0.489 0 3.0 1e-06 
3.0 0.489 0 3.0 1e-06 
0.05 0.49 0 3.0 1e-06 
3.0 0.49 0 3.0 1e-06 
0.05 0.491 0 3.0 1e-06 
3.0 0.491 0 3.0 1e-06 
0.05 0.492 0 3.0 1e-06 
3.0 0.492 0 3.0 1e-06 
0.05 0.493 0 3.0 1e-06 
3.0 0.493 0 3.0 1e-06 
0.05 0.494 0 3.0 1e-06 
3.0 0.494 0 3.0 1e-06 
0.05 0.495 0 3.0 1e-06 
3.0 0.495 0 3.0 1e-06 
0.05 0.496 0 3.0 1e-06 
3.0 0.496 0 3.0 1e-06 
0.05 0.497 0 3.0 1e-06 
3.0 0.497 0 3.0 1e-06 
0.05 0.498 0 3.0 1e-06 
3.0 0.498 0 3.0 1e-06 
0.05 0.499 0 3.0 1e-06 
3.0 0.499 0 3.0 1e-06 
0.05 0.5 0 3.0 1e-06 
3.0 0.5 0 3.0 1e-06 
0.05 0.501 0 3.0 1e-06 
3.0 0.501 0 3.0 1e-06 
0.05 0.502 0 3.0 1e-06 
3.0 0.502 0 3.0 1e-06 
0.05 0.503 0 3.0 1e-06 
3.0 0.503 0 3.0 1e-06 
0.05 0.504 0 3.0 1e-06 
3.0 0.504 0 3.0 1e-06 
0.05 0.505 0 3.0 1e-06 
3.0 0.505 0 3.0 1e-06 
0.05 0.506 0 3.0 1e-06 
3.0 0.506 0 3.0 1e-06 
0.05 0.507 0 3.0 1e-06 
3.0 0.507 0 3.0 1e-06 
0.05 0.508 0 3.0 1e-06 
3.0 0.508 0 3.0 1e-06 
0.05 0.509 0 3.0 1e-06 
3.0 0.509 0 3.0 1e-06 
0.05 0.51 0 3.0 1e-06 
3.0 0.51 0 3.0 1e-06 
0.05 0.511 0 3.0 1e-06 
3.0 0.511 0 3.0 1e-06 
0.05 0.512 0 3.0 1e-06 
3.0 0.512 0 3.0 1e-06 
0.05 0.513 0 3.0 1e-06 
3.0 0.513 0 3.0 1e-06 
0.05 0.514 0 3.0 1e-06 
3.0 0.514 0 3.0 1e-06 
0.05 0.515 0 3.0 1e-06 
3.0 0.515 0 3.0 1e-06 
0.05 0.516 0 3.0 1e-06 
3.0 0.516 0 3.0 1e-06 
0.05 0.517 0 3.0 1e-06 
3.0 0.517 0 3.0 1e-06 
0.05 0.518 0 3.0 1e-06 
3.0 0.518 0 3.0 1e-06 
0.05 0.519 0 3.0 1e-06 
3.0 0.519 0 3.0 1e-06 
0.05 0.52 0 3.0 1e-06 
3.0 0.52 0 3.0 1e-06 
0.05 0.521 0 3.0 1e-06 
3.0 0.521 0 3.0 1e-06 
0.05 0.522 0 3.0 1e-06 
3.0 0.522 0 3.0 1e-06 
0.05 0.523 0 3.0 1e-06 
3.0 0.523 0 3.0 1e-06 
0.05 0.524 0 3.0 1e-06 
3.0 0.524 0 3.0 1e-06 
0.05 0.525 0 3.0 1e-06 
3.0 0.525 0 3.0 1e-06 
0.05 0.526 0 3.0 1e-06 
3.0 0.526 0 3.0 1e-06 
0.05 0.527 0 3.0 1e-06 
3.0 0.527 0 3.0 1e-06 
0.05 0.528 0 3.0 1e-06 
3.0 0.528 0 3.0 1e-06 
0.05 0.529 0 3.0 1e-06 
3.0 0.529 0 3.0 1e-06 
0.05 0.53 0 3.0 1e-06 
3.0 0.53 0 3.0 1e-06 
0.05 0.531 0 3.0 1e-06 
3.0 0.531 0 3.0 1e-06 
0.05 0.532 0 3.0 1e-06 
3.0 0.532 0 3.0 1e-06 
0.05 0.533 0 3.0 1e-06 
3.0 0.533 0 3.0 1e-06 
0.05 0.534 0 3.0 1e-06 
3.0 0.534 0 3.0 1e-06 
0.05 0.535 0 3.0 1e-06 
3.0 0.535 0 3.0 1e-06 
0.05 0.536 0 3.0 1e-06 
3.0 0.536 0 3.0 1e-06 
0.05 0.537 0 3.0 1e-06 
3.0 0.537 0 3.0 1e-06 
0.05 0.538 0 3.0 1e-06 
3.0 0.538 0 3.0 1e-06 
0.05 0.539 0 3.0 1e-06 
3.0 0.539 0 3.0 1e-06 
0.05 0.54 0 3.0 1e-06 
3.0 0.54 0 3.0 1e-06 
0.05 0.541 0 3.0 1e-06 
3.0 0.541 0 3.0 1e-06 
0.05 0.542 0 3.0 1e-06 
3.0 0.542 0 3.0 1e-06 
0.05 0.543 0 3.0 1e-06 
3.0 0.543 0 3.0 1e-06 
0.05 0.544 0 3.0 1e-06 
3.0 0.544 0 3.0 1e-06 
0.05 0.545 0 3.0 1e-06 
3.0 0.545 0 3.0 1e-06 
0.05 0.546 0 3.0 1e-06 
3.0 0.546 0 3.0 1e-06 
0.05 0.547 0 3.0 1e-06 
3.0 0.547 0 3.0 1e-06 
0.05 0.548 0 3.0 1e-06 
3.0 0.548 0 3.0 1e-06 
0.05 0.549 0 3.0 1e-06 
3.0 0.549 0 3.0 1e-06 
0.05 0.55 0 3.0 1e-06 
3.0 0.55 0 3.0 1e-06 
0.05 0.551 0 3.0 1e-06 
3.0 0.551 0 3.0 1e-06 
0.05 0.552 0 3.0 1e-06 
3.0 0.552 0 3.0 1e-06 
0.05 0.553 0 3.0 1e-06 
3.0 0.553 0 3.0 1e-06 
0.05 0.554 0 3.0 1e-06 
3.0 0.554 0 3.0 1e-06 
0.05 0.555 0 3.0 1e-06 
3.0 0.555 0 3.0 1e-06 
0.05 0.556 0 3.0 1e-06 
3.0 0.556 0 3.0 1e-06 
0.05 0.557 0 3.0 1e-06 
3.0 0.557 0 3.0 1e-06 
0.05 0.558 0 3.0 1e-06 
3.0 0.558 0 3.0 1e-06 
0.05 0.559 0 3.0 1e-06 
3.0 0.559 0 3.0 1e-06 
0.05 0.56 0 3.0 1e-06 
3.0 0.56 0 3.0 1e-06 
0.05 0.561 0 3.0 1e-06 
3.0 0.561 0 3.0 1e-06 
0.05 0.562 0 3.0 1e-06 
3.0 0.562 0 3.0 1e-06 
0.05 0.563 0 3.0 1e-06 
3.0 0.563 0 3.0 1e-06 
0.05 0.564 0 3.0 1e-06 
3.0 0.564 0 3.0 1e-06 
0.05 0.565 0 3.0 1e-06 
3.0 0.565 0 3.0 1e-06 
0.05 0.566 0 3.0 1e-06 
3.0 0.566 0 3.0 1e-06 
0.05 0.567 0 3.0 1e-06 
3.0 0.567 0 3.0 1e-06 
0.05 0.568 0 3.0 1e-06 
3.0 0.568 0 3.0 1e-06 
0.05 0.569 0 3.0 1e-06 
3.0 0.569 0 3.0 1e-06 
0.05 0.57 0 3.0 1e-06 
3.0 0.57 0 3.0 1e-06 
0.05 0.571 0 3.0 1e-06 
3.0 0.571 0 3.0 1e-06 
0.05 0.572 0 3.0 1e-06 
3.0 0.572 0 3.0 1e-06 
0.05 0.573 0 3.0 1e-06 
3.0 0.573 0 3.0 1e-06 
0.05 0.574 0 3.0 1e-06 
3.0 0.574 0 3.0 1e-06 
0.05 0.575 0 3.0 1e-06 
3.0 0.575 0 3.0 1e-06 
0.05 0.576 0 3.0 1e-06 
3.0 0.576 0 3.0 1e-06 
0.05 0.577 0 3.0 1e-06 
3.0 0.577 0 3.0 1e-06 
0.05 0.578 0 3.0 1e-06 
3.0 0.578 0 3.0 1e-06 
0.05 0.579 0 3.0 1e-06 
3.0 0.579 0 3.0 1e-06 
0.05 0.58 0 3.0 1e-06 
3.0 0.58 0 3.0 1e-06 
0.05 0.581 0 3.0 1e-06 
3.0 0.581 0 3.0 1e-06 
0.05 0.582 0 3.0 1e-06 
3.0 0.582 0 3.0 1e-06 
0.05 0.583 0 3.0 1e-06 
3.0 0.583 0 3.0 1e-06 
0.05 0.584 0 3.0 1e-06 
3.0 0.584 0 3.0 1e-06 
0.05 0.585 0 3.0 1e-06 
3.0 0.585 0 3.0 1e-06 
0.05 0.586 0 3.0 1e-06 
3.0 0.586 0 3.0 1e-06 
0.05 0.587 0 3.0 1e-06 
3.0 0.587 0 3.0 1e-06 
0.05 0.588 0 3.0 1e-06 
3.0 0.588 0 3.0 1e-06 
0.05 0.589 0 3.0 1e-06 
3.0 0.589 0 3.0 1e-06 
0.05 0.59 0 3.0 1e-06 
3.0 0.59 0 3.0 1e-06 
0.05 0.591 0 3.0 1e-06 
3.0 0.591 0 3.0 1e-06 
0.05 0.592 0 3.0 1e-06 
3.0 0.592 0 3.0 1e-06 
0.05 0.593 0 3.0 1e-06 
3.0 0.593 0 3.0 1e-06 
0.05 0.594 0 3.0 1e-06 
3.0 0.594 0 3.0 1e-06 
0.05 0.595 0 3.0 1e-06 
3.0 0.595 0 3.0 1e-06 
0.05 0.596 0 3.0 1e-06 
3.0 0.596 0 3.0 1e-06 
0.05 0.597 0 3.0 1e-06 
3.0 0.597 0 3.0 1e-06 
0.05 0.598 0 3.0 1e-06 
3.0 0.598 0 3.0 1e-06 
0.05 0.599 0 3.0 1e-06 
3.0 0.599 0 3.0 1e-06 
0.05 0.6 0 3.0 1e-06 
3.0 0.6 0 3.0 1e-06 
0.05 0.601 0 3.0 1e-06 
3.0 0.601 0 3.0 1e-06 
0.05 0.602 0 3.0 1e-06 
3.0 0.602 0 3.0 1e-06 
0.05 0.603 0 3.0 1e-06 
3.0 0.603 0 3.0 1e-06 
0.05 0.604 0 3.0 1e-06 
3.0 0.604 0 3.0 1e-06 
0.05 0.605 0 3.0 1e-06 
3.0 0.605 0 3.0 1e-06 
0.05 0.606 0 3.0 1e-06 
3.0 0.606 0 3.0 1e-06 
0.05 0.607 0 3.0 1e-06 
3.0 0.607 0 3.0 1e-06 
0.05 0.608 0 3.0 1e-06 
3.0 0.608 0 3.0 1e-06 
0.05 0.609 0 3.0 1e-06 
3.0 0.609 0 3.0 1e-06 
0.05 0.61 0 3.0 1e-06 
3.0 0.61 0 3.0 1e-06 
0.05 0.611 0 3.0 1e-06 
3.0 0.611 0 3.0 1e-06 
0.05 0.612 0 3.0 1e-06 
3.0 0.612 0 3.0 1e-06 
0.05 0.613 0 3.0 1e-06 
3.0 0.613 0 3.0 1e-06 
0.05 0.614 0 3.0 1e-06 
3.0 0.614 0 3.0 1e-06 
0.05 0.615 0 3.0 1e-06 
3.0 0.615 0 3.0 1e-06 
0.05 0.616 0 3.0 1e-06 
3.0 0.616 0 3.0 1e-06 
0.05 0.617 0 3.0 1e-06 
3.0 0.617 0 3.0 1e-06 
0.05 0.618 0 3.0 1e-06 
3.0 0.618 0 3.0 1e-06 
0.05 0.619 0 3.0 1e-06 
3.0 0.619 0 3.0 1e-06 
0.05 0.62 0 3.0 1e-06 
3.0 0.62 0 3.0 1e-06 
0.05 0.621 0 3.0 1e-06 
3.0 0.621 0 3.0 1e-06 
0.05 0.622 0 3.0 1e-06 
3.0 0.622 0 3.0 1e-06 
0.05 0.623 0 3.0 1e-06 
3.0 0.623 0 3.0 1e-06 
0.05 0.624 0 3.0 1e-06 
3.0 0.624 0 3.0 1e-06 
0.05 0.625 0 3.0 1e-06 
3.0 0.625 0 3.0 1e-06 
0.05 0.626 0 3.0 1e-06 
3.0 0.626 0 3.0 1e-06 
0.05 0.627 0 3.0 1e-06 
3.0 0.627 0 3.0 1e-06 
0.05 0.628 0 3.0 1e-06 
3.0 0.628 0 3.0 1e-06 
0.05 0.629 0 3.0 1e-06 
3.0 0.629 0 3.0 1e-06 
0.05 0.63 0 3.0 1e-06 
3.0 0.63 0 3.0 1e-06 
0.05 0.631 0 3.0 1e-06 
3.0 0.631 0 3.0 1e-06 
0.05 0.632 0 3.0 1e-06 
3.0 0.632 0 3.0 1e-06 
0.05 0.633 0 3.0 1e-06 
3.0 0.633 0 3.0 1e-06 
0.05 0.634 0 3.0 1e-06 
3.0 0.634 0 3.0 1e-06 
0.05 0.635 0 3.0 1e-06 
3.0 0.635 0 3.0 1e-06 
0.05 0.636 0 3.0 1e-06 
3.0 0.636 0 3.0 1e-06 
0.05 0.637 0 3.0 1e-06 
3.0 0.637 0 3.0 1e-06 
0.05 0.638 0 3.0 1e-06 
3.0 0.638 0 3.0 1e-06 
0.05 0.639 0 3.0 1e-06 
3.0 0.639 0 3.0 1e-06 
0.05 0.64 0 3.0 1e-06 
3.0 0.64 0 3.0 1e-06 
0.05 0.641 0 3.0 1e-06 
3.0 0.641 0 3.0 1e-06 
0.05 0.642 0 3.0 1e-06 
3.0 0.642 0 3.0 1e-06 
0.05 0.643 0 3.0 1e-06 
3.0 0.643 0 3.0 1e-06 
0.05 0.644 0 3.0 1e-06 
3.0 0.644 0 3.0 1e-06 
0.05 0.645 0 3.0 1e-06 
3.0 0.645 0 3.0 1e-06 
0.05 0.646 0 3.0 1e-06 
3.0 0.646 0 3.0 1e-06 
0.05 0.647 0 3.0 1e-06 
3.0 0.647 0 3.0 1e-06 
0.05 0.648 0 3.0 1e-06 
3.0 0.648 0 3.0 1e-06 
0.05 0.649 0 3.0 1e-06 
3.0 0.649 0 3.0 1e-06 
0.05 0.65 0 3.0 1e-06 
3.0 0.65 0 3.0 1e-06 
0.05 0.651 0 3.0 1e-06 
3.0 0.651 0 3.0 1e-06 
0.05 0.652 0 3.0 1e-06 
3.0 0.652 0 3.0 1e-06 
0.05 0.653 0 3.0 1e-06 
3.0 0.653 0 3.0 1e-06 
0.05 0.654 0 3.0 1e-06 
3.0 0.654 0 3.0 1e-06 
0.05 0.655 0 3.0 1e-06 
3.0 0.655 0 3.0 1e-06 
0.05 0.656 0 3.0 1e-06 
3.0 0.656 0 3.0 1e-06 
0.05 0.657 0 3.0 1e-06 
3.0 0.657 0 3.0 1e-06 
0.05 0.658 0 3.0 1e-06 
3.0 0.658 0 3.0 1e-06 
0.05 0.659 0 3.0 1e-06 
3.0 0.659 0 3.0 1e-06 
0.05 0.66 0 3.0 1e-06 
3.0 0.66 0 3.0 1e-06 
0.05 0.661 0 3.0 1e-06 
3.0 0.661 0 3.0 1e-06 
0.05 0.662 0 3.0 1e-06 
3.0 0.662 0 3.0 1e-06 
0.05 0.663 0 3.0 1e-06 
3.0 0.663 0 3.0 1e-06 
0.05 0.664 0 3.0 1e-06 
3.0 0.664 0 3.0 1e-06 
0.05 0.665 0 3.0 1e-06 
3.0 0.665 0 3.0 1e-06 
0.05 0.666 0 3.0 1e-06 
3.0 0.666 0 3.0 1e-06 
0.05 0.667 0 3.0 1e-06 
3.0 0.667 0 3.0 1e-06 
0.05 0.668 0 3.0 1e-06 
3.0 0.668 0 3.0 1e-06 
0.05 0.669 0 3.0 1e-06 
3.0 0.669 0 3.0 1e-06 
0.05 0.67 0 3.0 1e-06 
3.0 0.67 0 3.0 1e-06 
0.05 0.671 0 3.0 1e-06 
3.0 0.671 0 3.0 1e-06 
0.05 0.672 0 3.0 1e-06 
3.0 0.672 0 3.0 1e-06 
0.05 0.673 0 3.0 1e-06 
3.0 0.673 0 3.0 1e-06 
0.05 0.674 0 3.0 1e-06 
3.0 0.674 0 3.0 1e-06 
0.05 0.675 0 3.0 1e-06 
3.0 0.675 0 3.0 1e-06 
0.05 0.676 0 3.0 1e-06 
3.0 0.676 0 3.0 1e-06 
0.05 0.677 0 3.0 1e-06 
3.0 0.677 0 3.0 1e-06 
0.05 0.678 0 3.0 1e-06 
3.0 0.678 0 3.0 1e-06 
0.05 0.679 0 3.0 1e-06 
3.0 0.679 0 3.0 1e-06 
0.05 0.68 0 3.0 1e-06 
3.0 0.68 0 3.0 1e-06 
0.05 0.681 0 3.0 1e-06 
3.0 0.681 0 3.0 1e-06 
0.05 0.682 0 3.0 1e-06 
3.0 0.682 0 3.0 1e-06 
0.05 0.683 0 3.0 1e-06 
3.0 0.683 0 3.0 1e-06 
0.05 0.684 0 3.0 1e-06 
3.0 0.684 0 3.0 1e-06 
0.05 0.685 0 3.0 1e-06 
3.0 0.685 0 3.0 1e-06 
0.05 0.686 0 3.0 1e-06 
3.0 0.686 0 3.0 1e-06 
0.05 0.687 0 3.0 1e-06 
3.0 0.687 0 3.0 1e-06 
0.05 0.688 0 3.0 1e-06 
3.0 0.688 0 3.0 1e-06 
0.05 0.689 0 3.0 1e-06 
3.0 0.689 0 3.0 1e-06 
0.05 0.69 0 3.0 1e-06 
3.0 0.69 0 3.0 1e-06 
0.05 0.691 0 3.0 1e-06 
3.0 0.691 0 3.0 1e-06 
0.05 0.692 0 3.0 1e-06 
3.0 0.692 0 3.0 1e-06 
0.05 0.693 0 3.0 1e-06 
3.0 0.693 0 3.0 1e-06 
0.05 0.694 0 3.0 1e-06 
3.0 0.694 0 3.0 1e-06 
0.05 0.695 0 3.0 1e-06 
3.0 0.695 0 3.0 1e-06 
0.05 0.696 0 3.0 1e-06 
3.0 0.696 0 3.0 1e-06 
0.05 0.697 0 3.0 1e-06 
3.0 0.697 0 3.0 1e-06 
0.05 0.698 0 3.0 1e-06 
3.0 0.698 0 3.0 1e-06 
0.05 0.699 0 3.0 1e-06 
3.0 0.699 0 3.0 1e-06 
0.05 0.7 0 3.0 1e-06 
3.0 0.7 0 3.0 1e-06 
0.05 0.701 0 3.0 1e-06 
3.0 0.701 0 3.0 1e-06 
0.05 0.702 0 3.0 1e-06 
3.0 0.702 0 3.0 1e-06 
0.05 0.703 0 3.0 1e-06 
3.0 0.703 0 3.0 1e-06 
0.05 0.704 0 3.0 1e-06 
3.0 0.704 0 3.0 1e-06 
0.05 0.705 0 3.0 1e-06 
3.0 0.705 0 3.0 1e-06 
0.05 0.706 0 3.0 1e-06 
3.0 0.706 0 3.0 1e-06 
0.05 0.707 0 3.0 1e-06 
3.0 0.707 0 3.0 1e-06 
0.05 0.708 0 3.0 1e-06 
3.0 0.708 0 3.0 1e-06 
0.05 0.709 0 3.0 1e-06 
3.0 0.709 0 3.0 1e-06 
0.05 0.71 0 3.0 1e-06 
3.0 0.71 0 3.0 1e-06 
0.05 0.711 0 3.0 1e-06 
3.0 0.711 0 3.0 1e-06 
0.05 0.712 0 3.0 1e-06 
3.0 0.712 0 3.0 1e-06 
0.05 0.713 0 3.0 1e-06 
3.0 0.713 0 3.0 1e-06 
0.05 0.714 0 3.0 1e-06 
3.0 0.714 0 3.0 1e-06 
0.05 0.715 0 3.0 1e-06 
3.0 0.715 0 3.0 1e-06 
0.05 0.716 0 3.0 1e-06 
3.0 0.716 0 3.0 1e-06 
0.05 0.717 0 3.0 1e-06 
3.0 0.717 0 3.0 1e-06 
0.05 0.718 0 3.0 1e-06 
3.0 0.718 0 3.0 1e-06 
0.05 0.719 0 3.0 1e-06 
3.0 0.719 0 3.0 1e-06 
0.05 0.72 0 3.0 1e-06 
3.0 0.72 0 3.0 1e-06 
0.05 0.721 0 3.0 1e-06 
3.0 0.721 0 3.0 1e-06 
0.05 0.722 0 3.0 1e-06 
3.0 0.722 0 3.0 1e-06 
0.05 0.723 0 3.0 1e-06 
3.0 0.723 0 3.0 1e-06 
0.05 0.724 0 3.0 1e-06 
3.0 0.724 0 3.0 1e-06 
0.05 0.725 0 3.0 1e-06 
3.0 0.725 0 3.0 1e-06 
0.05 0.726 0 3.0 1e-06 
3.0 0.726 0 3.0 1e-06 
0.05 0.727 0 3.0 1e-06 
3.0 0.727 0 3.0 1e-06 
0.05 0.728 0 3.0 1e-06 
3.0 0.728 0 3.0 1e-06 
0.05 0.729 0 3.0 1e-06 
3.0 0.729 0 3.0 1e-06 
0.05 0.73 0 3.0 1e-06 
3.0 0.73 0 3.0 1e-06 
0.05 0.731 0 3.0 1e-06 
3.0 0.731 0 3.0 1e-06 
0.05 0.732 0 3.0 1e-06 
3.0 0.732 0 3.0 1e-06 
0.05 0.733 0 3.0 1e-06 
3.0 0.733 0 3.0 1e-06 
0.05 0.734 0 3.0 1e-06 
3.0 0.734 0 3.0 1e-06 
0.05 0.735 0 3.0 1e-06 
3.0 0.735 0 3.0 1e-06 
0.05 0.736 0 3.0 1e-06 
3.0 0.736 0 3.0 1e-06 
0.05 0.737 0 3.0 1e-06 
3.0 0.737 0 3.0 1e-06 
0.05 0.738 0 3.0 1e-06 
3.0 0.738 0 3.0 1e-06 
0.05 0.739 0 3.0 1e-06 
3.0 0.739 0 3.0 1e-06 
0.05 0.74 0 3.0 1e-06 
3.0 0.74 0 3.0 1e-06 
0.05 0.741 0 3.0 1e-06 
3.0 0.741 0 3.0 1e-06 
0.05 0.742 0 3.0 1e-06 
3.0 0.742 0 3.0 1e-06 
0.05 0.743 0 3.0 1e-06 
3.0 0.743 0 3.0 1e-06 
0.05 0.744 0 3.0 1e-06 
3.0 0.744 0 3.0 1e-06 
0.05 0.745 0 3.0 1e-06 
3.0 0.745 0 3.0 1e-06 
0.05 0.746 0 3.0 1e-06 
3.0 0.746 0 3.0 1e-06 
0.05 0.747 0 3.0 1e-06 
3.0 0.747 0 3.0 1e-06 
0.05 0.748 0 3.0 1e-06 
3.0 0.748 0 3.0 1e-06 
0.05 0.749 0 3.0 1e-06 
3.0 0.749 0 3.0 1e-06 
0.05 0.75 0 3.0 1e-06 
3.0 0.75 0 3.0 1e-06 
0.05 0.751 0 3.0 1e-06 
3.0 0.751 0 3.0 1e-06 
0.05 0.752 0 3.0 1e-06 
3.0 0.752 0 3.0 1e-06 
0.05 0.753 0 3.0 1e-06 
3.0 0.753 0 3.0 1e-06 
0.05 0.754 0 3.0 1e-06 
3.0 0.754 0 3.0 1e-06 
0.05 0.755 0 3.0 1e-06 
3.0 0.755 0 3.0 1e-06 
0.05 0.756 0 3.0 1e-06 
3.0 0.756 0 3.0 1e-06 
0.05 0.757 0 3.0 1e-06 
3.0 0.757 0 3.0 1e-06 
0.05 0.758 0 3.0 1e-06 
3.0 0.758 0 3.0 1e-06 
0.05 0.759 0 3.0 1e-06 
3.0 0.759 0 3.0 1e-06 
0.05 0.76 0 3.0 1e-06 
3.0 0.76 0 3.0 1e-06 
0.05 0.761 0 3.0 1e-06 
3.0 0.761 0 3.0 1e-06 
0.05 0.762 0 3.0 1e-06 
3.0 0.762 0 3.0 1e-06 
0.05 0.763 0 3.0 1e-06 
3.0 0.763 0 3.0 1e-06 
0.05 0.764 0 3.0 1e-06 
3.0 0.764 0 3.0 1e-06 
0.05 0.765 0 3.0 1e-06 
3.0 0.765 0 3.0 1e-06 
0.05 0.766 0 3.0 1e-06 
3.0 0.766 0 3.0 1e-06 
0.05 0.767 0 3.0 1e-06 
3.0 0.767 0 3.0 1e-06 
0.05 0.768 0 3.0 1e-06 
3.0 0.768 0 3.0 1e-06 
0.05 0.769 0 3.0 1e-06 
3.0 0.769 0 3.0 1e-06 
0.05 0.77 0 3.0 1e-06 
3.0 0.77 0 3.0 1e-06 
0.05 0.771 0 3.0 1e-06 
3.0 0.771 0 3.0 1e-06 
0.05 0.772 0 3.0 1e-06 
3.0 0.772 0 3.0 1e-06 
0.05 0.773 0 3.0 1e-06 
3.0 0.773 0 3.0 1e-06 
0.05 0.774 0 3.0 1e-06 
3.0 0.774 0 3.0 1e-06 
0.05 0.775 0 3.0 1e-06 
3.0 0.775 0 3.0 1e-06 
0.05 0.776 0 3.0 1e-06 
3.0 0.776 0 3.0 1e-06 
0.05 0.777 0 3.0 1e-06 
3.0 0.777 0 3.0 1e-06 
0.05 0.778 0 3.0 1e-06 
3.0 0.778 0 3.0 1e-06 
0.05 0.779 0 3.0 1e-06 
3.0 0.779 0 3.0 1e-06 
0.05 0.78 0 3.0 1e-06 
3.0 0.78 0 3.0 1e-06 
0.05 0.781 0 3.0 1e-06 
3.0 0.781 0 3.0 1e-06 
0.05 0.782 0 3.0 1e-06 
3.0 0.782 0 3.0 1e-06 
0.05 0.783 0 3.0 1e-06 
3.0 0.783 0 3.0 1e-06 
0.05 0.784 0 3.0 1e-06 
3.0 0.784 0 3.0 1e-06 
0.05 0.785 0 3.0 1e-06 
3.0 0.785 0 3.0 1e-06 
0.05 0.786 0 3.0 1e-06 
3.0 0.786 0 3.0 1e-06 
0.05 0.787 0 3.0 1e-06 
3.0 0.787 0 3.0 1e-06 
0.05 0.788 0 3.0 1e-06 
3.0 0.788 0 3.0 1e-06 
0.05 0.789 0 3.0 1e-06 
3.0 0.789 0 3.0 1e-06 
0.05 0.79 0 3.0 1e-06 
3.0 0.79 0 3.0 1e-06 
0.05 0.791 0 3.0 1e-06 
3.0 0.791 0 3.0 1e-06 
0.05 0.792 0 3.0 1e-06 
3.0 0.792 0 3.0 1e-06 
0.05 0.793 0 3.0 1e-06 
3.0 0.793 0 3.0 1e-06 
0.05 0.794 0 3.0 1e-06 
3.0 0.794 0 3.0 1e-06 
0.05 0.795 0 3.0 1e-06 
3.0 0.795 0 3.0 1e-06 
0.05 0.796 0 3.0 1e-06 
3.0 0.796 0 3.0 1e-06 
0.05 0.797 0 3.0 1e-06 
3.0 0.797 0 3.0 1e-06 
0.05 0.798 0 3.0 1e-06 
3.0 0.798 0 3.0 1e-06 
0.05 0.799 0 3.0 1e-06 
3.0 0.799 0 3.0 1e-06 
0.05 0.8 0 3.0 1e-06 
3.0 0.8 0 3.0 1e-06 
0.05 0.801 0 3.0 1e-06 
3.0 0.801 0 3.0 1e-06 
0.05 0.802 0 3.0 1e-06 
3.0 0.802 0 3.0 1e-06 
0.05 0.803 0 3.0 1e-06 
3.0 0.803 0 3.0 1e-06 
0.05 0.804 0 3.0 1e-06 
3.0 0.804 0 3.0 1e-06 
0.05 0.805 0 3.0 1e-06 
3.0 0.805 0 3.0 1e-06 
0.05 0.806 0 3.0 1e-06 
3.0 0.806 0 3.0 1e-06 
0.05 0.807 0 3.0 1e-06 
3.0 0.807 0 3.0 1e-06 
0.05 0.808 0 3.0 1e-06 
3.0 0.808 0 3.0 1e-06 
0.05 0.809 0 3.0 1e-06 
3.0 0.809 0 3.0 1e-06 
0.05 0.81 0 3.0 1e-06 
3.0 0.81 0 3.0 1e-06 
0.05 0.811 0 3.0 1e-06 
3.0 0.811 0 3.0 1e-06 
0.05 0.812 0 3.0 1e-06 
3.0 0.812 0 3.0 1e-06 
0.05 0.813 0 3.0 1e-06 
3.0 0.813 0 3.0 1e-06 
0.05 0.814 0 3.0 1e-06 
3.0 0.814 0 3.0 1e-06 
0.05 0.815 0 3.0 1e-06 
3.0 0.815 0 3.0 1e-06 
0.05 0.816 0 3.0 1e-06 
3.0 0.816 0 3.0 1e-06 
0.05 0.817 0 3.0 1e-06 
3.0 0.817 0 3.0 1e-06 
0.05 0.818 0 3.0 1e-06 
3.0 0.818 0 3.0 1e-06 
0.05 0.819 0 3.0 1e-06 
3.0 0.819 0 3.0 1e-06 
0.05 0.82 0 3.0 1e-06 
3.0 0.82 0 3.0 1e-06 
0.05 0.821 0 3.0 1e-06 
3.0 0.821 0 3.0 1e-06 
0.05 0.822 0 3.0 1e-06 
3.0 0.822 0 3.0 1e-06 
0.05 0.823 0 3.0 1e-06 
3.0 0.823 0 3.0 1e-06 
0.05 0.824 0 3.0 1e-06 
3.0 0.824 0 3.0 1e-06 
0.05 0.825 0 3.0 1e-06 
3.0 0.825 0 3.0 1e-06 
0.05 0.826 0 3.0 1e-06 
3.0 0.826 0 3.0 1e-06 
0.05 0.827 0 3.0 1e-06 
3.0 0.827 0 3.0 1e-06 
0.05 0.828 0 3.0 1e-06 
3.0 0.828 0 3.0 1e-06 
0.05 0.829 0 3.0 1e-06 
3.0 0.829 0 3.0 1e-06 
0.05 0.83 0 3.0 1e-06 
3.0 0.83 0 3.0 1e-06 
0.05 0.831 0 3.0 1e-06 
3.0 0.831 0 3.0 1e-06 
0.05 0.832 0 3.0 1e-06 
3.0 0.832 0 3.0 1e-06 
0.05 0.833 0 3.0 1e-06 
3.0 0.833 0 3.0 1e-06 
0.05 0.834 0 3.0 1e-06 
3.0 0.834 0 3.0 1e-06 
0.05 0.835 0 3.0 1e-06 
3.0 0.835 0 3.0 1e-06 
0.05 0.836 0 3.0 1e-06 
3.0 0.836 0 3.0 1e-06 
0.05 0.837 0 3.0 1e-06 
3.0 0.837 0 3.0 1e-06 
0.05 0.838 0 3.0 1e-06 
3.0 0.838 0 3.0 1e-06 
0.05 0.839 0 3.0 1e-06 
3.0 0.839 0 3.0 1e-06 
0.05 0.84 0 3.0 1e-06 
3.0 0.84 0 3.0 1e-06 
0.05 0.841 0 3.0 1e-06 
3.0 0.841 0 3.0 1e-06 
0.05 0.842 0 3.0 1e-06 
3.0 0.842 0 3.0 1e-06 
0.05 0.843 0 3.0 1e-06 
3.0 0.843 0 3.0 1e-06 
0.05 0.844 0 3.0 1e-06 
3.0 0.844 0 3.0 1e-06 
0.05 0.845 0 3.0 1e-06 
3.0 0.845 0 3.0 1e-06 
0.05 0.846 0 3.0 1e-06 
3.0 0.846 0 3.0 1e-06 
0.05 0.847 0 3.0 1e-06 
3.0 0.847 0 3.0 1e-06 
0.05 0.848 0 3.0 1e-06 
3.0 0.848 0 3.0 1e-06 
0.05 0.849 0 3.0 1e-06 
3.0 0.849 0 3.0 1e-06 
0.05 0.85 0 3.0 1e-06 
3.0 0.85 0 3.0 1e-06 
0.05 0.851 0 3.0 1e-06 
3.0 0.851 0 3.0 1e-06 
0.05 0.852 0 3.0 1e-06 
3.0 0.852 0 3.0 1e-06 
0.05 0.853 0 3.0 1e-06 
3.0 0.853 0 3.0 1e-06 
0.05 0.854 0 3.0 1e-06 
3.0 0.854 0 3.0 1e-06 
0.05 0.855 0 3.0 1e-06 
3.0 0.855 0 3.0 1e-06 
0.05 0.856 0 3.0 1e-06 
3.0 0.856 0 3.0 1e-06 
0.05 0.857 0 3.0 1e-06 
3.0 0.857 0 3.0 1e-06 
0.05 0.858 0 3.0 1e-06 
3.0 0.858 0 3.0 1e-06 
0.05 0.859 0 3.0 1e-06 
3.0 0.859 0 3.0 1e-06 
0.05 0.86 0 3.0 1e-06 
3.0 0.86 0 3.0 1e-06 
0.05 0.861 0 3.0 1e-06 
3.0 0.861 0 3.0 1e-06 
0.05 0.862 0 3.0 1e-06 
3.0 0.862 0 3.0 1e-06 
0.05 0.863 0 3.0 1e-06 
3.0 0.863 0 3.0 1e-06 
0.05 0.864 0 3.0 1e-06 
3.0 0.864 0 3.0 1e-06 
0.05 0.865 0 3.0 1e-06 
3.0 0.865 0 3.0 1e-06 
0.05 0.866 0 3.0 1e-06 
3.0 0.866 0 3.0 1e-06 
0.05 0.867 0 3.0 1e-06 
3.0 0.867 0 3.0 1e-06 
0.05 0.868 0 3.0 1e-06 
3.0 0.868 0 3.0 1e-06 
0.05 0.869 0 3.0 1e-06 
3.0 0.869 0 3.0 1e-06 
0.05 0.87 0 3.0 1e-06 
3.0 0.87 0 3.0 1e-06 
0.05 0.871 0 3.0 1e-06 
3.0 0.871 0 3.0 1e-06 
0.05 0.872 0 3.0 1e-06 
3.0 0.872 0 3.0 1e-06 
0.05 0.873 0 3.0 1e-06 
3.0 0.873 0 3.0 1e-06 
0.05 0.874 0 3.0 1e-06 
3.0 0.874 0 3.0 1e-06 
0.05 0.875 0 3.0 1e-06 
3.0 0.875 0 3.0 1e-06 
0.05 0.876 0 3.0 1e-06 
3.0 0.876 0 3.0 1e-06 
0.05 0.877 0 3.0 1e-06 
3.0 0.877 0 3.0 1e-06 
0.05 0.878 0 3.0 1e-06 
3.0 0.878 0 3.0 1e-06 
0.05 0.879 0 3.0 1e-06 
3.0 0.879 0 3.0 1e-06 
0.05 0.88 0 3.0 1e-06 
3.0 0.88 0 3.0 1e-06 
0.05 0.881 0 3.0 1e-06 
3.0 0.881 0 3.0 1e-06 
0.05 0.882 0 3.0 1e-06 
3.0 0.882 0 3.0 1e-06 
0.05 0.883 0 3.0 1e-06 
3.0 0.883 0 3.0 1e-06 
0.05 0.884 0 3.0 1e-06 
3.0 0.884 0 3.0 1e-06 
0.05 0.885 0 3.0 1e-06 
3.0 0.885 0 3.0 1e-06 
0.05 0.886 0 3.0 1e-06 
3.0 0.886 0 3.0 1e-06 
0.05 0.887 0 3.0 1e-06 
3.0 0.887 0 3.0 1e-06 
0.05 0.888 0 3.0 1e-06 
3.0 0.888 0 3.0 1e-06 
0.05 0.889 0 3.0 1e-06 
3.0 0.889 0 3.0 1e-06 
0.05 0.89 0 3.0 1e-06 
3.0 0.89 0 3.0 1e-06 
0.05 0.891 0 3.0 1e-06 
3.0 0.891 0 3.0 1e-06 
0.05 0.892 0 3.0 1e-06 
3.0 0.892 0 3.0 1e-06 
0.05 0.893 0 3.0 1e-06 
3.0 0.893 0 3.0 1e-06 
0.05 0.894 0 3.0 1e-06 
3.0 0.894 0 3.0 1e-06 
0.05 0.895 0 3.0 1e-06 
3.0 0.895 0 3.0 1e-06 
0.05 0.896 0 3.0 1e-06 
3.0 0.896 0 3.0 1e-06 
0.05 0.897 0 3.0 1e-06 
3.0 0.897 0 3.0 1e-06 
0.05 0.898 0 3.0 1e-06 
3.0 0.898 0 3.0 1e-06 
0.05 0.899 0 3.0 1e-06 
3.0 0.899 0 3.0 1e-06 
0.05 0.9 0 3.0 1e-06 
3.0 0.9 0 3.0 1e-06 
0.05 0.901 0 3.0 1e-06 
3.0 0.901 0 3.0 1e-06 
0.05 0.902 0 3.0 1e-06 
3.0 0.902 0 3.0 1e-06 
0.05 0.903 0 3.0 1e-06 
3.0 0.903 0 3.0 1e-06 
0.05 0.904 0 3.0 1e-06 
3.0 0.904 0 3.0 1e-06 
0.05 0.905 0 3.0 1e-06 
3.0 0.905 0 3.0 1e-06 
0.05 0.906 0 3.0 1e-06 
3.0 0.906 0 3.0 1e-06 
0.05 0.907 0 3.0 1e-06 
3.0 0.907 0 3.0 1e-06 
0.05 0.908 0 3.0 1e-06 
3.0 0.908 0 3.0 1e-06 
0.05 0.909 0 3.0 1e-06 
3.0 0.909 0 3.0 1e-06 
0.05 0.91 0 3.0 1e-06 
3.0 0.91 0 3.0 1e-06 
0.05 0.911 0 3.0 1e-06 
3.0 0.911 0 3.0 1e-06 
0.05 0.912 0 3.0 1e-06 
3.0 0.912 0 3.0 1e-06 
0.05 0.913 0 3.0 1e-06 
3.0 0.913 0 3.0 1e-06 
0.05 0.914 0 3.0 1e-06 
3.0 0.914 0 3.0 1e-06 
0.05 0.915 0 3.0 1e-06 
3.0 0.915 0 3.0 1e-06 
0.05 0.916 0 3.0 1e-06 
3.0 0.916 0 3.0 1e-06 
0.05 0.917 0 3.0 1e-06 
3.0 0.917 0 3.0 1e-06 
0.05 0.918 0 3.0 1e-06 
3.0 0.918 0 3.0 1e-06 
0.05 0.919 0 3.0 1e-06 
3.0 0.919 0 3.0 1e-06 
0.05 0.92 0 3.0 1e-06 
3.0 0.92 0 3.0 1e-06 
0.05 0.921 0 3.0 1e-06 
3.0 0.921 0 3.0 1e-06 
0.05 0.922 0 3.0 1e-06 
3.0 0.922 0 3.0 1e-06 
0.05 0.923 0 3.0 1e-06 
3.0 0.923 0 3.0 1e-06 
0.05 0.924 0 3.0 1e-06 
3.0 0.924 0 3.0 1e-06 
0.05 0.925 0 3.0 1e-06 
3.0 0.925 0 3.0 1e-06 
0.05 0.926 0 3.0 1e-06 
3.0 0.926 0 3.0 1e-06 
0.05 0.927 0 3.0 1e-06 
3.0 0.927 0 3.0 1e-06 
0.05 0.928 0 3.0 1e-06 
3.0 0.928 0 3.0 1e-06 
0.05 0.929 0 3.0 1e-06 
3.0 0.929 0 3.0 1e-06 
0.05 0.93 0 3.0 1e-06 
3.0 0.93 0 3.0 1e-06 
0.05 0.931 0 3.0 1e-06 
3.0 0.931 0 3.0 1e-06 
0.05 0.932 0 3.0 1e-06 
3.0 0.932 0 3.0 1e-06 
0.05 0.933 0 3.0 1e-06 
3.0 0.933 0 3.0 1e-06 
0.05 0.934 0 3.0 1e-06 
3.0 0.934 0 3.0 1e-06 
0.05 0.935 0 3.0 1e-06 
3.0 0.935 0 3.0 1e-06 
0.05 0.936 0 3.0 1e-06 
3.0 0.936 0 3.0 1e-06 
0.05 0.937 0 3.0 1e-06 
3.0 0.937 0 3.0 1e-06 
0.05 0.938 0 3.0 1e-06 
3.0 0.938 0 3.0 1e-06 
0.05 0.939 0 3.0 1e-06 
3.0 0.939 0 3.0 1e-06 
0.05 0.94 0 3.0 1e-06 
3.0 0.94 0 3.0 1e-06 
0.05 0.941 0 3.0 1e-06 
3.0 0.941 0 3.0 1e-06 
0.05 0.942 0 3.0 1e-06 
3.0 0.942 0 3.0 1e-06 
0.05 0.943 0 3.0 1e-06 
3.0 0.943 0 3.0 1e-06 
0.05 0.944 0 3.0 1e-06 
3.0 0.944 0 3.0 1e-06 
0.05 0.945 0 3.0 1e-06 
3.0 0.945 0 3.0 1e-06 
0.05 0.946 0 3.0 1e-06 
3.0 0.946 0 3.0 1e-06 
0.05 0.947 0 3.0 1e-06 
3.0 0.947 0 3.0 1e-06 
0.05 0.948 0 3.0 1e-06 
3.0 0.948 0 3.0 1e-06 
0.05 0.949 0 3.0 1e-06 
3.0 0.949 0 3.0 1e-06 
0.05 0.95 0 3.0 1e-06 
3.0 0.95 0 3.0 1e-06 
0.05 0.951 0 3.0 1e-06 
3.0 0.951 0 3.0 1e-06 
0.05 0.952 0 3.0 1e-06 
3.0 0.952 0 3.0 1e-06 
0.05 0.953 0 3.0 1e-06 
3.0 0.953 0 3.0 1e-06 
0.05 0.954 0 3.0 1e-06 
3.0 0.954 0 3.0 1e-06 
0.05 0.955 0 3.0 1e-06 
3.0 0.955 0 3.0 1e-06 
0.05 0.956 0 3.0 1e-06 
3.0 0.956 0 3.0 1e-06 
0.05 0.957 0 3.0 1e-06 
3.0 0.957 0 3.0 1e-06 
0.05 0.958 0 3.0 1e-06 
3.0 0.958 0 3.0 1e-06 
0.05 0.959 0 3.0 1e-06 
3.0 0.959 0 3.0 1e-06 
0.05 0.96 0 3.0 1e-06 
3.0 0.96 0 3.0 1e-06 
0.05 0.961 0 3.0 1e-06 
3.0 0.961 0 3.0 1e-06 
0.05 0.962 0 3.0 1e-06 
3.0 0.962 0 3.0 1e-06 
0.05 0.963 0 3.0 1e-06 
3.0 0.963 0 3.0 1e-06 
0.05 0.964 0 3.0 1e-06 
3.0 0.964 0 3.0 1e-06 
0.05 0.965 0 3.0 1e-06 
3.0 0.965 0 3.0 1e-06 
0.05 0.966 0 3.0 1e-06 
3.0 0.966 0 3.0 1e-06 
0.05 0.967 0 3.0 1e-06 
3.0 0.967 0 3.0 1e-06 
0.05 0.968 0 3.0 1e-06 
3.0 0.968 0 3.0 1e-06 
0.05 0.969 0 3.0 1e-06 
3.0 0.969 0 3.0 1e-06 
0.05 0.97 0 3.0 1e-06 
3.0 0.97 0 3.0 1e-06 
0.05 0.971 0 3.0 1e-06 
3.0 0.971 0 3.0 1e-06 
0.05 0.972 0 3.0 1e-06 
3.0 0.972 0 3.0 1e-06 
0.05 0.973 0 3.0 1e-06 
3.0 0.973 0 3.0 1e-06 
0.05 0.974 0 3.0 1e-06 
3.0 0.974 0 3.0 1e-06 
0.05 0.975 0 3.0 1e-06 
3.0 0.975 0 3.0 1e-06 
0.05 0.976 0 3.0 1e-06 
3.0 0.976 0 3.0 1e-06 
0.05 0.977 0 3.0 1e-06 
3.0 0.977 0 3.0 1e-06 
0.05 0.978 0 3.0 1e-06 
3.0 0.978 0 3.0 1e-06 
0.05 0.979 0 3.0 1e-06 
3.0 0.979 0 3.0 1e-06 
0.05 0.98 0 3.0 1e-06 
3.0 0.98 0 3.0 1e-06 
0.05 0.981 0 3.0 1e-06 
3.0 0.981 0 3.0 1e-06 
0.05 0.982 0 3.0 1e-06 
3.0 0.982 0 3.0 1e-06 
0.05 0.983 0 3.0 1e-06 
3.0 0.983 0 3.0 1e-06 
0.05 0.984 0 3.0 1e-06 
3.0 0.984 0 3.0 1e-06 
0.05 0.985 0 3.0 1e-06 
3.0 0.985 0 3.0 1e-06 
0.05 0.986 0 3.0 1e-06 
3.0 0.986 0 3.0 1e-06 
0.05 0.987 0 3.0 1e-06 
3.0 0.987 0 3.0 1e-06 
0.05 0.988 0 3.0 1e-06 
3.0 0.988 0 3.0 1e-06 
0.05 0.989 0 3.0 1e-06 
3.0 0.989 0 3.0 1e-06 
0.05 0.99 0 3.0 1e-06 
3.0 0.99 0 3.0 1e-06 
0.05 0.991 0 3.0 1e-06 
3.0 0.991 0 3.0 1e-06 
0.05 0.992 0 3.0 1e-06 
3.0 0.992 0 3.0 1e-06 
0.05 0.993 0 3.0 1e-06 
3.0 0.993 0 3.0 1e-06 
0.05 0.994 0 3.0 1e-06 
3.0 0.994 0 3.0 1e-06 
0.05 0.995 0 3.0 1e-06 
3.0 0.995 0 3.0 1e-06 
0.05 0.996 0 3.0 1e-06 
3.0 0.996 0 3.0 1e-06 
0.05 0.997 0 3.0 1e-06 
3.0 0.997 0 3.0 1e-06 
0.05 0.998 0 3.0 1e-06 
3.0 0.998 0 3.0 1e-06 
0.05 0.999 0 3.0 1e-06 
3.0 0.999 0 3.0 1e-06 
0.05 1.0 0 3.0 1e-06 
3.0 1.0 0 3.0 1e-06 
0.05 1.001 0 3.0 1e-06 
3.0 1.001 0 3.0 1e-06 
0.05 1.002 0 3.0 1e-06 
3.0 1.002 0 3.0 1e-06 
0.05 1.003 0 3.0 1e-06 
3.0 1.003 0 3.0 1e-06 
0.05 1.004 0 3.0 1e-06 
3.0 1.004 0 3.0 1e-06 
0.05 1.005 0 3.0 1e-06 
3.0 1.005 0 3.0 1e-06 
0.05 1.006 0 3.0 1e-06 
3.0 1.006 0 3.0 1e-06 
0.05 1.007 0 3.0 1e-06 
3.0 1.007 0 3.0 1e-06 
0.05 1.008 0 3.0 1e-06 
3.0 1.008 0 3.0 1e-06 
0.05 1.009 0 3.0 1e-06 
3.0 1.009 0 3.0 1e-06 
0.05 1.01 0 3.0 1e-06 
3.0 1.01 0 3.0 1e-06 
0.05 1.011 0 3.0 1e-06 
3.0 1.011 0 3.0 1e-06 
0.05 1.012 0 3.0 1e-06 
3.0 1.012 0 3.0 1e-06 
0.05 1.013 0 3.0 1e-06 
3.0 1.013 0 3.0 1e-06 
0.05 1.014 0 3.0 1e-06 
3.0 1.014 0 3.0 1e-06 
0.05 1.015 0 3.0 1e-06 
3.0 1.015 0 3.0 1e-06 
0.05 1.016 0 3.0 1e-06 
3.0 1.016 0 3.0 1e-06 
0.05 1.017 0 3.0 1e-06 
3.0 1.017 0 3.0 1e-06 
0.05 1.018 0 3.0 1e-06 
3.0 1.018 0 3.0 1e-06 
0.05 1.019 0 3.0 1e-06 
3.0 1.019 0 3.0 1e-06 
0.05 1.02 0 3.0 1e-06 
3.0 1.02 0 3.0 1e-06 
0.05 1.021 0 3.0 1e-06 
3.0 1.021 0 3.0 1e-06 
0.05 1.022 0 3.0 1e-06 
3.0 1.022 0 3.0 1e-06 
0.05 1.023 0 3.0 1e-06 
3.0 1.023 0 3.0 1e-06 
0.05 1.024 0 3.0 1e-06 
3.0 1.024 0 3.0 1e-06 
0.05 1.025 0 3.0 1e-06 
3.0 1.025 0 3.0 1e-06 
0.05 1.026 0 3.0 1e-06 
3.0 1.026 0 3.0 1e-06 
0.05 1.027 0 3.0 1e-06 
3.0 1.027 0 3.0 1e-06 
0.05 1.028 0 3.0 1e-06 
3.0 1.028 0 3.0 1e-06 
0.05 1.029 0 3.0 1e-06 
3.0 1.029 0 3.0 1e-06 
0.05 1.03 0 3.0 1e-06 
3.0 1.03 0 3.0 1e-06 
0.05 1.031 0 3.0 1e-06 
3.0 1.031 0 3.0 1e-06 
0.05 1.032 0 3.0 1e-06 
3.0 1.032 0 3.0 1e-06 
0.05 1.033 0 3.0 1e-06 
3.0 1.033 0 3.0 1e-06 
0.05 1.034 0 3.0 1e-06 
3.0 1.034 0 3.0 1e-06 
0.05 1.035 0 3.0 1e-06 
3.0 1.035 0 3.0 1e-06 
0.05 1.036 0 3.0 1e-06 
3.0 1.036 0 3.0 1e-06 
0.05 1.037 0 3.0 1e-06 
3.0 1.037 0 3.0 1e-06 
0.05 1.038 0 3.0 1e-06 
3.0 1.038 0 3.0 1e-06 
0.05 1.039 0 3.0 1e-06 
3.0 1.039 0 3.0 1e-06 
0.05 1.04 0 3.0 1e-06 
3.0 1.04 0 3.0 1e-06 
0.05 1.041 0 3.0 1e-06 
3.0 1.041 0 3.0 1e-06 
0.05 1.042 0 3.0 1e-06 
3.0 1.042 0 3.0 1e-06 
0.05 1.043 0 3.0 1e-06 
3.0 1.043 0 3.0 1e-06 
0.05 1.044 0 3.0 1e-06 
3.0 1.044 0 3.0 1e-06 
0.05 1.045 0 3.0 1e-06 
3.0 1.045 0 3.0 1e-06 
0.05 1.046 0 3.0 1e-06 
3.0 1.046 0 3.0 1e-06 
0.05 1.047 0 3.0 1e-06 
3.0 1.047 0 3.0 1e-06 
0.05 1.048 0 3.0 1e-06 
3.0 1.048 0 3.0 1e-06 
0.05 1.049 0 3.0 1e-06 
3.0 1.049 0 3.0 1e-06 
0.05 1.05 0 3.0 1e-06 
3.0 1.05 0 3.0 1e-06 
0.05 1.051 0 3.0 1e-06 
3.0 1.051 0 3.0 1e-06 
0.05 1.052 0 3.0 1e-06 
3.0 1.052 0 3.0 1e-06 
0.05 1.053 0 3.0 1e-06 
3.0 1.053 0 3.0 1e-06 
0.05 1.054 0 3.0 1e-06 
3.0 1.054 0 3.0 1e-06 
0.05 1.055 0 3.0 1e-06 
3.0 1.055 0 3.0 1e-06 
0.05 1.056 0 3.0 1e-06 
3.0 1.056 0 3.0 1e-06 
0.05 1.057 0 3.0 1e-06 
3.0 1.057 0 3.0 1e-06 
0.05 1.058 0 3.0 1e-06 
3.0 1.058 0 3.0 1e-06 
0.05 1.059 0 3.0 1e-06 
3.0 1.059 0 3.0 1e-06 
0.05 1.06 0 3.0 1e-06 
3.0 1.06 0 3.0 1e-06 
0.05 1.061 0 3.0 1e-06 
3.0 1.061 0 3.0 1e-06 
0.05 1.062 0 3.0 1e-06 
3.0 1.062 0 3.0 1e-06 
0.05 1.063 0 3.0 1e-06 
3.0 1.063 0 3.0 1e-06 
0.05 1.064 0 3.0 1e-06 
3.0 1.064 0 3.0 1e-06 
0.05 1.065 0 3.0 1e-06 
3.0 1.065 0 3.0 1e-06 
0.05 1.066 0 3.0 1e-06 
3.0 1.066 0 3.0 1e-06 
0.05 1.067 0 3.0 1e-06 
3.0 1.067 0 3.0 1e-06 
0.05 1.068 0 3.0 1e-06 
3.0 1.068 0 3.0 1e-06 
0.05 1.069 0 3.0 1e-06 
3.0 1.069 0 3.0 1e-06 
0.05 1.07 0 3.0 1e-06 
3.0 1.07 0 3.0 1e-06 
0.05 1.071 0 3.0 1e-06 
3.0 1.071 0 3.0 1e-06 
0.05 1.072 0 3.0 1e-06 
3.0 1.072 0 3.0 1e-06 
0.05 1.073 0 3.0 1e-06 
3.0 1.073 0 3.0 1e-06 
0.05 1.074 0 3.0 1e-06 
3.0 1.074 0 3.0 1e-06 
0.05 1.075 0 3.0 1e-06 
3.0 1.075 0 3.0 1e-06 
0.05 1.076 0 3.0 1e-06 
3.0 1.076 0 3.0 1e-06 
0.05 1.077 0 3.0 1e-06 
3.0 1.077 0 3.0 1e-06 
0.05 1.078 0 3.0 1e-06 
3.0 1.078 0 3.0 1e-06 
0.05 1.079 0 3.0 1e-06 
3.0 1.079 0 3.0 1e-06 
0.05 1.08 0 3.0 1e-06 
3.0 1.08 0 3.0 1e-06 
0.05 1.081 0 3.0 1e-06 
3.0 1.081 0 3.0 1e-06 
0.05 1.082 0 3.0 1e-06 
3.0 1.082 0 3.0 1e-06 
0.05 1.083 0 3.0 1e-06 
3.0 1.083 0 3.0 1e-06 
0.05 1.084 0 3.0 1e-06 
3.0 1.084 0 3.0 1e-06 
0.05 1.085 0 3.0 1e-06 
3.0 1.085 0 3.0 1e-06 
0.05 1.086 0 3.0 1e-06 
3.0 1.086 0 3.0 1e-06 
0.05 1.087 0 3.0 1e-06 
3.0 1.087 0 3.0 1e-06 
0.05 1.088 0 3.0 1e-06 
3.0 1.088 0 3.0 1e-06 
0.05 1.089 0 3.0 1e-06 
3.0 1.089 0 3.0 1e-06 
0.05 1.09 0 3.0 1e-06 
3.0 1.09 0 3.0 1e-06 
0.05 1.091 0 3.0 1e-06 
3.0 1.091 0 3.0 1e-06 
0.05 1.092 0 3.0 1e-06 
3.0 1.092 0 3.0 1e-06 
0.05 1.093 0 3.0 1e-06 
3.0 1.093 0 3.0 1e-06 
0.05 1.094 0 3.0 1e-06 
3.0 1.094 0 3.0 1e-06 
0.05 1.095 0 3.0 1e-06 
3.0 1.095 0 3.0 1e-06 
0.05 1.096 0 3.0 1e-06 
3.0 1.096 0 3.0 1e-06 
0.05 1.097 0 3.0 1e-06 
3.0 1.097 0 3.0 1e-06 
0.05 1.098 0 3.0 1e-06 
3.0 1.098 0 3.0 1e-06 
0.05 1.099 0 3.0 1e-06 
3.0 1.099 0 3.0 1e-06 
0.05 1.1 0 3.0 1e-06 
3.0 1.1 0 3.0 1e-06 
0.05 1.101 0 3.0 1e-06 
3.0 1.101 0 3.0 1e-06 
0.05 1.102 0 3.0 1e-06 
3.0 1.102 0 3.0 1e-06 
0.05 1.103 0 3.0 1e-06 
3.0 1.103 0 3.0 1e-06 
0.05 1.104 0 3.0 1e-06 
3.0 1.104 0 3.0 1e-06 
0.05 1.105 0 3.0 1e-06 
3.0 1.105 0 3.0 1e-06 
0.05 1.106 0 3.0 1e-06 
3.0 1.106 0 3.0 1e-06 
0.05 1.107 0 3.0 1e-06 
3.0 1.107 0 3.0 1e-06 
0.05 1.108 0 3.0 1e-06 
3.0 1.108 0 3.0 1e-06 
0.05 1.109 0 3.0 1e-06 
3.0 1.109 0 3.0 1e-06 
0.05 1.11 0 3.0 1e-06 
3.0 1.11 0 3.0 1e-06 
0.05 1.111 0 3.0 1e-06 
3.0 1.111 0 3.0 1e-06 
0.05 1.112 0 3.0 1e-06 
3.0 1.112 0 3.0 1e-06 
0.05 1.113 0 3.0 1e-06 
3.0 1.113 0 3.0 1e-06 
0.05 1.114 0 3.0 1e-06 
3.0 1.114 0 3.0 1e-06 
0.05 1.115 0 3.0 1e-06 
3.0 1.115 0 3.0 1e-06 
0.05 1.116 0 3.0 1e-06 
3.0 1.116 0 3.0 1e-06 
0.05 1.117 0 3.0 1e-06 
3.0 1.117 0 3.0 1e-06 
0.05 1.118 0 3.0 1e-06 
3.0 1.118 0 3.0 1e-06 
0.05 1.119 0 3.0 1e-06 
3.0 1.119 0 3.0 1e-06 
0.05 1.12 0 3.0 1e-06 
3.0 1.12 0 3.0 1e-06 
0.05 1.121 0 3.0 1e-06 
3.0 1.121 0 3.0 1e-06 
0.05 1.122 0 3.0 1e-06 
3.0 1.122 0 3.0 1e-06 
0.05 1.123 0 3.0 1e-06 
3.0 1.123 0 3.0 1e-06 
0.05 1.124 0 3.0 1e-06 
3.0 1.124 0 3.0 1e-06 
0.05 1.125 0 3.0 1e-06 
3.0 1.125 0 3.0 1e-06 
0.05 1.126 0 3.0 1e-06 
3.0 1.126 0 3.0 1e-06 
0.05 1.127 0 3.0 1e-06 
3.0 1.127 0 3.0 1e-06 
0.05 1.128 0 3.0 1e-06 
3.0 1.128 0 3.0 1e-06 
0.05 1.129 0 3.0 1e-06 
3.0 1.129 0 3.0 1e-06 
0.05 1.13 0 3.0 1e-06 
3.0 1.13 0 3.0 1e-06 
0.05 1.131 0 3.0 1e-06 
3.0 1.131 0 3.0 1e-06 
0.05 1.132 0 3.0 1e-06 
3.0 1.132 0 3.0 1e-06 
0.05 1.133 0 3.0 1e-06 
3.0 1.133 0 3.0 1e-06 
0.05 1.134 0 3.0 1e-06 
3.0 1.134 0 3.0 1e-06 
0.05 1.135 0 3.0 1e-06 
3.0 1.135 0 3.0 1e-06 
0.05 1.136 0 3.0 1e-06 
3.0 1.136 0 3.0 1e-06 
0.05 1.137 0 3.0 1e-06 
3.0 1.137 0 3.0 1e-06 
0.05 1.138 0 3.0 1e-06 
3.0 1.138 0 3.0 1e-06 
0.05 1.139 0 3.0 1e-06 
3.0 1.139 0 3.0 1e-06 
0.05 1.14 0 3.0 1e-06 
3.0 1.14 0 3.0 1e-06 
0.05 1.141 0 3.0 1e-06 
3.0 1.141 0 3.0 1e-06 
0.05 1.142 0 3.0 1e-06 
3.0 1.142 0 3.0 1e-06 
0.05 1.143 0 3.0 1e-06 
3.0 1.143 0 3.0 1e-06 
0.05 1.144 0 3.0 1e-06 
3.0 1.144 0 3.0 1e-06 
0.05 1.145 0 3.0 1e-06 
3.0 1.145 0 3.0 1e-06 
0.05 1.146 0 3.0 1e-06 
3.0 1.146 0 3.0 1e-06 
0.05 1.147 0 3.0 1e-06 
3.0 1.147 0 3.0 1e-06 
0.05 1.148 0 3.0 1e-06 
3.0 1.148 0 3.0 1e-06 
0.05 1.149 0 3.0 1e-06 
3.0 1.149 0 3.0 1e-06 
0.05 1.15 0 3.0 1e-06 
3.0 1.15 0 3.0 1e-06 
0.05 1.151 0 3.0 1e-06 
3.0 1.151 0 3.0 1e-06 
0.05 1.152 0 3.0 1e-06 
3.0 1.152 0 3.0 1e-06 
0.05 1.153 0 3.0 1e-06 
3.0 1.153 0 3.0 1e-06 
0.05 1.154 0 3.0 1e-06 
3.0 1.154 0 3.0 1e-06 
0.05 1.155 0 3.0 1e-06 
3.0 1.155 0 3.0 1e-06 
0.05 1.156 0 3.0 1e-06 
3.0 1.156 0 3.0 1e-06 
0.05 1.157 0 3.0 1e-06 
3.0 1.157 0 3.0 1e-06 
0.05 1.158 0 3.0 1e-06 
3.0 1.158 0 3.0 1e-06 
0.05 1.159 0 3.0 1e-06 
3.0 1.159 0 3.0 1e-06 
0.05 1.16 0 3.0 1e-06 
3.0 1.16 0 3.0 1e-06 
0.05 1.161 0 3.0 1e-06 
3.0 1.161 0 3.0 1e-06 
0.05 1.162 0 3.0 1e-06 
3.0 1.162 0 3.0 1e-06 
0.05 1.163 0 3.0 1e-06 
3.0 1.163 0 3.0 1e-06 
0.05 1.164 0 3.0 1e-06 
3.0 1.164 0 3.0 1e-06 
0.05 1.165 0 3.0 1e-06 
3.0 1.165 0 3.0 1e-06 
0.05 1.166 0 3.0 1e-06 
3.0 1.166 0 3.0 1e-06 
0.05 1.167 0 3.0 1e-06 
3.0 1.167 0 3.0 1e-06 
0.05 1.168 0 3.0 1e-06 
3.0 1.168 0 3.0 1e-06 
0.05 1.169 0 3.0 1e-06 
3.0 1.169 0 3.0 1e-06 
0.05 1.17 0 3.0 1e-06 
3.0 1.17 0 3.0 1e-06 
0.05 1.171 0 3.0 1e-06 
3.0 1.171 0 3.0 1e-06 
0.05 1.172 0 3.0 1e-06 
3.0 1.172 0 3.0 1e-06 
0.05 1.173 0 3.0 1e-06 
3.0 1.173 0 3.0 1e-06 
0.05 1.174 0 3.0 1e-06 
3.0 1.174 0 3.0 1e-06 
0.05 1.175 0 3.0 1e-06 
3.0 1.175 0 3.0 1e-06 
0.05 1.176 0 3.0 1e-06 
3.0 1.176 0 3.0 1e-06 
0.05 1.177 0 3.0 1e-06 
3.0 1.177 0 3.0 1e-06 
0.05 1.178 0 3.0 1e-06 
3.0 1.178 0 3.0 1e-06 
0.05 1.179 0 3.0 1e-06 
3.0 1.179 0 3.0 1e-06 
0.05 1.18 0 3.0 1e-06 
3.0 1.18 0 3.0 1e-06 
0.05 1.181 0 3.0 1e-06 
3.0 1.181 0 3.0 1e-06 
0.05 1.182 0 3.0 1e-06 
3.0 1.182 0 3.0 1e-06 
0.05 1.183 0 3.0 1e-06 
3.0 1.183 0 3.0 1e-06 
0.05 1.184 0 3.0 1e-06 
3.0 1.184 0 3.0 1e-06 
0.05 1.185 0 3.0 1e-06 
3.0 1.185 0 3.0 1e-06 
0.05 1.186 0 3.0 1e-06 
3.0 1.186 0 3.0 1e-06 
0.05 1.187 0 3.0 1e-06 
3.0 1.187 0 3.0 1e-06 
0.05 1.188 0 3.0 1e-06 
3.0 1.188 0 3.0 1e-06 
0.05 1.189 0 3.0 1e-06 
3.0 1.189 0 3.0 1e-06 
0.05 1.19 0 3.0 1e-06 
3.0 1.19 0 3.0 1e-06 
0.05 1.191 0 3.0 1e-06 
3.0 1.191 0 3.0 1e-06 
0.05 1.192 0 3.0 1e-06 
3.0 1.192 0 3.0 1e-06 
0.05 1.193 0 3.0 1e-06 
3.0 1.193 0 3.0 1e-06 
0.05 1.194 0 3.0 1e-06 
3.0 1.194 0 3.0 1e-06 
0.05 1.195 0 3.0 1e-06 
3.0 1.195 0 3.0 1e-06 
0.05 1.196 0 3.0 1e-06 
3.0 1.196 0 3.0 1e-06 
0.05 1.197 0 3.0 1e-06 
3.0 1.197 0 3.0 1e-06 
0.05 1.198 0 3.0 1e-06 
3.0 1.198 0 3.0 1e-06 
0.05 1.199 0 3.0 1e-06 
3.0 1.199 0 3.0 1e-06 
0.05 1.2 0 3.0 1e-06 
3.0 1.2 0 3.0 1e-06 
0.05 1.201 0 3.0 1e-06 
3.0 1.201 0 3.0 1e-06 
0.05 1.202 0 3.0 1e-06 
3.0 1.202 0 3.0 1e-06 
0.05 1.203 0 3.0 1e-06 
3.0 1.203 0 3.0 1e-06 
0.05 1.204 0 3.0 1e-06 
3.0 1.204 0 3.0 1e-06 
0.05 1.205 0 3.0 1e-06 
3.0 1.205 0 3.0 1e-06 
0.05 1.206 0 3.0 1e-06 
3.0 1.206 0 3.0 1e-06 
0.05 1.207 0 3.0 1e-06 
3.0 1.207 0 3.0 1e-06 
0.05 1.208 0 3.0 1e-06 
3.0 1.208 0 3.0 1e-06 
0.05 1.209 0 3.0 1e-06 
3.0 1.209 0 3.0 1e-06 
0.05 1.21 0 3.0 1e-06 
3.0 1.21 0 3.0 1e-06 
0.05 1.211 0 3.0 1e-06 
3.0 1.211 0 3.0 1e-06 
0.05 1.212 0 3.0 1e-06 
3.0 1.212 0 3.0 1e-06 
0.05 1.213 0 3.0 1e-06 
3.0 1.213 0 3.0 1e-06 
0.05 1.214 0 3.0 1e-06 
3.0 1.214 0 3.0 1e-06 
0.05 1.215 0 3.0 1e-06 
3.0 1.215 0 3.0 1e-06 
0.05 1.216 0 3.0 1e-06 
3.0 1.216 0 3.0 1e-06 
0.05 1.217 0 3.0 1e-06 
3.0 1.217 0 3.0 1e-06 
0.05 1.218 0 3.0 1e-06 
3.0 1.218 0 3.0 1e-06 
0.05 1.219 0 3.0 1e-06 
3.0 1.219 0 3.0 1e-06 
0.05 1.22 0 3.0 1e-06 
3.0 1.22 0 3.0 1e-06 
0.05 1.221 0 3.0 1e-06 
3.0 1.221 0 3.0 1e-06 
0.05 1.222 0 3.0 1e-06 
3.0 1.222 0 3.0 1e-06 
0.05 1.223 0 3.0 1e-06 
3.0 1.223 0 3.0 1e-06 
0.05 1.224 0 3.0 1e-06 
3.0 1.224 0 3.0 1e-06 
0.05 1.225 0 3.0 1e-06 
3.0 1.225 0 3.0 1e-06 
0.05 1.226 0 3.0 1e-06 
3.0 1.226 0 3.0 1e-06 
0.05 1.227 0 3.0 1e-06 
3.0 1.227 0 3.0 1e-06 
0.05 1.228 0 3.0 1e-06 
3.0 1.228 0 3.0 1e-06 
0.05 1.229 0 3.0 1e-06 
3.0 1.229 0 3.0 1e-06 
0.05 1.23 0 3.0 1e-06 
3.0 1.23 0 3.0 1e-06 
0.05 1.231 0 3.0 1e-06 
3.0 1.231 0 3.0 1e-06 
0.05 1.232 0 3.0 1e-06 
3.0 1.232 0 3.0 1e-06 
0.05 1.233 0 3.0 1e-06 
3.0 1.233 0 3.0 1e-06 
0.05 1.234 0 3.0 1e-06 
3.0 1.234 0 3.0 1e-06 
0.05 1.235 0 3.0 1e-06 
3.0 1.235 0 3.0 1e-06 
0.05 1.236 0 3.0 1e-06 
3.0 1.236 0 3.0 1e-06 
0.05 1.237 0 3.0 1e-06 
3.0 1.237 0 3.0 1e-06 
0.05 1.238 0 3.0 1e-06 
3.0 1.238 0 3.0 1e-06 
0.05 1.239 0 3.0 1e-06 
3.0 1.239 0 3.0 1e-06 
0.05 1.24 0 3.0 1e-06 
3.0 1.24 0 3.0 1e-06 
0.05 1.241 0 3.0 1e-06 
3.0 1.241 0 3.0 1e-06 
0.05 1.242 0 3.0 1e-06 
3.0 1.242 0 3.0 1e-06 
0.05 1.243 0 3.0 1e-06 
3.0 1.243 0 3.0 1e-06 
0.05 1.244 0 3.0 1e-06 
3.0 1.244 0 3.0 1e-06 
0.05 1.245 0 3.0 1e-06 
3.0 1.245 0 3.0 1e-06 
0.05 1.246 0 3.0 1e-06 
3.0 1.246 0 3.0 1e-06 
0.05 1.247 0 3.0 1e-06 
3.0 1.247 0 3.0 1e-06 
0.05 1.248 0 3.0 1e-06 
3.0 1.248 0 3.0 1e-06 
0.05 1.249 0 3.0 1e-06 
3.0 1.249 0 3.0 1e-06 
0.05 1.25 0 3.0 1e-06 
3.0 1.25 0 3.0 1e-06 
0.05 1.251 0 3.0 1e-06 
3.0 1.251 0 3.0 1e-06 
0.05 1.252 0 3.0 1e-06 
3.0 1.252 0 3.0 1e-06 
0.05 1.253 0 3.0 1e-06 
3.0 1.253 0 3.0 1e-06 
0.05 1.254 0 3.0 1e-06 
3.0 1.254 0 3.0 1e-06 
0.05 1.255 0 3.0 1e-06 
3.0 1.255 0 3.0 1e-06 
0.05 1.256 0 3.0 1e-06 
3.0 1.256 0 3.0 1e-06 
0.05 1.257 0 3.0 1e-06 
3.0 1.257 0 3.0 1e-06 
0.05 1.258 0 3.0 1e-06 
3.0 1.258 0 3.0 1e-06 
0.05 1.259 0 3.0 1e-06 
3.0 1.259 0 3.0 1e-06 
0.05 1.26 0 3.0 1e-06 
3.0 1.26 0 3.0 1e-06 
0.05 1.261 0 3.0 1e-06 
3.0 1.261 0 3.0 1e-06 
0.05 1.262 0 3.0 1e-06 
3.0 1.262 0 3.0 1e-06 
0.05 1.263 0 3.0 1e-06 
3.0 1.263 0 3.0 1e-06 
0.05 1.264 0 3.0 1e-06 
3.0 1.264 0 3.0 1e-06 
0.05 1.265 0 3.0 1e-06 
3.0 1.265 0 3.0 1e-06 
0.05 1.266 0 3.0 1e-06 
3.0 1.266 0 3.0 1e-06 
0.05 1.267 0 3.0 1e-06 
3.0 1.267 0 3.0 1e-06 
0.05 1.268 0 3.0 1e-06 
3.0 1.268 0 3.0 1e-06 
0.05 1.269 0 3.0 1e-06 
3.0 1.269 0 3.0 1e-06 
0.05 1.27 0 3.0 1e-06 
3.0 1.27 0 3.0 1e-06 
0.05 1.271 0 3.0 1e-06 
3.0 1.271 0 3.0 1e-06 
0.05 1.272 0 3.0 1e-06 
3.0 1.272 0 3.0 1e-06 
0.05 1.273 0 3.0 1e-06 
3.0 1.273 0 3.0 1e-06 
0.05 1.274 0 3.0 1e-06 
3.0 1.274 0 3.0 1e-06 
0.05 1.275 0 3.0 1e-06 
3.0 1.275 0 3.0 1e-06 
0.05 1.276 0 3.0 1e-06 
3.0 1.276 0 3.0 1e-06 
0.05 1.277 0 3.0 1e-06 
3.0 1.277 0 3.0 1e-06 
0.05 1.278 0 3.0 1e-06 
3.0 1.278 0 3.0 1e-06 
0.05 1.279 0 3.0 1e-06 
3.0 1.279 0 3.0 1e-06 
0.05 1.28 0 3.0 1e-06 
3.0 1.28 0 3.0 1e-06 
0.05 1.281 0 3.0 1e-06 
3.0 1.281 0 3.0 1e-06 
0.05 1.282 0 3.0 1e-06 
3.0 1.282 0 3.0 1e-06 
0.05 1.283 0 3.0 1e-06 
3.0 1.283 0 3.0 1e-06 
0.05 1.284 0 3.0 1e-06 
3.0 1.284 0 3.0 1e-06 
0.05 1.285 0 3.0 1e-06 
3.0 1.285 0 3.0 1e-06 
0.05 1.286 0 3.0 1e-06 
3.0 1.286 0 3.0 1e-06 
0.05 1.287 0 3.0 1e-06 
3.0 1.287 0 3.0 1e-06 
0.05 1.288 0 3.0 1e-06 
3.0 1.288 0 3.0 1e-06 
0.05 1.289 0 3.0 1e-06 
3.0 1.289 0 3.0 1e-06 
0.05 1.29 0 3.0 1e-06 
3.0 1.29 0 3.0 1e-06 
0.05 1.291 0 3.0 1e-06 
3.0 1.291 0 3.0 1e-06 
0.05 1.292 0 3.0 1e-06 
3.0 1.292 0 3.0 1e-06 
0.05 1.293 0 3.0 1e-06 
3.0 1.293 0 3.0 1e-06 
0.05 1.294 0 3.0 1e-06 
3.0 1.294 0 3.0 1e-06 
0.05 1.295 0 3.0 1e-06 
3.0 1.295 0 3.0 1e-06 
0.05 1.296 0 3.0 1e-06 
3.0 1.296 0 3.0 1e-06 
0.05 1.297 0 3.0 1e-06 
3.0 1.297 0 3.0 1e-06 
0.05 1.298 0 3.0 1e-06 
3.0 1.298 0 3.0 1e-06 
0.05 1.299 0 3.0 1e-06 
3.0 1.299 0 3.0 1e-06 
0.05 1.3 0 3.0 1e-06 
3.0 1.3 0 3.0 1e-06 
0.05 1.301 0 3.0 1e-06 
3.0 1.301 0 3.0 1e-06 
0.05 1.302 0 3.0 1e-06 
3.0 1.302 0 3.0 1e-06 
0.05 1.303 0 3.0 1e-06 
3.0 1.303 0 3.0 1e-06 
0.05 1.304 0 3.0 1e-06 
3.0 1.304 0 3.0 1e-06 
0.05 1.305 0 3.0 1e-06 
3.0 1.305 0 3.0 1e-06 
0.05 1.306 0 3.0 1e-06 
3.0 1.306 0 3.0 1e-06 
0.05 1.307 0 3.0 1e-06 
3.0 1.307 0 3.0 1e-06 
0.05 1.308 0 3.0 1e-06 
3.0 1.308 0 3.0 1e-06 
0.05 1.309 0 3.0 1e-06 
3.0 1.309 0 3.0 1e-06 
0.05 1.31 0 3.0 1e-06 
3.0 1.31 0 3.0 1e-06 
0.05 1.311 0 3.0 1e-06 
3.0 1.311 0 3.0 1e-06 
0.05 1.312 0 3.0 1e-06 
3.0 1.312 0 3.0 1e-06 
0.05 1.313 0 3.0 1e-06 
3.0 1.313 0 3.0 1e-06 
0.05 1.314 0 3.0 1e-06 
3.0 1.314 0 3.0 1e-06 
0.05 1.315 0 3.0 1e-06 
3.0 1.315 0 3.0 1e-06 
0.05 1.316 0 3.0 1e-06 
3.0 1.316 0 3.0 1e-06 
0.05 1.317 0 3.0 1e-06 
3.0 1.317 0 3.0 1e-06 
0.05 1.318 0 3.0 1e-06 
3.0 1.318 0 3.0 1e-06 
0.05 1.319 0 3.0 1e-06 
3.0 1.319 0 3.0 1e-06 
0.05 1.32 0 3.0 1e-06 
3.0 1.32 0 3.0 1e-06 
0.05 1.321 0 3.0 1e-06 
3.0 1.321 0 3.0 1e-06 
0.05 1.322 0 3.0 1e-06 
3.0 1.322 0 3.0 1e-06 
0.05 1.323 0 3.0 1e-06 
3.0 1.323 0 3.0 1e-06 
0.05 1.324 0 3.0 1e-06 
3.0 1.324 0 3.0 1e-06 
0.05 1.325 0 3.0 1e-06 
3.0 1.325 0 3.0 1e-06 
0.05 1.326 0 3.0 1e-06 
3.0 1.326 0 3.0 1e-06 
0.05 1.327 0 3.0 1e-06 
3.0 1.327 0 3.0 1e-06 
0.05 1.328 0 3.0 1e-06 
3.0 1.328 0 3.0 1e-06 
0.05 1.329 0 3.0 1e-06 
3.0 1.329 0 3.0 1e-06 
0.05 1.33 0 3.0 1e-06 
3.0 1.33 0 3.0 1e-06 
0.05 1.331 0 3.0 1e-06 
3.0 1.331 0 3.0 1e-06 
0.05 1.332 0 3.0 1e-06 
3.0 1.332 0 3.0 1e-06 
0.05 1.333 0 3.0 1e-06 
3.0 1.333 0 3.0 1e-06 
0.05 1.334 0 3.0 1e-06 
3.0 1.334 0 3.0 1e-06 
0.05 1.335 0 3.0 1e-06 
3.0 1.335 0 3.0 1e-06 
0.05 1.336 0 3.0 1e-06 
3.0 1.336 0 3.0 1e-06 
0.05 1.337 0 3.0 1e-06 
3.0 1.337 0 3.0 1e-06 
0.05 1.338 0 3.0 1e-06 
3.0 1.338 0 3.0 1e-06 
0.05 1.339 0 3.0 1e-06 
3.0 1.339 0 3.0 1e-06 
0.05 1.34 0 3.0 1e-06 
3.0 1.34 0 3.0 1e-06 
0.05 1.341 0 3.0 1e-06 
3.0 1.341 0 3.0 1e-06 
0.05 1.342 0 3.0 1e-06 
3.0 1.342 0 3.0 1e-06 
0.05 1.343 0 3.0 1e-06 
3.0 1.343 0 3.0 1e-06 
0.05 1.344 0 3.0 1e-06 
3.0 1.344 0 3.0 1e-06 
0.05 1.345 0 3.0 1e-06 
3.0 1.345 0 3.0 1e-06 
0.05 1.346 0 3.0 1e-06 
3.0 1.346 0 3.0 1e-06 
0.05 1.347 0 3.0 1e-06 
3.0 1.347 0 3.0 1e-06 
0.05 1.348 0 3.0 1e-06 
3.0 1.348 0 3.0 1e-06 
0.05 1.349 0 3.0 1e-06 
3.0 1.349 0 3.0 1e-06 
0.05 1.35 0 3.0 1e-06 
3.0 1.35 0 3.0 1e-06 
0.05 1.351 0 3.0 1e-06 
3.0 1.351 0 3.0 1e-06 
0.05 1.352 0 3.0 1e-06 
3.0 1.352 0 3.0 1e-06 
0.05 1.353 0 3.0 1e-06 
3.0 1.353 0 3.0 1e-06 
0.05 1.354 0 3.0 1e-06 
3.0 1.354 0 3.0 1e-06 
0.05 1.355 0 3.0 1e-06 
3.0 1.355 0 3.0 1e-06 
0.05 1.356 0 3.0 1e-06 
3.0 1.356 0 3.0 1e-06 
0.05 1.357 0 3.0 1e-06 
3.0 1.357 0 3.0 1e-06 
0.05 1.358 0 3.0 1e-06 
3.0 1.358 0 3.0 1e-06 
0.05 1.359 0 3.0 1e-06 
3.0 1.359 0 3.0 1e-06 
0.05 1.36 0 3.0 1e-06 
3.0 1.36 0 3.0 1e-06 
0.05 1.361 0 3.0 1e-06 
3.0 1.361 0 3.0 1e-06 
0.05 1.362 0 3.0 1e-06 
3.0 1.362 0 3.0 1e-06 
0.05 1.363 0 3.0 1e-06 
3.0 1.363 0 3.0 1e-06 
0.05 1.364 0 3.0 1e-06 
3.0 1.364 0 3.0 1e-06 
0.05 1.365 0 3.0 1e-06 
3.0 1.365 0 3.0 1e-06 
0.05 1.366 0 3.0 1e-06 
3.0 1.366 0 3.0 1e-06 
0.05 1.367 0 3.0 1e-06 
3.0 1.367 0 3.0 1e-06 
0.05 1.368 0 3.0 1e-06 
3.0 1.368 0 3.0 1e-06 
0.05 1.369 0 3.0 1e-06 
3.0 1.369 0 3.0 1e-06 
0.05 1.37 0 3.0 1e-06 
3.0 1.37 0 3.0 1e-06 
0.05 1.371 0 3.0 1e-06 
3.0 1.371 0 3.0 1e-06 
0.05 1.372 0 3.0 1e-06 
3.0 1.372 0 3.0 1e-06 
0.05 1.373 0 3.0 1e-06 
3.0 1.373 0 3.0 1e-06 
0.05 1.374 0 3.0 1e-06 
3.0 1.374 0 3.0 1e-06 
0.05 1.375 0 3.0 1e-06 
3.0 1.375 0 3.0 1e-06 
0.05 1.376 0 3.0 1e-06 
3.0 1.376 0 3.0 1e-06 
0.05 1.377 0 3.0 1e-06 
3.0 1.377 0 3.0 1e-06 
0.05 1.378 0 3.0 1e-06 
3.0 1.378 0 3.0 1e-06 
0.05 1.379 0 3.0 1e-06 
3.0 1.379 0 3.0 1e-06 
0.05 1.38 0 3.0 1e-06 
3.0 1.38 0 3.0 1e-06 
0.05 1.381 0 3.0 1e-06 
3.0 1.381 0 3.0 1e-06 
0.05 1.382 0 3.0 1e-06 
3.0 1.382 0 3.0 1e-06 
0.05 1.383 0 3.0 1e-06 
3.0 1.383 0 3.0 1e-06 
0.05 1.384 0 3.0 1e-06 
3.0 1.384 0 3.0 1e-06 
0.05 1.385 0 3.0 1e-06 
3.0 1.385 0 3.0 1e-06 
0.05 1.386 0 3.0 1e-06 
3.0 1.386 0 3.0 1e-06 
0.05 1.387 0 3.0 1e-06 
3.0 1.387 0 3.0 1e-06 
0.05 1.388 0 3.0 1e-06 
3.0 1.388 0 3.0 1e-06 
0.05 1.389 0 3.0 1e-06 
3.0 1.389 0 3.0 1e-06 
0.05 1.39 0 3.0 1e-06 
3.0 1.39 0 3.0 1e-06 
0.05 1.391 0 3.0 1e-06 
3.0 1.391 0 3.0 1e-06 
0.05 1.392 0 3.0 1e-06 
3.0 1.392 0 3.0 1e-06 
0.05 1.393 0 3.0 1e-06 
3.0 1.393 0 3.0 1e-06 
0.05 1.394 0 3.0 1e-06 
3.0 1.394 0 3.0 1e-06 
0.05 1.395 0 3.0 1e-06 
3.0 1.395 0 3.0 1e-06 
0.05 1.396 0 3.0 1e-06 
3.0 1.396 0 3.0 1e-06 
0.05 1.397 0 3.0 1e-06 
3.0 1.397 0 3.0 1e-06 
0.05 1.398 0 3.0 1e-06 
3.0 1.398 0 3.0 1e-06 
0.05 1.399 0 3.0 1e-06 
3.0 1.399 0 3.0 1e-06 
0.05 1.4 0 3.0 1e-06 
3.0 1.4 0 3.0 1e-06 
0.05 1.401 0 3.0 1e-06 
3.0 1.401 0 3.0 1e-06 
0.05 1.402 0 3.0 1e-06 
3.0 1.402 0 3.0 1e-06 
0.05 1.403 0 3.0 1e-06 
3.0 1.403 0 3.0 1e-06 
0.05 1.404 0 3.0 1e-06 
3.0 1.404 0 3.0 1e-06 
0.05 1.405 0 3.0 1e-06 
3.0 1.405 0 3.0 1e-06 
0.05 1.406 0 3.0 1e-06 
3.0 1.406 0 3.0 1e-06 
0.05 1.407 0 3.0 1e-06 
3.0 1.407 0 3.0 1e-06 
0.05 1.408 0 3.0 1e-06 
3.0 1.408 0 3.0 1e-06 
0.05 1.409 0 3.0 1e-06 
3.0 1.409 0 3.0 1e-06 
0.05 1.41 0 3.0 1e-06 
3.0 1.41 0 3.0 1e-06 
0.05 1.411 0 3.0 1e-06 
3.0 1.411 0 3.0 1e-06 
0.05 1.412 0 3.0 1e-06 
3.0 1.412 0 3.0 1e-06 
0.05 1.413 0 3.0 1e-06 
3.0 1.413 0 3.0 1e-06 
0.05 1.414 0 3.0 1e-06 
3.0 1.414 0 3.0 1e-06 
0.05 1.415 0 3.0 1e-06 
3.0 1.415 0 3.0 1e-06 
0.05 1.416 0 3.0 1e-06 
3.0 1.416 0 3.0 1e-06 
0.05 1.417 0 3.0 1e-06 
3.0 1.417 0 3.0 1e-06 
0.05 1.418 0 3.0 1e-06 
3.0 1.418 0 3.0 1e-06 
0.05 1.419 0 3.0 1e-06 
3.0 1.419 0 3.0 1e-06 
0.05 1.42 0 3.0 1e-06 
3.0 1.42 0 3.0 1e-06 
0.05 1.421 0 3.0 1e-06 
3.0 1.421 0 3.0 1e-06 
0.05 1.422 0 3.0 1e-06 
3.0 1.422 0 3.0 1e-06 
0.05 1.423 0 3.0 1e-06 
3.0 1.423 0 3.0 1e-06 
0.05 1.424 0 3.0 1e-06 
3.0 1.424 0 3.0 1e-06 
0.05 1.425 0 3.0 1e-06 
3.0 1.425 0 3.0 1e-06 
0.05 1.426 0 3.0 1e-06 
3.0 1.426 0 3.0 1e-06 
0.05 1.427 0 3.0 1e-06 
3.0 1.427 0 3.0 1e-06 
0.05 1.428 0 3.0 1e-06 
3.0 1.428 0 3.0 1e-06 
0.05 1.429 0 3.0 1e-06 
3.0 1.429 0 3.0 1e-06 
0.05 1.43 0 3.0 1e-06 
3.0 1.43 0 3.0 1e-06 
0.05 1.431 0 3.0 1e-06 
3.0 1.431 0 3.0 1e-06 
0.05 1.432 0 3.0 1e-06 
3.0 1.432 0 3.0 1e-06 
0.05 1.433 0 3.0 1e-06 
3.0 1.433 0 3.0 1e-06 
0.05 1.434 0 3.0 1e-06 
3.0 1.434 0 3.0 1e-06 
0.05 1.435 0 3.0 1e-06 
3.0 1.435 0 3.0 1e-06 
0.05 1.436 0 3.0 1e-06 
3.0 1.436 0 3.0 1e-06 
0.05 1.437 0 3.0 1e-06 
3.0 1.437 0 3.0 1e-06 
0.05 1.438 0 3.0 1e-06 
3.0 1.438 0 3.0 1e-06 
0.05 1.439 0 3.0 1e-06 
3.0 1.439 0 3.0 1e-06 
0.05 1.44 0 3.0 1e-06 
3.0 1.44 0 3.0 1e-06 
0.05 1.441 0 3.0 1e-06 
3.0 1.441 0 3.0 1e-06 
0.05 1.442 0 3.0 1e-06 
3.0 1.442 0 3.0 1e-06 
0.05 1.443 0 3.0 1e-06 
3.0 1.443 0 3.0 1e-06 
0.05 1.444 0 3.0 1e-06 
3.0 1.444 0 3.0 1e-06 
0.05 1.445 0 3.0 1e-06 
3.0 1.445 0 3.0 1e-06 
0.05 1.446 0 3.0 1e-06 
3.0 1.446 0 3.0 1e-06 
0.05 1.447 0 3.0 1e-06 
3.0 1.447 0 3.0 1e-06 
0.05 1.448 0 3.0 1e-06 
3.0 1.448 0 3.0 1e-06 
0.05 1.449 0 3.0 1e-06 
3.0 1.449 0 3.0 1e-06 
0.05 1.45 0 3.0 1e-06 
3.0 1.45 0 3.0 1e-06 
0.05 1.451 0 3.0 1e-06 
3.0 1.451 0 3.0 1e-06 
0.05 1.452 0 3.0 1e-06 
3.0 1.452 0 3.0 1e-06 
0.05 1.453 0 3.0 1e-06 
3.0 1.453 0 3.0 1e-06 
0.05 1.454 0 3.0 1e-06 
3.0 1.454 0 3.0 1e-06 
0.05 1.455 0 3.0 1e-06 
3.0 1.455 0 3.0 1e-06 
0.05 1.456 0 3.0 1e-06 
3.0 1.456 0 3.0 1e-06 
0.05 1.457 0 3.0 1e-06 
3.0 1.457 0 3.0 1e-06 
0.05 1.458 0 3.0 1e-06 
3.0 1.458 0 3.0 1e-06 
0.05 1.459 0 3.0 1e-06 
3.0 1.459 0 3.0 1e-06 
0.05 1.46 0 3.0 1e-06 
3.0 1.46 0 3.0 1e-06 
0.05 1.461 0 3.0 1e-06 
3.0 1.461 0 3.0 1e-06 
0.05 1.462 0 3.0 1e-06 
3.0 1.462 0 3.0 1e-06 
0.05 1.463 0 3.0 1e-06 
3.0 1.463 0 3.0 1e-06 
0.05 1.464 0 3.0 1e-06 
3.0 1.464 0 3.0 1e-06 
0.05 1.465 0 3.0 1e-06 
3.0 1.465 0 3.0 1e-06 
0.05 1.466 0 3.0 1e-06 
3.0 1.466 0 3.0 1e-06 
0.05 1.467 0 3.0 1e-06 
3.0 1.467 0 3.0 1e-06 
0.05 1.468 0 3.0 1e-06 
3.0 1.468 0 3.0 1e-06 
0.05 1.469 0 3.0 1e-06 
3.0 1.469 0 3.0 1e-06 
0.05 1.47 0 3.0 1e-06 
3.0 1.47 0 3.0 1e-06 
0.05 1.471 0 3.0 1e-06 
3.0 1.471 0 3.0 1e-06 
0.05 1.472 0 3.0 1e-06 
3.0 1.472 0 3.0 1e-06 
0.05 1.473 0 3.0 1e-06 
3.0 1.473 0 3.0 1e-06 
0.05 1.474 0 3.0 1e-06 
3.0 1.474 0 3.0 1e-06 
0.05 1.475 0 3.0 1e-06 
3.0 1.475 0 3.0 1e-06 
0.05 1.476 0 3.0 1e-06 
3.0 1.476 0 3.0 1e-06 
0.05 1.477 0 3.0 1e-06 
3.0 1.477 0 3.0 1e-06 
0.05 1.478 0 3.0 1e-06 
3.0 1.478 0 3.0 1e-06 
0.05 1.479 0 3.0 1e-06 
3.0 1.479 0 3.0 1e-06 
0.05 1.48 0 3.0 1e-06 
3.0 1.48 0 3.0 1e-06 
0.05 1.481 0 3.0 1e-06 
3.0 1.481 0 3.0 1e-06 
0.05 1.482 0 3.0 1e-06 
3.0 1.482 0 3.0 1e-06 
0.05 1.483 0 3.0 1e-06 
3.0 1.483 0 3.0 1e-06 
0.05 1.484 0 3.0 1e-06 
3.0 1.484 0 3.0 1e-06 
0.05 1.485 0 3.0 1e-06 
3.0 1.485 0 3.0 1e-06 
0.05 1.486 0 3.0 1e-06 
3.0 1.486 0 3.0 1e-06 
0.05 1.487 0 3.0 1e-06 
3.0 1.487 0 3.0 1e-06 
0.05 1.488 0 3.0 1e-06 
3.0 1.488 0 3.0 1e-06 
0.05 1.489 0 3.0 1e-06 
3.0 1.489 0 3.0 1e-06 
0.05 1.49 0 3.0 1e-06 
3.0 1.49 0 3.0 1e-06 
0.05 1.491 0 3.0 1e-06 
3.0 1.491 0 3.0 1e-06 
0.05 1.492 0 3.0 1e-06 
3.0 1.492 0 3.0 1e-06 
0.05 1.493 0 3.0 1e-06 
3.0 1.493 0 3.0 1e-06 
0.05 1.494 0 3.0 1e-06 
3.0 1.494 0 3.0 1e-06 
0.05 1.495 0 3.0 1e-06 
3.0 1.495 0 3.0 1e-06 
0.05 1.496 0 3.0 1e-06 
3.0 1.496 0 3.0 1e-06 
0.05 1.497 0 3.0 1e-06 
3.0 1.497 0 3.0 1e-06 
0.05 1.498 0 3.0 1e-06 
3.0 1.498 0 3.0 1e-06 
0.05 1.499 0 3.0 1e-06 
3.0 1.499 0 3.0 1e-06 
0.05 1.5 0 3.0 1e-06 
3.0 1.5 0 3.0 1e-06 
0.05 1.501 0 3.0 1e-06 
3.0 1.501 0 3.0 1e-06 
0.05 1.502 0 3.0 1e-06 
3.0 1.502 0 3.0 1e-06 
0.05 1.503 0 3.0 1e-06 
3.0 1.503 0 3.0 1e-06 
0.05 1.504 0 3.0 1e-06 
3.0 1.504 0 3.0 1e-06 
0.05 1.505 0 3.0 1e-06 
3.0 1.505 0 3.0 1e-06 
0.05 1.506 0 3.0 1e-06 
3.0 1.506 0 3.0 1e-06 
0.05 1.507 0 3.0 1e-06 
3.0 1.507 0 3.0 1e-06 
0.05 1.508 0 3.0 1e-06 
3.0 1.508 0 3.0 1e-06 
0.05 1.509 0 3.0 1e-06 
3.0 1.509 0 3.0 1e-06 
0.05 1.51 0 3.0 1e-06 
3.0 1.51 0 3.0 1e-06 
0.05 1.511 0 3.0 1e-06 
3.0 1.511 0 3.0 1e-06 
0.05 1.512 0 3.0 1e-06 
3.0 1.512 0 3.0 1e-06 
0.05 1.513 0 3.0 1e-06 
3.0 1.513 0 3.0 1e-06 
0.05 1.514 0 3.0 1e-06 
3.0 1.514 0 3.0 1e-06 
0.05 1.515 0 3.0 1e-06 
3.0 1.515 0 3.0 1e-06 
0.05 1.516 0 3.0 1e-06 
3.0 1.516 0 3.0 1e-06 
0.05 1.517 0 3.0 1e-06 
3.0 1.517 0 3.0 1e-06 
0.05 1.518 0 3.0 1e-06 
3.0 1.518 0 3.0 1e-06 
0.05 1.519 0 3.0 1e-06 
3.0 1.519 0 3.0 1e-06 
0.05 1.52 0 3.0 1e-06 
3.0 1.52 0 3.0 1e-06 
0.05 1.521 0 3.0 1e-06 
3.0 1.521 0 3.0 1e-06 
0.05 1.522 0 3.0 1e-06 
3.0 1.522 0 3.0 1e-06 
0.05 1.523 0 3.0 1e-06 
3.0 1.523 0 3.0 1e-06 
0.05 1.524 0 3.0 1e-06 
3.0 1.524 0 3.0 1e-06 
0.05 1.525 0 3.0 1e-06 
3.0 1.525 0 3.0 1e-06 
0.05 1.526 0 3.0 1e-06 
3.0 1.526 0 3.0 1e-06 
0.05 1.527 0 3.0 1e-06 
3.0 1.527 0 3.0 1e-06 
0.05 1.528 0 3.0 1e-06 
3.0 1.528 0 3.0 1e-06 
0.05 1.529 0 3.0 1e-06 
3.0 1.529 0 3.0 1e-06 
0.05 1.53 0 3.0 1e-06 
3.0 1.53 0 3.0 1e-06 
0.05 1.531 0 3.0 1e-06 
3.0 1.531 0 3.0 1e-06 
0.05 1.532 0 3.0 1e-06 
3.0 1.532 0 3.0 1e-06 
0.05 1.533 0 3.0 1e-06 
3.0 1.533 0 3.0 1e-06 
0.05 1.534 0 3.0 1e-06 
3.0 1.534 0 3.0 1e-06 
0.05 1.535 0 3.0 1e-06 
3.0 1.535 0 3.0 1e-06 
0.05 1.536 0 3.0 1e-06 
3.0 1.536 0 3.0 1e-06 
0.05 1.537 0 3.0 1e-06 
3.0 1.537 0 3.0 1e-06 
0.05 1.538 0 3.0 1e-06 
3.0 1.538 0 3.0 1e-06 
0.05 1.539 0 3.0 1e-06 
3.0 1.539 0 3.0 1e-06 
0.05 1.54 0 3.0 1e-06 
3.0 1.54 0 3.0 1e-06 
0.05 1.541 0 3.0 1e-06 
3.0 1.541 0 3.0 1e-06 
0.05 1.542 0 3.0 1e-06 
3.0 1.542 0 3.0 1e-06 
0.05 1.543 0 3.0 1e-06 
3.0 1.543 0 3.0 1e-06 
0.05 1.544 0 3.0 1e-06 
3.0 1.544 0 3.0 1e-06 
0.05 1.545 0 3.0 1e-06 
3.0 1.545 0 3.0 1e-06 
0.05 1.546 0 3.0 1e-06 
3.0 1.546 0 3.0 1e-06 
0.05 1.547 0 3.0 1e-06 
3.0 1.547 0 3.0 1e-06 
0.05 1.548 0 3.0 1e-06 
3.0 1.548 0 3.0 1e-06 
0.05 1.549 0 3.0 1e-06 
3.0 1.549 0 3.0 1e-06 
0.05 1.55 0 3.0 1e-06 
3.0 1.55 0 3.0 1e-06 
0.05 1.551 0 3.0 1e-06 
3.0 1.551 0 3.0 1e-06 
0.05 1.552 0 3.0 1e-06 
3.0 1.552 0 3.0 1e-06 
0.05 1.553 0 3.0 1e-06 
3.0 1.553 0 3.0 1e-06 
0.05 1.554 0 3.0 1e-06 
3.0 1.554 0 3.0 1e-06 
0.05 1.555 0 3.0 1e-06 
3.0 1.555 0 3.0 1e-06 
0.05 1.556 0 3.0 1e-06 
3.0 1.556 0 3.0 1e-06 
0.05 1.557 0 3.0 1e-06 
3.0 1.557 0 3.0 1e-06 
0.05 1.558 0 3.0 1e-06 
3.0 1.558 0 3.0 1e-06 
0.05 1.559 0 3.0 1e-06 
3.0 1.559 0 3.0 1e-06 
0.05 1.56 0 3.0 1e-06 
3.0 1.56 0 3.0 1e-06 
0.05 1.561 0 3.0 1e-06 
3.0 1.561 0 3.0 1e-06 
0.05 1.562 0 3.0 1e-06 
3.0 1.562 0 3.0 1e-06 
0.05 1.563 0 3.0 1e-06 
3.0 1.563 0 3.0 1e-06 
0.05 1.564 0 3.0 1e-06 
3.0 1.564 0 3.0 1e-06 
0.05 1.565 0 3.0 1e-06 
3.0 1.565 0 3.0 1e-06 
0.05 1.566 0 3.0 1e-06 
3.0 1.566 0 3.0 1e-06 
0.05 1.567 0 3.0 1e-06 
3.0 1.567 0 3.0 1e-06 
0.05 1.568 0 3.0 1e-06 
3.0 1.568 0 3.0 1e-06 
0.05 1.569 0 3.0 1e-06 
3.0 1.569 0 3.0 1e-06 
0.05 1.57 0 3.0 1e-06 
3.0 1.57 0 3.0 1e-06 
0.05 1.571 0 3.0 1e-06 
3.0 1.571 0 3.0 1e-06 
0.05 1.572 0 3.0 1e-06 
3.0 1.572 0 3.0 1e-06 
0.05 1.573 0 3.0 1e-06 
3.0 1.573 0 3.0 1e-06 
0.05 1.574 0 3.0 1e-06 
3.0 1.574 0 3.0 1e-06 
0.05 1.575 0 3.0 1e-06 
3.0 1.575 0 3.0 1e-06 
0.05 1.576 0 3.0 1e-06 
3.0 1.576 0 3.0 1e-06 
0.05 1.577 0 3.0 1e-06 
3.0 1.577 0 3.0 1e-06 
0.05 1.578 0 3.0 1e-06 
3.0 1.578 0 3.0 1e-06 
0.05 1.579 0 3.0 1e-06 
3.0 1.579 0 3.0 1e-06 
0.05 1.58 0 3.0 1e-06 
3.0 1.58 0 3.0 1e-06 
0.05 1.581 0 3.0 1e-06 
3.0 1.581 0 3.0 1e-06 
0.05 1.582 0 3.0 1e-06 
3.0 1.582 0 3.0 1e-06 
0.05 1.583 0 3.0 1e-06 
3.0 1.583 0 3.0 1e-06 
0.05 1.584 0 3.0 1e-06 
3.0 1.584 0 3.0 1e-06 
0.05 1.585 0 3.0 1e-06 
3.0 1.585 0 3.0 1e-06 
0.05 1.586 0 3.0 1e-06 
3.0 1.586 0 3.0 1e-06 
0.05 1.587 0 3.0 1e-06 
3.0 1.587 0 3.0 1e-06 
0.05 1.588 0 3.0 1e-06 
3.0 1.588 0 3.0 1e-06 
0.05 1.589 0 3.0 1e-06 
3.0 1.589 0 3.0 1e-06 
0.05 1.59 0 3.0 1e-06 
3.0 1.59 0 3.0 1e-06 
0.05 1.591 0 3.0 1e-06 
3.0 1.591 0 3.0 1e-06 
0.05 1.592 0 3.0 1e-06 
3.0 1.592 0 3.0 1e-06 
0.05 1.593 0 3.0 1e-06 
3.0 1.593 0 3.0 1e-06 
0.05 1.594 0 3.0 1e-06 
3.0 1.594 0 3.0 1e-06 
0.05 1.595 0 3.0 1e-06 
3.0 1.595 0 3.0 1e-06 
0.05 1.596 0 3.0 1e-06 
3.0 1.596 0 3.0 1e-06 
0.05 1.597 0 3.0 1e-06 
3.0 1.597 0 3.0 1e-06 
0.05 1.598 0 3.0 1e-06 
3.0 1.598 0 3.0 1e-06 
0.05 1.599 0 3.0 1e-06 
3.0 1.599 0 3.0 1e-06 
0.05 1.6 0 3.0 1e-06 
3.0 1.6 0 3.0 1e-06 
0.05 1.601 0 3.0 1e-06 
3.0 1.601 0 3.0 1e-06 
0.05 1.602 0 3.0 1e-06 
3.0 1.602 0 3.0 1e-06 
0.05 1.603 0 3.0 1e-06 
3.0 1.603 0 3.0 1e-06 
0.05 1.604 0 3.0 1e-06 
3.0 1.604 0 3.0 1e-06 
0.05 1.605 0 3.0 1e-06 
3.0 1.605 0 3.0 1e-06 
0.05 1.606 0 3.0 1e-06 
3.0 1.606 0 3.0 1e-06 
0.05 1.607 0 3.0 1e-06 
3.0 1.607 0 3.0 1e-06 
0.05 1.608 0 3.0 1e-06 
3.0 1.608 0 3.0 1e-06 
0.05 1.609 0 3.0 1e-06 
3.0 1.609 0 3.0 1e-06 
0.05 1.61 0 3.0 1e-06 
3.0 1.61 0 3.0 1e-06 
0.05 1.611 0 3.0 1e-06 
3.0 1.611 0 3.0 1e-06 
0.05 1.612 0 3.0 1e-06 
3.0 1.612 0 3.0 1e-06 
0.05 1.613 0 3.0 1e-06 
3.0 1.613 0 3.0 1e-06 
0.05 1.614 0 3.0 1e-06 
3.0 1.614 0 3.0 1e-06 
0.05 1.615 0 3.0 1e-06 
3.0 1.615 0 3.0 1e-06 
0.05 1.616 0 3.0 1e-06 
3.0 1.616 0 3.0 1e-06 
0.05 1.617 0 3.0 1e-06 
3.0 1.617 0 3.0 1e-06 
0.05 1.618 0 3.0 1e-06 
3.0 1.618 0 3.0 1e-06 
0.05 1.619 0 3.0 1e-06 
3.0 1.619 0 3.0 1e-06 
0.05 1.62 0 3.0 1e-06 
3.0 1.62 0 3.0 1e-06 
0.05 1.621 0 3.0 1e-06 
3.0 1.621 0 3.0 1e-06 
0.05 1.622 0 3.0 1e-06 
3.0 1.622 0 3.0 1e-06 
0.05 1.623 0 3.0 1e-06 
3.0 1.623 0 3.0 1e-06 
0.05 1.624 0 3.0 1e-06 
3.0 1.624 0 3.0 1e-06 
0.05 1.625 0 3.0 1e-06 
3.0 1.625 0 3.0 1e-06 
0.05 1.626 0 3.0 1e-06 
3.0 1.626 0 3.0 1e-06 
0.05 1.627 0 3.0 1e-06 
3.0 1.627 0 3.0 1e-06 
0.05 1.628 0 3.0 1e-06 
3.0 1.628 0 3.0 1e-06 
0.05 1.629 0 3.0 1e-06 
3.0 1.629 0 3.0 1e-06 
0.05 1.63 0 3.0 1e-06 
3.0 1.63 0 3.0 1e-06 
0.05 1.631 0 3.0 1e-06 
3.0 1.631 0 3.0 1e-06 
0.05 1.632 0 3.0 1e-06 
3.0 1.632 0 3.0 1e-06 
0.05 1.633 0 3.0 1e-06 
3.0 1.633 0 3.0 1e-06 
0.05 1.634 0 3.0 1e-06 
3.0 1.634 0 3.0 1e-06 
0.05 1.635 0 3.0 1e-06 
3.0 1.635 0 3.0 1e-06 
0.05 1.636 0 3.0 1e-06 
3.0 1.636 0 3.0 1e-06 
0.05 1.637 0 3.0 1e-06 
3.0 1.637 0 3.0 1e-06 
0.05 1.638 0 3.0 1e-06 
3.0 1.638 0 3.0 1e-06 
0.05 1.639 0 3.0 1e-06 
3.0 1.639 0 3.0 1e-06 
0.05 1.64 0 3.0 1e-06 
3.0 1.64 0 3.0 1e-06 
0.05 1.641 0 3.0 1e-06 
3.0 1.641 0 3.0 1e-06 
0.05 1.642 0 3.0 1e-06 
3.0 1.642 0 3.0 1e-06 
0.05 1.643 0 3.0 1e-06 
3.0 1.643 0 3.0 1e-06 
0.05 1.644 0 3.0 1e-06 
3.0 1.644 0 3.0 1e-06 
0.05 1.645 0 3.0 1e-06 
3.0 1.645 0 3.0 1e-06 
0.05 1.646 0 3.0 1e-06 
3.0 1.646 0 3.0 1e-06 
0.05 1.647 0 3.0 1e-06 
3.0 1.647 0 3.0 1e-06 
0.05 1.648 0 3.0 1e-06 
3.0 1.648 0 3.0 1e-06 
0.05 1.649 0 3.0 1e-06 
3.0 1.649 0 3.0 1e-06 
0.05 1.65 0 3.0 1e-06 
3.0 1.65 0 3.0 1e-06 
0.05 1.651 0 3.0 1e-06 
3.0 1.651 0 3.0 1e-06 
0.05 1.652 0 3.0 1e-06 
3.0 1.652 0 3.0 1e-06 
0.05 1.653 0 3.0 1e-06 
3.0 1.653 0 3.0 1e-06 
0.05 1.654 0 3.0 1e-06 
3.0 1.654 0 3.0 1e-06 
0.05 1.655 0 3.0 1e-06 
3.0 1.655 0 3.0 1e-06 
0.05 1.656 0 3.0 1e-06 
3.0 1.656 0 3.0 1e-06 
0.05 1.657 0 3.0 1e-06 
3.0 1.657 0 3.0 1e-06 
0.05 1.658 0 3.0 1e-06 
3.0 1.658 0 3.0 1e-06 
0.05 1.659 0 3.0 1e-06 
3.0 1.659 0 3.0 1e-06 
0.05 1.66 0 3.0 1e-06 
3.0 1.66 0 3.0 1e-06 
0.05 1.661 0 3.0 1e-06 
3.0 1.661 0 3.0 1e-06 
0.05 1.662 0 3.0 1e-06 
3.0 1.662 0 3.0 1e-06 
0.05 1.663 0 3.0 1e-06 
3.0 1.663 0 3.0 1e-06 
0.05 1.664 0 3.0 1e-06 
3.0 1.664 0 3.0 1e-06 
0.05 1.665 0 3.0 1e-06 
3.0 1.665 0 3.0 1e-06 
0.05 1.666 0 3.0 1e-06 
3.0 1.666 0 3.0 1e-06 
0.05 1.667 0 3.0 1e-06 
3.0 1.667 0 3.0 1e-06 
0.05 1.668 0 3.0 1e-06 
3.0 1.668 0 3.0 1e-06 
0.05 1.669 0 3.0 1e-06 
3.0 1.669 0 3.0 1e-06 
0.05 1.67 0 3.0 1e-06 
3.0 1.67 0 3.0 1e-06 
0.05 1.671 0 3.0 1e-06 
3.0 1.671 0 3.0 1e-06 
0.05 1.672 0 3.0 1e-06 
3.0 1.672 0 3.0 1e-06 
0.05 1.673 0 3.0 1e-06 
3.0 1.673 0 3.0 1e-06 
0.05 1.674 0 3.0 1e-06 
3.0 1.674 0 3.0 1e-06 
0.05 1.675 0 3.0 1e-06 
3.0 1.675 0 3.0 1e-06 
0.05 1.676 0 3.0 1e-06 
3.0 1.676 0 3.0 1e-06 
0.05 1.677 0 3.0 1e-06 
3.0 1.677 0 3.0 1e-06 
0.05 1.678 0 3.0 1e-06 
3.0 1.678 0 3.0 1e-06 
0.05 1.679 0 3.0 1e-06 
3.0 1.679 0 3.0 1e-06 
0.05 1.68 0 3.0 1e-06 
3.0 1.68 0 3.0 1e-06 
0.05 1.681 0 3.0 1e-06 
3.0 1.681 0 3.0 1e-06 
0.05 1.682 0 3.0 1e-06 
3.0 1.682 0 3.0 1e-06 
0.05 1.683 0 3.0 1e-06 
3.0 1.683 0 3.0 1e-06 
0.05 1.684 0 3.0 1e-06 
3.0 1.684 0 3.0 1e-06 
0.05 1.685 0 3.0 1e-06 
3.0 1.685 0 3.0 1e-06 
0.05 1.686 0 3.0 1e-06 
3.0 1.686 0 3.0 1e-06 
0.05 1.687 0 3.0 1e-06 
3.0 1.687 0 3.0 1e-06 
0.05 1.688 0 3.0 1e-06 
3.0 1.688 0 3.0 1e-06 
0.05 1.689 0 3.0 1e-06 
3.0 1.689 0 3.0 1e-06 
0.05 1.69 0 3.0 1e-06 
3.0 1.69 0 3.0 1e-06 
0.05 1.691 0 3.0 1e-06 
3.0 1.691 0 3.0 1e-06 
0.05 1.692 0 3.0 1e-06 
3.0 1.692 0 3.0 1e-06 
0.05 1.693 0 3.0 1e-06 
3.0 1.693 0 3.0 1e-06 
0.05 1.694 0 3.0 1e-06 
3.0 1.694 0 3.0 1e-06 
0.05 1.695 0 3.0 1e-06 
3.0 1.695 0 3.0 1e-06 
0.05 1.696 0 3.0 1e-06 
3.0 1.696 0 3.0 1e-06 
0.05 1.697 0 3.0 1e-06 
3.0 1.697 0 3.0 1e-06 
0.05 1.698 0 3.0 1e-06 
3.0 1.698 0 3.0 1e-06 
0.05 1.699 0 3.0 1e-06 
3.0 1.699 0 3.0 1e-06 
0.05 1.7 0 3.0 1e-06 
3.0 1.7 0 3.0 1e-06 
0.05 1.701 0 3.0 1e-06 
3.0 1.701 0 3.0 1e-06 
0.05 1.702 0 3.0 1e-06 
3.0 1.702 0 3.0 1e-06 
0.05 1.703 0 3.0 1e-06 
3.0 1.703 0 3.0 1e-06 
0.05 1.704 0 3.0 1e-06 
3.0 1.704 0 3.0 1e-06 
0.05 1.705 0 3.0 1e-06 
3.0 1.705 0 3.0 1e-06 
0.05 1.706 0 3.0 1e-06 
3.0 1.706 0 3.0 1e-06 
0.05 1.707 0 3.0 1e-06 
3.0 1.707 0 3.0 1e-06 
0.05 1.708 0 3.0 1e-06 
3.0 1.708 0 3.0 1e-06 
0.05 1.709 0 3.0 1e-06 
3.0 1.709 0 3.0 1e-06 
0.05 1.71 0 3.0 1e-06 
3.0 1.71 0 3.0 1e-06 
0.05 1.711 0 3.0 1e-06 
3.0 1.711 0 3.0 1e-06 
0.05 1.712 0 3.0 1e-06 
3.0 1.712 0 3.0 1e-06 
0.05 1.713 0 3.0 1e-06 
3.0 1.713 0 3.0 1e-06 
0.05 1.714 0 3.0 1e-06 
3.0 1.714 0 3.0 1e-06 
0.05 1.715 0 3.0 1e-06 
3.0 1.715 0 3.0 1e-06 
0.05 1.716 0 3.0 1e-06 
3.0 1.716 0 3.0 1e-06 
0.05 1.717 0 3.0 1e-06 
3.0 1.717 0 3.0 1e-06 
0.05 1.718 0 3.0 1e-06 
3.0 1.718 0 3.0 1e-06 
0.05 1.719 0 3.0 1e-06 
3.0 1.719 0 3.0 1e-06 
0.05 1.72 0 3.0 1e-06 
3.0 1.72 0 3.0 1e-06 
0.05 1.721 0 3.0 1e-06 
3.0 1.721 0 3.0 1e-06 
0.05 1.722 0 3.0 1e-06 
3.0 1.722 0 3.0 1e-06 
0.05 1.723 0 3.0 1e-06 
3.0 1.723 0 3.0 1e-06 
0.05 1.724 0 3.0 1e-06 
3.0 1.724 0 3.0 1e-06 
0.05 1.725 0 3.0 1e-06 
3.0 1.725 0 3.0 1e-06 
0.05 1.726 0 3.0 1e-06 
3.0 1.726 0 3.0 1e-06 
0.05 1.727 0 3.0 1e-06 
3.0 1.727 0 3.0 1e-06 
0.05 1.728 0 3.0 1e-06 
3.0 1.728 0 3.0 1e-06 
0.05 1.729 0 3.0 1e-06 
3.0 1.729 0 3.0 1e-06 
0.05 1.73 0 3.0 1e-06 
3.0 1.73 0 3.0 1e-06 
0.05 1.731 0 3.0 1e-06 
3.0 1.731 0 3.0 1e-06 
0.05 1.732 0 3.0 1e-06 
3.0 1.732 0 3.0 1e-06 
0.05 1.733 0 3.0 1e-06 
3.0 1.733 0 3.0 1e-06 
0.05 1.734 0 3.0 1e-06 
3.0 1.734 0 3.0 1e-06 
0.05 1.735 0 3.0 1e-06 
3.0 1.735 0 3.0 1e-06 
0.05 1.736 0 3.0 1e-06 
3.0 1.736 0 3.0 1e-06 
0.05 1.737 0 3.0 1e-06 
3.0 1.737 0 3.0 1e-06 
0.05 1.738 0 3.0 1e-06 
3.0 1.738 0 3.0 1e-06 
0.05 1.739 0 3.0 1e-06 
3.0 1.739 0 3.0 1e-06 
0.05 1.74 0 3.0 1e-06 
3.0 1.74 0 3.0 1e-06 
0.05 1.741 0 3.0 1e-06 
3.0 1.741 0 3.0 1e-06 
0.05 1.742 0 3.0 1e-06 
3.0 1.742 0 3.0 1e-06 
0.05 1.743 0 3.0 1e-06 
3.0 1.743 0 3.0 1e-06 
0.05 1.744 0 3.0 1e-06 
3.0 1.744 0 3.0 1e-06 
0.05 1.745 0 3.0 1e-06 
3.0 1.745 0 3.0 1e-06 
0.05 1.746 0 3.0 1e-06 
3.0 1.746 0 3.0 1e-06 
0.05 1.747 0 3.0 1e-06 
3.0 1.747 0 3.0 1e-06 
0.05 1.748 0 3.0 1e-06 
3.0 1.748 0 3.0 1e-06 
0.05 1.749 0 3.0 1e-06 
3.0 1.749 0 3.0 1e-06 
0.05 1.75 0 3.0 1e-06 
3.0 1.75 0 3.0 1e-06 
0.05 1.751 0 3.0 1e-06 
3.0 1.751 0 3.0 1e-06 
0.05 1.752 0 3.0 1e-06 
3.0 1.752 0 3.0 1e-06 
0.05 1.753 0 3.0 1e-06 
3.0 1.753 0 3.0 1e-06 
0.05 1.754 0 3.0 1e-06 
3.0 1.754 0 3.0 1e-06 
0.05 1.755 0 3.0 1e-06 
3.0 1.755 0 3.0 1e-06 
0.05 1.756 0 3.0 1e-06 
3.0 1.756 0 3.0 1e-06 
0.05 1.757 0 3.0 1e-06 
3.0 1.757 0 3.0 1e-06 
0.05 1.758 0 3.0 1e-06 
3.0 1.758 0 3.0 1e-06 
0.05 1.759 0 3.0 1e-06 
3.0 1.759 0 3.0 1e-06 
0.05 1.76 0 3.0 1e-06 
3.0 1.76 0 3.0 1e-06 
0.05 1.761 0 3.0 1e-06 
3.0 1.761 0 3.0 1e-06 
0.05 1.762 0 3.0 1e-06 
3.0 1.762 0 3.0 1e-06 
0.05 1.763 0 3.0 1e-06 
3.0 1.763 0 3.0 1e-06 
0.05 1.764 0 3.0 1e-06 
3.0 1.764 0 3.0 1e-06 
0.05 1.765 0 3.0 1e-06 
3.0 1.765 0 3.0 1e-06 
0.05 1.766 0 3.0 1e-06 
3.0 1.766 0 3.0 1e-06 
0.05 1.767 0 3.0 1e-06 
3.0 1.767 0 3.0 1e-06 
0.05 1.768 0 3.0 1e-06 
3.0 1.768 0 3.0 1e-06 
0.05 1.769 0 3.0 1e-06 
3.0 1.769 0 3.0 1e-06 
0.05 1.77 0 3.0 1e-06 
3.0 1.77 0 3.0 1e-06 
0.05 1.771 0 3.0 1e-06 
3.0 1.771 0 3.0 1e-06 
0.05 1.772 0 3.0 1e-06 
3.0 1.772 0 3.0 1e-06 
0.05 1.773 0 3.0 1e-06 
3.0 1.773 0 3.0 1e-06 
0.05 1.774 0 3.0 1e-06 
3.0 1.774 0 3.0 1e-06 
0.05 1.775 0 3.0 1e-06 
3.0 1.775 0 3.0 1e-06 
0.05 1.776 0 3.0 1e-06 
3.0 1.776 0 3.0 1e-06 
0.05 1.777 0 3.0 1e-06 
3.0 1.777 0 3.0 1e-06 
0.05 1.778 0 3.0 1e-06 
3.0 1.778 0 3.0 1e-06 
0.05 1.779 0 3.0 1e-06 
3.0 1.779 0 3.0 1e-06 
0.05 1.78 0 3.0 1e-06 
3.0 1.78 0 3.0 1e-06 
0.05 1.781 0 3.0 1e-06 
3.0 1.781 0 3.0 1e-06 
0.05 1.782 0 3.0 1e-06 
3.0 1.782 0 3.0 1e-06 
0.05 1.783 0 3.0 1e-06 
3.0 1.783 0 3.0 1e-06 
0.05 1.784 0 3.0 1e-06 
3.0 1.784 0 3.0 1e-06 
0.05 1.785 0 3.0 1e-06 
3.0 1.785 0 3.0 1e-06 
0.05 1.786 0 3.0 1e-06 
3.0 1.786 0 3.0 1e-06 
0.05 1.787 0 3.0 1e-06 
3.0 1.787 0 3.0 1e-06 
0.05 1.788 0 3.0 1e-06 
3.0 1.788 0 3.0 1e-06 
0.05 1.789 0 3.0 1e-06 
3.0 1.789 0 3.0 1e-06 
0.05 1.79 0 3.0 1e-06 
3.0 1.79 0 3.0 1e-06 
0.05 1.791 0 3.0 1e-06 
3.0 1.791 0 3.0 1e-06 
0.05 1.792 0 3.0 1e-06 
3.0 1.792 0 3.0 1e-06 
0.05 1.793 0 3.0 1e-06 
3.0 1.793 0 3.0 1e-06 
0.05 1.794 0 3.0 1e-06 
3.0 1.794 0 3.0 1e-06 
0.05 1.795 0 3.0 1e-06 
3.0 1.795 0 3.0 1e-06 
0.05 1.796 0 3.0 1e-06 
3.0 1.796 0 3.0 1e-06 
0.05 1.797 0 3.0 1e-06 
3.0 1.797 0 3.0 1e-06 
0.05 1.798 0 3.0 1e-06 
3.0 1.798 0 3.0 1e-06 
0.05 1.799 0 3.0 1e-06 
3.0 1.799 0 3.0 1e-06 
0.05 1.8 0 3.0 1e-06 
3.0 1.8 0 3.0 1e-06 
0.05 1.801 0 3.0 1e-06 
3.0 1.801 0 3.0 1e-06 
0.05 1.802 0 3.0 1e-06 
3.0 1.802 0 3.0 1e-06 
0.05 1.803 0 3.0 1e-06 
3.0 1.803 0 3.0 1e-06 
0.05 1.804 0 3.0 1e-06 
3.0 1.804 0 3.0 1e-06 
0.05 1.805 0 3.0 1e-06 
3.0 1.805 0 3.0 1e-06 
0.05 1.806 0 3.0 1e-06 
3.0 1.806 0 3.0 1e-06 
0.05 1.807 0 3.0 1e-06 
3.0 1.807 0 3.0 1e-06 
0.05 1.808 0 3.0 1e-06 
3.0 1.808 0 3.0 1e-06 
0.05 1.809 0 3.0 1e-06 
3.0 1.809 0 3.0 1e-06 
0.05 1.81 0 3.0 1e-06 
3.0 1.81 0 3.0 1e-06 
0.05 1.811 0 3.0 1e-06 
3.0 1.811 0 3.0 1e-06 
0.05 1.812 0 3.0 1e-06 
3.0 1.812 0 3.0 1e-06 
0.05 1.813 0 3.0 1e-06 
3.0 1.813 0 3.0 1e-06 
0.05 1.814 0 3.0 1e-06 
3.0 1.814 0 3.0 1e-06 
0.05 1.815 0 3.0 1e-06 
3.0 1.815 0 3.0 1e-06 
0.05 1.816 0 3.0 1e-06 
3.0 1.816 0 3.0 1e-06 
0.05 1.817 0 3.0 1e-06 
3.0 1.817 0 3.0 1e-06 
0.05 1.818 0 3.0 1e-06 
3.0 1.818 0 3.0 1e-06 
0.05 1.819 0 3.0 1e-06 
3.0 1.819 0 3.0 1e-06 
0.05 1.82 0 3.0 1e-06 
3.0 1.82 0 3.0 1e-06 
0.05 1.821 0 3.0 1e-06 
3.0 1.821 0 3.0 1e-06 
0.05 1.822 0 3.0 1e-06 
3.0 1.822 0 3.0 1e-06 
0.05 1.823 0 3.0 1e-06 
3.0 1.823 0 3.0 1e-06 
0.05 1.824 0 3.0 1e-06 
3.0 1.824 0 3.0 1e-06 
0.05 1.825 0 3.0 1e-06 
3.0 1.825 0 3.0 1e-06 
0.05 1.826 0 3.0 1e-06 
3.0 1.826 0 3.0 1e-06 
0.05 1.827 0 3.0 1e-06 
3.0 1.827 0 3.0 1e-06 
0.05 1.828 0 3.0 1e-06 
3.0 1.828 0 3.0 1e-06 
0.05 1.829 0 3.0 1e-06 
3.0 1.829 0 3.0 1e-06 
0.05 1.83 0 3.0 1e-06 
3.0 1.83 0 3.0 1e-06 
0.05 1.831 0 3.0 1e-06 
3.0 1.831 0 3.0 1e-06 
0.05 1.832 0 3.0 1e-06 
3.0 1.832 0 3.0 1e-06 
0.05 1.833 0 3.0 1e-06 
3.0 1.833 0 3.0 1e-06 
0.05 1.834 0 3.0 1e-06 
3.0 1.834 0 3.0 1e-06 
0.05 1.835 0 3.0 1e-06 
3.0 1.835 0 3.0 1e-06 
0.05 1.836 0 3.0 1e-06 
3.0 1.836 0 3.0 1e-06 
0.05 1.837 0 3.0 1e-06 
3.0 1.837 0 3.0 1e-06 
0.05 1.838 0 3.0 1e-06 
3.0 1.838 0 3.0 1e-06 
0.05 1.839 0 3.0 1e-06 
3.0 1.839 0 3.0 1e-06 
0.05 1.84 0 3.0 1e-06 
3.0 1.84 0 3.0 1e-06 
0.05 1.841 0 3.0 1e-06 
3.0 1.841 0 3.0 1e-06 
0.05 1.842 0 3.0 1e-06 
3.0 1.842 0 3.0 1e-06 
0.05 1.843 0 3.0 1e-06 
3.0 1.843 0 3.0 1e-06 
0.05 1.844 0 3.0 1e-06 
3.0 1.844 0 3.0 1e-06 
0.05 1.845 0 3.0 1e-06 
3.0 1.845 0 3.0 1e-06 
0.05 1.846 0 3.0 1e-06 
3.0 1.846 0 3.0 1e-06 
0.05 1.847 0 3.0 1e-06 
3.0 1.847 0 3.0 1e-06 
0.05 1.848 0 3.0 1e-06 
3.0 1.848 0 3.0 1e-06 
0.05 1.849 0 3.0 1e-06 
3.0 1.849 0 3.0 1e-06 
0.05 1.85 0 3.0 1e-06 
3.0 1.85 0 3.0 1e-06 
0.05 1.851 0 3.0 1e-06 
3.0 1.851 0 3.0 1e-06 
0.05 1.852 0 3.0 1e-06 
3.0 1.852 0 3.0 1e-06 
0.05 1.853 0 3.0 1e-06 
3.0 1.853 0 3.0 1e-06 
0.05 1.854 0 3.0 1e-06 
3.0 1.854 0 3.0 1e-06 
0.05 1.855 0 3.0 1e-06 
3.0 1.855 0 3.0 1e-06 
0.05 1.856 0 3.0 1e-06 
3.0 1.856 0 3.0 1e-06 
0.05 1.857 0 3.0 1e-06 
3.0 1.857 0 3.0 1e-06 
0.05 1.858 0 3.0 1e-06 
3.0 1.858 0 3.0 1e-06 
0.05 1.859 0 3.0 1e-06 
3.0 1.859 0 3.0 1e-06 
0.05 1.86 0 3.0 1e-06 
3.0 1.86 0 3.0 1e-06 
0.05 1.861 0 3.0 1e-06 
3.0 1.861 0 3.0 1e-06 
0.05 1.862 0 3.0 1e-06 
3.0 1.862 0 3.0 1e-06 
0.05 1.863 0 3.0 1e-06 
3.0 1.863 0 3.0 1e-06 
0.05 1.864 0 3.0 1e-06 
3.0 1.864 0 3.0 1e-06 
0.05 1.865 0 3.0 1e-06 
3.0 1.865 0 3.0 1e-06 
0.05 1.866 0 3.0 1e-06 
3.0 1.866 0 3.0 1e-06 
0.05 1.867 0 3.0 1e-06 
3.0 1.867 0 3.0 1e-06 
0.05 1.868 0 3.0 1e-06 
3.0 1.868 0 3.0 1e-06 
0.05 1.869 0 3.0 1e-06 
3.0 1.869 0 3.0 1e-06 
0.05 1.87 0 3.0 1e-06 
3.0 1.87 0 3.0 1e-06 
0.05 1.871 0 3.0 1e-06 
3.0 1.871 0 3.0 1e-06 
0.05 1.872 0 3.0 1e-06 
3.0 1.872 0 3.0 1e-06 
0.05 1.873 0 3.0 1e-06 
3.0 1.873 0 3.0 1e-06 
0.05 1.874 0 3.0 1e-06 
3.0 1.874 0 3.0 1e-06 
0.05 1.875 0 3.0 1e-06 
3.0 1.875 0 3.0 1e-06 
0.05 1.876 0 3.0 1e-06 
3.0 1.876 0 3.0 1e-06 
0.05 1.877 0 3.0 1e-06 
3.0 1.877 0 3.0 1e-06 
0.05 1.878 0 3.0 1e-06 
3.0 1.878 0 3.0 1e-06 
0.05 1.879 0 3.0 1e-06 
3.0 1.879 0 3.0 1e-06 
0.05 1.88 0 3.0 1e-06 
3.0 1.88 0 3.0 1e-06 
0.05 1.881 0 3.0 1e-06 
3.0 1.881 0 3.0 1e-06 
0.05 1.882 0 3.0 1e-06 
3.0 1.882 0 3.0 1e-06 
0.05 1.883 0 3.0 1e-06 
3.0 1.883 0 3.0 1e-06 
0.05 1.884 0 3.0 1e-06 
3.0 1.884 0 3.0 1e-06 
0.05 1.885 0 3.0 1e-06 
3.0 1.885 0 3.0 1e-06 
0.05 1.886 0 3.0 1e-06 
3.0 1.886 0 3.0 1e-06 
0.05 1.887 0 3.0 1e-06 
3.0 1.887 0 3.0 1e-06 
0.05 1.888 0 3.0 1e-06 
3.0 1.888 0 3.0 1e-06 
0.05 1.889 0 3.0 1e-06 
3.0 1.889 0 3.0 1e-06 
0.05 1.89 0 3.0 1e-06 
3.0 1.89 0 3.0 1e-06 
0.05 1.891 0 3.0 1e-06 
3.0 1.891 0 3.0 1e-06 
0.05 1.892 0 3.0 1e-06 
3.0 1.892 0 3.0 1e-06 
0.05 1.893 0 3.0 1e-06 
3.0 1.893 0 3.0 1e-06 
0.05 1.894 0 3.0 1e-06 
3.0 1.894 0 3.0 1e-06 
0.05 1.895 0 3.0 1e-06 
3.0 1.895 0 3.0 1e-06 
0.05 1.896 0 3.0 1e-06 
3.0 1.896 0 3.0 1e-06 
0.05 1.897 0 3.0 1e-06 
3.0 1.897 0 3.0 1e-06 
0.05 1.898 0 3.0 1e-06 
3.0 1.898 0 3.0 1e-06 
0.05 1.899 0 3.0 1e-06 
3.0 1.899 0 3.0 1e-06 
0.05 1.9 0 3.0 1e-06 
3.0 1.9 0 3.0 1e-06 
0.05 1.901 0 3.0 1e-06 
3.0 1.901 0 3.0 1e-06 
0.05 1.902 0 3.0 1e-06 
3.0 1.902 0 3.0 1e-06 
0.05 1.903 0 3.0 1e-06 
3.0 1.903 0 3.0 1e-06 
0.05 1.904 0 3.0 1e-06 
3.0 1.904 0 3.0 1e-06 
0.05 1.905 0 3.0 1e-06 
3.0 1.905 0 3.0 1e-06 
0.05 1.906 0 3.0 1e-06 
3.0 1.906 0 3.0 1e-06 
0.05 1.907 0 3.0 1e-06 
3.0 1.907 0 3.0 1e-06 
0.05 1.908 0 3.0 1e-06 
3.0 1.908 0 3.0 1e-06 
0.05 1.909 0 3.0 1e-06 
3.0 1.909 0 3.0 1e-06 
0.05 1.91 0 3.0 1e-06 
3.0 1.91 0 3.0 1e-06 
0.05 1.911 0 3.0 1e-06 
3.0 1.911 0 3.0 1e-06 
0.05 1.912 0 3.0 1e-06 
3.0 1.912 0 3.0 1e-06 
0.05 1.913 0 3.0 1e-06 
3.0 1.913 0 3.0 1e-06 
0.05 1.914 0 3.0 1e-06 
3.0 1.914 0 3.0 1e-06 
0.05 1.915 0 3.0 1e-06 
3.0 1.915 0 3.0 1e-06 
0.05 1.916 0 3.0 1e-06 
3.0 1.916 0 3.0 1e-06 
0.05 1.917 0 3.0 1e-06 
3.0 1.917 0 3.0 1e-06 
0.05 1.918 0 3.0 1e-06 
3.0 1.918 0 3.0 1e-06 
0.05 1.919 0 3.0 1e-06 
3.0 1.919 0 3.0 1e-06 
0.05 1.92 0 3.0 1e-06 
3.0 1.92 0 3.0 1e-06 
0.05 1.921 0 3.0 1e-06 
3.0 1.921 0 3.0 1e-06 
0.05 1.922 0 3.0 1e-06 
3.0 1.922 0 3.0 1e-06 
0.05 1.923 0 3.0 1e-06 
3.0 1.923 0 3.0 1e-06 
0.05 1.924 0 3.0 1e-06 
3.0 1.924 0 3.0 1e-06 
0.05 1.925 0 3.0 1e-06 
3.0 1.925 0 3.0 1e-06 
0.05 1.926 0 3.0 1e-06 
3.0 1.926 0 3.0 1e-06 
0.05 1.927 0 3.0 1e-06 
3.0 1.927 0 3.0 1e-06 
0.05 1.928 0 3.0 1e-06 
3.0 1.928 0 3.0 1e-06 
0.05 1.929 0 3.0 1e-06 
3.0 1.929 0 3.0 1e-06 
0.05 1.93 0 3.0 1e-06 
3.0 1.93 0 3.0 1e-06 
0.05 1.931 0 3.0 1e-06 
3.0 1.931 0 3.0 1e-06 
0.05 1.932 0 3.0 1e-06 
3.0 1.932 0 3.0 1e-06 
0.05 1.933 0 3.0 1e-06 
3.0 1.933 0 3.0 1e-06 
0.05 1.934 0 3.0 1e-06 
3.0 1.934 0 3.0 1e-06 
0.05 1.935 0 3.0 1e-06 
3.0 1.935 0 3.0 1e-06 
0.05 1.936 0 3.0 1e-06 
3.0 1.936 0 3.0 1e-06 
0.05 1.937 0 3.0 1e-06 
3.0 1.937 0 3.0 1e-06 
0.05 1.938 0 3.0 1e-06 
3.0 1.938 0 3.0 1e-06 
0.05 1.939 0 3.0 1e-06 
3.0 1.939 0 3.0 1e-06 
0.05 1.94 0 3.0 1e-06 
3.0 1.94 0 3.0 1e-06 
0.05 1.941 0 3.0 1e-06 
3.0 1.941 0 3.0 1e-06 
0.05 1.942 0 3.0 1e-06 
3.0 1.942 0 3.0 1e-06 
0.05 1.943 0 3.0 1e-06 
3.0 1.943 0 3.0 1e-06 
0.05 1.944 0 3.0 1e-06 
3.0 1.944 0 3.0 1e-06 
0.05 1.945 0 3.0 1e-06 
3.0 1.945 0 3.0 1e-06 
0.05 1.946 0 3.0 1e-06 
3.0 1.946 0 3.0 1e-06 
0.05 1.947 0 3.0 1e-06 
3.0 1.947 0 3.0 1e-06 
0.05 1.948 0 3.0 1e-06 
3.0 1.948 0 3.0 1e-06 
0.05 1.949 0 3.0 1e-06 
3.0 1.949 0 3.0 1e-06 
0.05 1.95 0 3.0 1e-06 
3.0 1.95 0 3.0 1e-06 
0.05 1.951 0 3.0 1e-06 
3.0 1.951 0 3.0 1e-06 
0.05 1.952 0 3.0 1e-06 
3.0 1.952 0 3.0 1e-06 
0.05 1.953 0 3.0 1e-06 
3.0 1.953 0 3.0 1e-06 
0.05 1.954 0 3.0 1e-06 
3.0 1.954 0 3.0 1e-06 
0.05 1.955 0 3.0 1e-06 
3.0 1.955 0 3.0 1e-06 
0.05 1.956 0 3.0 1e-06 
3.0 1.956 0 3.0 1e-06 
0.05 1.957 0 3.0 1e-06 
3.0 1.957 0 3.0 1e-06 
0.05 1.958 0 3.0 1e-06 
3.0 1.958 0 3.0 1e-06 
0.05 1.959 0 3.0 1e-06 
3.0 1.959 0 3.0 1e-06 
0.05 1.96 0 3.0 1e-06 
3.0 1.96 0 3.0 1e-06 
0.05 1.961 0 3.0 1e-06 
3.0 1.961 0 3.0 1e-06 
0.05 1.962 0 3.0 1e-06 
3.0 1.962 0 3.0 1e-06 
0.05 1.963 0 3.0 1e-06 
3.0 1.963 0 3.0 1e-06 
0.05 1.964 0 3.0 1e-06 
3.0 1.964 0 3.0 1e-06 
0.05 1.965 0 3.0 1e-06 
3.0 1.965 0 3.0 1e-06 
0.05 1.966 0 3.0 1e-06 
3.0 1.966 0 3.0 1e-06 
0.05 1.967 0 3.0 1e-06 
3.0 1.967 0 3.0 1e-06 
0.05 1.968 0 3.0 1e-06 
3.0 1.968 0 3.0 1e-06 
0.05 1.969 0 3.0 1e-06 
3.0 1.969 0 3.0 1e-06 
0.05 1.97 0 3.0 1e-06 
3.0 1.97 0 3.0 1e-06 
0.05 1.971 0 3.0 1e-06 
3.0 1.971 0 3.0 1e-06 
0.05 1.972 0 3.0 1e-06 
3.0 1.972 0 3.0 1e-06 
0.05 1.973 0 3.0 1e-06 
3.0 1.973 0 3.0 1e-06 
0.05 1.974 0 3.0 1e-06 
3.0 1.974 0 3.0 1e-06 
0.05 1.975 0 3.0 1e-06 
3.0 1.975 0 3.0 1e-06 
0.05 1.976 0 3.0 1e-06 
3.0 1.976 0 3.0 1e-06 
0.05 1.977 0 3.0 1e-06 
3.0 1.977 0 3.0 1e-06 
0.05 1.978 0 3.0 1e-06 
3.0 1.978 0 3.0 1e-06 
0.05 1.979 0 3.0 1e-06 
3.0 1.979 0 3.0 1e-06 
0.05 1.98 0 3.0 1e-06 
3.0 1.98 0 3.0 1e-06 
0.05 1.981 0 3.0 1e-06 
3.0 1.981 0 3.0 1e-06 
0.05 1.982 0 3.0 1e-06 
3.0 1.982 0 3.0 1e-06 
0.05 1.983 0 3.0 1e-06 
3.0 1.983 0 3.0 1e-06 
0.05 1.984 0 3.0 1e-06 
3.0 1.984 0 3.0 1e-06 
0.05 1.985 0 3.0 1e-06 
3.0 1.985 0 3.0 1e-06 
0.05 1.986 0 3.0 1e-06 
3.0 1.986 0 3.0 1e-06 
0.05 1.987 0 3.0 1e-06 
3.0 1.987 0 3.0 1e-06 
0.05 1.988 0 3.0 1e-06 
3.0 1.988 0 3.0 1e-06 
0.05 1.989 0 3.0 1e-06 
3.0 1.989 0 3.0 1e-06 
0.05 1.99 0 3.0 1e-06 
3.0 1.99 0 3.0 1e-06 
0.05 1.991 0 3.0 1e-06 
3.0 1.991 0 3.0 1e-06 
0.05 1.992 0 3.0 1e-06 
3.0 1.992 0 3.0 1e-06 
0.05 1.993 0 3.0 1e-06 
3.0 1.993 0 3.0 1e-06 
0.05 1.994 0 3.0 1e-06 
3.0 1.994 0 3.0 1e-06 
0.05 1.995 0 3.0 1e-06 
3.0 1.995 0 3.0 1e-06 
0.05 1.996 0 3.0 1e-06 
3.0 1.996 0 3.0 1e-06 
0.05 1.997 0 3.0 1e-06 
3.0 1.997 0 3.0 1e-06 
0.05 1.998 0 3.0 1e-06 
3.0 1.998 0 3.0 1e-06 
0.05 1.999 0 3.0 1e-06 
3.0 1.999 0 3.0 1e-06 
0.05 2.0 0 3.0 1e-06 
3.0 2.0 0 3.0 1e-06 
0.05 2.001 0 3.0 1e-06 
3.0 2.001 0 3.0 1e-06 
0.05 2.002 0 3.0 1e-06 
3.0 2.002 0 3.0 1e-06 
0.05 2.003 0 3.0 1e-06 
3.0 2.003 0 3.0 1e-06 
0.05 2.004 0 3.0 1e-06 
3.0 2.004 0 3.0 1e-06 
0.05 2.005 0 3.0 1e-06 
3.0 2.005 0 3.0 1e-06 
0.05 2.006 0 3.0 1e-06 
3.0 2.006 0 3.0 1e-06 
0.05 2.007 0 3.0 1e-06 
3.0 2.007 0 3.0 1e-06 
0.05 2.008 0 3.0 1e-06 
3.0 2.008 0 3.0 1e-06 
0.05 2.009 0 3.0 1e-06 
3.0 2.009 0 3.0 1e-06 
0.05 2.01 0 3.0 1e-06 
3.0 2.01 0 3.0 1e-06 
0.05 2.011 0 3.0 1e-06 
3.0 2.011 0 3.0 1e-06 
0.05 2.012 0 3.0 1e-06 
3.0 2.012 0 3.0 1e-06 
0.05 2.013 0 3.0 1e-06 
3.0 2.013 0 3.0 1e-06 
0.05 2.014 0 3.0 1e-06 
3.0 2.014 0 3.0 1e-06 
0.05 2.015 0 3.0 1e-06 
3.0 2.015 0 3.0 1e-06 
0.05 2.016 0 3.0 1e-06 
3.0 2.016 0 3.0 1e-06 
0.05 2.017 0 3.0 1e-06 
3.0 2.017 0 3.0 1e-06 
0.05 2.018 0 3.0 1e-06 
3.0 2.018 0 3.0 1e-06 
0.05 2.019 0 3.0 1e-06 
3.0 2.019 0 3.0 1e-06 
0.05 2.02 0 3.0 1e-06 
3.0 2.02 0 3.0 1e-06 
0.05 2.021 0 3.0 1e-06 
3.0 2.021 0 3.0 1e-06 
0.05 2.022 0 3.0 1e-06 
3.0 2.022 0 3.0 1e-06 
0.05 2.023 0 3.0 1e-06 
3.0 2.023 0 3.0 1e-06 
0.05 2.024 0 3.0 1e-06 
3.0 2.024 0 3.0 1e-06 
0.05 2.025 0 3.0 1e-06 
3.0 2.025 0 3.0 1e-06 
0.05 2.026 0 3.0 1e-06 
3.0 2.026 0 3.0 1e-06 
0.05 2.027 0 3.0 1e-06 
3.0 2.027 0 3.0 1e-06 
0.05 2.028 0 3.0 1e-06 
3.0 2.028 0 3.0 1e-06 
0.05 2.029 0 3.0 1e-06 
3.0 2.029 0 3.0 1e-06 
0.05 2.03 0 3.0 1e-06 
3.0 2.03 0 3.0 1e-06 
0.05 2.031 0 3.0 1e-06 
3.0 2.031 0 3.0 1e-06 
0.05 2.032 0 3.0 1e-06 
3.0 2.032 0 3.0 1e-06 
0.05 2.033 0 3.0 1e-06 
3.0 2.033 0 3.0 1e-06 
0.05 2.034 0 3.0 1e-06 
3.0 2.034 0 3.0 1e-06 
0.05 2.035 0 3.0 1e-06 
3.0 2.035 0 3.0 1e-06 
0.05 2.036 0 3.0 1e-06 
3.0 2.036 0 3.0 1e-06 
0.05 2.037 0 3.0 1e-06 
3.0 2.037 0 3.0 1e-06 
0.05 2.038 0 3.0 1e-06 
3.0 2.038 0 3.0 1e-06 
0.05 2.039 0 3.0 1e-06 
3.0 2.039 0 3.0 1e-06 
0.05 2.04 0 3.0 1e-06 
3.0 2.04 0 3.0 1e-06 
0.05 2.041 0 3.0 1e-06 
3.0 2.041 0 3.0 1e-06 
0.05 2.042 0 3.0 1e-06 
3.0 2.042 0 3.0 1e-06 
0.05 2.043 0 3.0 1e-06 
3.0 2.043 0 3.0 1e-06 
0.05 2.044 0 3.0 1e-06 
3.0 2.044 0 3.0 1e-06 
0.05 2.045 0 3.0 1e-06 
3.0 2.045 0 3.0 1e-06 
0.05 2.046 0 3.0 1e-06 
3.0 2.046 0 3.0 1e-06 
0.05 2.047 0 3.0 1e-06 
3.0 2.047 0 3.0 1e-06 
0.05 2.048 0 3.0 1e-06 
3.0 2.048 0 3.0 1e-06 
0.05 2.049 0 3.0 1e-06 
3.0 2.049 0 3.0 1e-06 
0.05 2.05 0 3.0 1e-06 
3.0 2.05 0 3.0 1e-06 
0.05 2.051 0 3.0 1e-06 
3.0 2.051 0 3.0 1e-06 
0.05 2.052 0 3.0 1e-06 
3.0 2.052 0 3.0 1e-06 
0.05 2.053 0 3.0 1e-06 
3.0 2.053 0 3.0 1e-06 
0.05 2.054 0 3.0 1e-06 
3.0 2.054 0 3.0 1e-06 
0.05 2.055 0 3.0 1e-06 
3.0 2.055 0 3.0 1e-06 
0.05 2.056 0 3.0 1e-06 
3.0 2.056 0 3.0 1e-06 
0.05 2.057 0 3.0 1e-06 
3.0 2.057 0 3.0 1e-06 
0.05 2.058 0 3.0 1e-06 
3.0 2.058 0 3.0 1e-06 
0.05 2.059 0 3.0 1e-06 
3.0 2.059 0 3.0 1e-06 
0.05 2.06 0 3.0 1e-06 
3.0 2.06 0 3.0 1e-06 
0.05 2.061 0 3.0 1e-06 
3.0 2.061 0 3.0 1e-06 
0.05 2.062 0 3.0 1e-06 
3.0 2.062 0 3.0 1e-06 
0.05 2.063 0 3.0 1e-06 
3.0 2.063 0 3.0 1e-06 
0.05 2.064 0 3.0 1e-06 
3.0 2.064 0 3.0 1e-06 
0.05 2.065 0 3.0 1e-06 
3.0 2.065 0 3.0 1e-06 
0.05 2.066 0 3.0 1e-06 
3.0 2.066 0 3.0 1e-06 
0.05 2.067 0 3.0 1e-06 
3.0 2.067 0 3.0 1e-06 
0.05 2.068 0 3.0 1e-06 
3.0 2.068 0 3.0 1e-06 
0.05 2.069 0 3.0 1e-06 
3.0 2.069 0 3.0 1e-06 
0.05 2.07 0 3.0 1e-06 
3.0 2.07 0 3.0 1e-06 
0.05 2.071 0 3.0 1e-06 
3.0 2.071 0 3.0 1e-06 
0.05 2.072 0 3.0 1e-06 
3.0 2.072 0 3.0 1e-06 
0.05 2.073 0 3.0 1e-06 
3.0 2.073 0 3.0 1e-06 
0.05 2.074 0 3.0 1e-06 
3.0 2.074 0 3.0 1e-06 
0.05 2.075 0 3.0 1e-06 
3.0 2.075 0 3.0 1e-06 
0.05 2.076 0 3.0 1e-06 
3.0 2.076 0 3.0 1e-06 
0.05 2.077 0 3.0 1e-06 
3.0 2.077 0 3.0 1e-06 
0.05 2.078 0 3.0 1e-06 
3.0 2.078 0 3.0 1e-06 
0.05 2.079 0 3.0 1e-06 
3.0 2.079 0 3.0 1e-06 
0.05 2.08 0 3.0 1e-06 
3.0 2.08 0 3.0 1e-06 
0.05 2.081 0 3.0 1e-06 
3.0 2.081 0 3.0 1e-06 
0.05 2.082 0 3.0 1e-06 
3.0 2.082 0 3.0 1e-06 
0.05 2.083 0 3.0 1e-06 
3.0 2.083 0 3.0 1e-06 
0.05 2.084 0 3.0 1e-06 
3.0 2.084 0 3.0 1e-06 
0.05 2.085 0 3.0 1e-06 
3.0 2.085 0 3.0 1e-06 
0.05 2.086 0 3.0 1e-06 
3.0 2.086 0 3.0 1e-06 
0.05 2.087 0 3.0 1e-06 
3.0 2.087 0 3.0 1e-06 
0.05 2.088 0 3.0 1e-06 
3.0 2.088 0 3.0 1e-06 
0.05 2.089 0 3.0 1e-06 
3.0 2.089 0 3.0 1e-06 
0.05 2.09 0 3.0 1e-06 
3.0 2.09 0 3.0 1e-06 
0.05 2.091 0 3.0 1e-06 
3.0 2.091 0 3.0 1e-06 
0.05 2.092 0 3.0 1e-06 
3.0 2.092 0 3.0 1e-06 
0.05 2.093 0 3.0 1e-06 
3.0 2.093 0 3.0 1e-06 
0.05 2.094 0 3.0 1e-06 
3.0 2.094 0 3.0 1e-06 
0.05 2.095 0 3.0 1e-06 
3.0 2.095 0 3.0 1e-06 
0.05 2.096 0 3.0 1e-06 
3.0 2.096 0 3.0 1e-06 
0.05 2.097 0 3.0 1e-06 
3.0 2.097 0 3.0 1e-06 
0.05 2.098 0 3.0 1e-06 
3.0 2.098 0 3.0 1e-06 
0.05 2.099 0 3.0 1e-06 
3.0 2.099 0 3.0 1e-06 
0.05 2.1 0 3.0 1e-06 
3.0 2.1 0 3.0 1e-06 
0.05 2.101 0 3.0 1e-06 
3.0 2.101 0 3.0 1e-06 
0.05 2.102 0 3.0 1e-06 
3.0 2.102 0 3.0 1e-06 
0.05 2.103 0 3.0 1e-06 
3.0 2.103 0 3.0 1e-06 
0.05 2.104 0 3.0 1e-06 
3.0 2.104 0 3.0 1e-06 
0.05 2.105 0 3.0 1e-06 
3.0 2.105 0 3.0 1e-06 
0.05 2.106 0 3.0 1e-06 
3.0 2.106 0 3.0 1e-06 
0.05 2.107 0 3.0 1e-06 
3.0 2.107 0 3.0 1e-06 
0.05 2.108 0 3.0 1e-06 
3.0 2.108 0 3.0 1e-06 
0.05 2.109 0 3.0 1e-06 
3.0 2.109 0 3.0 1e-06 
0.05 2.11 0 3.0 1e-06 
3.0 2.11 0 3.0 1e-06 
0.05 2.111 0 3.0 1e-06 
3.0 2.111 0 3.0 1e-06 
0.05 2.112 0 3.0 1e-06 
3.0 2.112 0 3.0 1e-06 
0.05 2.113 0 3.0 1e-06 
3.0 2.113 0 3.0 1e-06 
0.05 2.114 0 3.0 1e-06 
3.0 2.114 0 3.0 1e-06 
0.05 2.115 0 3.0 1e-06 
3.0 2.115 0 3.0 1e-06 
0.05 2.116 0 3.0 1e-06 
3.0 2.116 0 3.0 1e-06 
0.05 2.117 0 3.0 1e-06 
3.0 2.117 0 3.0 1e-06 
0.05 2.118 0 3.0 1e-06 
3.0 2.118 0 3.0 1e-06 
0.05 2.119 0 3.0 1e-06 
3.0 2.119 0 3.0 1e-06 
0.05 2.12 0 3.0 1e-06 
3.0 2.12 0 3.0 1e-06 
0.05 2.121 0 3.0 1e-06 
3.0 2.121 0 3.0 1e-06 
0.05 2.122 0 3.0 1e-06 
3.0 2.122 0 3.0 1e-06 
0.05 2.123 0 3.0 1e-06 
3.0 2.123 0 3.0 1e-06 
0.05 2.124 0 3.0 1e-06 
3.0 2.124 0 3.0 1e-06 
0.05 2.125 0 3.0 1e-06 
3.0 2.125 0 3.0 1e-06 
0.05 2.126 0 3.0 1e-06 
3.0 2.126 0 3.0 1e-06 
0.05 2.127 0 3.0 1e-06 
3.0 2.127 0 3.0 1e-06 
0.05 2.128 0 3.0 1e-06 
3.0 2.128 0 3.0 1e-06 
0.05 2.129 0 3.0 1e-06 
3.0 2.129 0 3.0 1e-06 
0.05 2.13 0 3.0 1e-06 
3.0 2.13 0 3.0 1e-06 
0.05 2.131 0 3.0 1e-06 
3.0 2.131 0 3.0 1e-06 
0.05 2.132 0 3.0 1e-06 
3.0 2.132 0 3.0 1e-06 
0.05 2.133 0 3.0 1e-06 
3.0 2.133 0 3.0 1e-06 
0.05 2.134 0 3.0 1e-06 
3.0 2.134 0 3.0 1e-06 
0.05 2.135 0 3.0 1e-06 
3.0 2.135 0 3.0 1e-06 
0.05 2.136 0 3.0 1e-06 
3.0 2.136 0 3.0 1e-06 
0.05 2.137 0 3.0 1e-06 
3.0 2.137 0 3.0 1e-06 
0.05 2.138 0 3.0 1e-06 
3.0 2.138 0 3.0 1e-06 
0.05 2.139 0 3.0 1e-06 
3.0 2.139 0 3.0 1e-06 
0.05 2.14 0 3.0 1e-06 
3.0 2.14 0 3.0 1e-06 
0.05 2.141 0 3.0 1e-06 
3.0 2.141 0 3.0 1e-06 
0.05 2.142 0 3.0 1e-06 
3.0 2.142 0 3.0 1e-06 
0.05 2.143 0 3.0 1e-06 
3.0 2.143 0 3.0 1e-06 
0.05 2.144 0 3.0 1e-06 
3.0 2.144 0 3.0 1e-06 
0.05 2.145 0 3.0 1e-06 
3.0 2.145 0 3.0 1e-06 
0.05 2.146 0 3.0 1e-06 
3.0 2.146 0 3.0 1e-06 
0.05 2.147 0 3.0 1e-06 
3.0 2.147 0 3.0 1e-06 
0.05 2.148 0 3.0 1e-06 
3.0 2.148 0 3.0 1e-06 
0.05 2.149 0 3.0 1e-06 
3.0 2.149 0 3.0 1e-06 
0.05 2.15 0 3.0 1e-06 
3.0 2.15 0 3.0 1e-06 
0.05 2.151 0 3.0 1e-06 
3.0 2.151 0 3.0 1e-06 
0.05 2.152 0 3.0 1e-06 
3.0 2.152 0 3.0 1e-06 
0.05 2.153 0 3.0 1e-06 
3.0 2.153 0 3.0 1e-06 
0.05 2.154 0 3.0 1e-06 
3.0 2.154 0 3.0 1e-06 
0.05 2.155 0 3.0 1e-06 
3.0 2.155 0 3.0 1e-06 
0.05 2.156 0 3.0 1e-06 
3.0 2.156 0 3.0 1e-06 
0.05 2.157 0 3.0 1e-06 
3.0 2.157 0 3.0 1e-06 
0.05 2.158 0 3.0 1e-06 
3.0 2.158 0 3.0 1e-06 
0.05 2.159 0 3.0 1e-06 
3.0 2.159 0 3.0 1e-06 
0.05 2.16 0 3.0 1e-06 
3.0 2.16 0 3.0 1e-06 
0.05 2.161 0 3.0 1e-06 
3.0 2.161 0 3.0 1e-06 
0.05 2.162 0 3.0 1e-06 
3.0 2.162 0 3.0 1e-06 
0.05 2.163 0 3.0 1e-06 
3.0 2.163 0 3.0 1e-06 
0.05 2.164 0 3.0 1e-06 
3.0 2.164 0 3.0 1e-06 
0.05 2.165 0 3.0 1e-06 
3.0 2.165 0 3.0 1e-06 
0.05 2.166 0 3.0 1e-06 
3.0 2.166 0 3.0 1e-06 
0.05 2.167 0 3.0 1e-06 
3.0 2.167 0 3.0 1e-06 
0.05 2.168 0 3.0 1e-06 
3.0 2.168 0 3.0 1e-06 
0.05 2.169 0 3.0 1e-06 
3.0 2.169 0 3.0 1e-06 
0.05 2.17 0 3.0 1e-06 
3.0 2.17 0 3.0 1e-06 
0.05 2.171 0 3.0 1e-06 
3.0 2.171 0 3.0 1e-06 
0.05 2.172 0 3.0 1e-06 
3.0 2.172 0 3.0 1e-06 
0.05 2.173 0 3.0 1e-06 
3.0 2.173 0 3.0 1e-06 
0.05 2.174 0 3.0 1e-06 
3.0 2.174 0 3.0 1e-06 
0.05 2.175 0 3.0 1e-06 
3.0 2.175 0 3.0 1e-06 
0.05 2.176 0 3.0 1e-06 
3.0 2.176 0 3.0 1e-06 
0.05 2.177 0 3.0 1e-06 
3.0 2.177 0 3.0 1e-06 
0.05 2.178 0 3.0 1e-06 
3.0 2.178 0 3.0 1e-06 
0.05 2.179 0 3.0 1e-06 
3.0 2.179 0 3.0 1e-06 
0.05 2.18 0 3.0 1e-06 
3.0 2.18 0 3.0 1e-06 
0.05 2.181 0 3.0 1e-06 
3.0 2.181 0 3.0 1e-06 
0.05 2.182 0 3.0 1e-06 
3.0 2.182 0 3.0 1e-06 
0.05 2.183 0 3.0 1e-06 
3.0 2.183 0 3.0 1e-06 
0.05 2.184 0 3.0 1e-06 
3.0 2.184 0 3.0 1e-06 
0.05 2.185 0 3.0 1e-06 
3.0 2.185 0 3.0 1e-06 
0.05 2.186 0 3.0 1e-06 
3.0 2.186 0 3.0 1e-06 
0.05 2.187 0 3.0 1e-06 
3.0 2.187 0 3.0 1e-06 
0.05 2.188 0 3.0 1e-06 
3.0 2.188 0 3.0 1e-06 
0.05 2.189 0 3.0 1e-06 
3.0 2.189 0 3.0 1e-06 
0.05 2.19 0 3.0 1e-06 
3.0 2.19 0 3.0 1e-06 
0.05 2.191 0 3.0 1e-06 
3.0 2.191 0 3.0 1e-06 
0.05 2.192 0 3.0 1e-06 
3.0 2.192 0 3.0 1e-06 
0.05 2.193 0 3.0 1e-06 
3.0 2.193 0 3.0 1e-06 
0.05 2.194 0 3.0 1e-06 
3.0 2.194 0 3.0 1e-06 
0.05 2.195 0 3.0 1e-06 
3.0 2.195 0 3.0 1e-06 
0.05 2.196 0 3.0 1e-06 
3.0 2.196 0 3.0 1e-06 
0.05 2.197 0 3.0 1e-06 
3.0 2.197 0 3.0 1e-06 
0.05 2.198 0 3.0 1e-06 
3.0 2.198 0 3.0 1e-06 
0.05 2.199 0 3.0 1e-06 
3.0 2.199 0 3.0 1e-06 
0.05 2.2 0 3.0 1e-06 
3.0 2.2 0 3.0 1e-06 
0.05 2.201 0 3.0 1e-06 
3.0 2.201 0 3.0 1e-06 
0.05 2.202 0 3.0 1e-06 
3.0 2.202 0 3.0 1e-06 
0.05 2.203 0 3.0 1e-06 
3.0 2.203 0 3.0 1e-06 
0.05 2.204 0 3.0 1e-06 
3.0 2.204 0 3.0 1e-06 
0.05 2.205 0 3.0 1e-06 
3.0 2.205 0 3.0 1e-06 
0.05 2.206 0 3.0 1e-06 
3.0 2.206 0 3.0 1e-06 
0.05 2.207 0 3.0 1e-06 
3.0 2.207 0 3.0 1e-06 
0.05 2.208 0 3.0 1e-06 
3.0 2.208 0 3.0 1e-06 
0.05 2.209 0 3.0 1e-06 
3.0 2.209 0 3.0 1e-06 
0.05 2.21 0 3.0 1e-06 
3.0 2.21 0 3.0 1e-06 
0.05 2.211 0 3.0 1e-06 
3.0 2.211 0 3.0 1e-06 
0.05 2.212 0 3.0 1e-06 
3.0 2.212 0 3.0 1e-06 
0.05 2.213 0 3.0 1e-06 
3.0 2.213 0 3.0 1e-06 
0.05 2.214 0 3.0 1e-06 
3.0 2.214 0 3.0 1e-06 
0.05 2.215 0 3.0 1e-06 
3.0 2.215 0 3.0 1e-06 
0.05 2.216 0 3.0 1e-06 
3.0 2.216 0 3.0 1e-06 
0.05 2.217 0 3.0 1e-06 
3.0 2.217 0 3.0 1e-06 
0.05 2.218 0 3.0 1e-06 
3.0 2.218 0 3.0 1e-06 
0.05 2.219 0 3.0 1e-06 
3.0 2.219 0 3.0 1e-06 
0.05 2.22 0 3.0 1e-06 
3.0 2.22 0 3.0 1e-06 
0.05 2.221 0 3.0 1e-06 
3.0 2.221 0 3.0 1e-06 
0.05 2.222 0 3.0 1e-06 
3.0 2.222 0 3.0 1e-06 
0.05 2.223 0 3.0 1e-06 
3.0 2.223 0 3.0 1e-06 
0.05 2.224 0 3.0 1e-06 
3.0 2.224 0 3.0 1e-06 
0.05 2.225 0 3.0 1e-06 
3.0 2.225 0 3.0 1e-06 
0.05 2.226 0 3.0 1e-06 
3.0 2.226 0 3.0 1e-06 
0.05 2.227 0 3.0 1e-06 
3.0 2.227 0 3.0 1e-06 
0.05 2.228 0 3.0 1e-06 
3.0 2.228 0 3.0 1e-06 
0.05 2.229 0 3.0 1e-06 
3.0 2.229 0 3.0 1e-06 
0.05 2.23 0 3.0 1e-06 
3.0 2.23 0 3.0 1e-06 
0.05 2.231 0 3.0 1e-06 
3.0 2.231 0 3.0 1e-06 
0.05 2.232 0 3.0 1e-06 
3.0 2.232 0 3.0 1e-06 
0.05 2.233 0 3.0 1e-06 
3.0 2.233 0 3.0 1e-06 
0.05 2.234 0 3.0 1e-06 
3.0 2.234 0 3.0 1e-06 
0.05 2.235 0 3.0 1e-06 
3.0 2.235 0 3.0 1e-06 
0.05 2.236 0 3.0 1e-06 
3.0 2.236 0 3.0 1e-06 
0.05 2.237 0 3.0 1e-06 
3.0 2.237 0 3.0 1e-06 
0.05 2.238 0 3.0 1e-06 
3.0 2.238 0 3.0 1e-06 
0.05 2.239 0 3.0 1e-06 
3.0 2.239 0 3.0 1e-06 
0.05 2.24 0 3.0 1e-06 
3.0 2.24 0 3.0 1e-06 
0.05 2.241 0 3.0 1e-06 
3.0 2.241 0 3.0 1e-06 
0.05 2.242 0 3.0 1e-06 
3.0 2.242 0 3.0 1e-06 
0.05 2.243 0 3.0 1e-06 
3.0 2.243 0 3.0 1e-06 
0.05 2.244 0 3.0 1e-06 
3.0 2.244 0 3.0 1e-06 
0.05 2.245 0 3.0 1e-06 
3.0 2.245 0 3.0 1e-06 
0.05 2.246 0 3.0 1e-06 
3.0 2.246 0 3.0 1e-06 
0.05 2.247 0 3.0 1e-06 
3.0 2.247 0 3.0 1e-06 
0.05 2.248 0 3.0 1e-06 
3.0 2.248 0 3.0 1e-06 
0.05 2.249 0 3.0 1e-06 
3.0 2.249 0 3.0 1e-06 
0.05 2.25 0 3.0 1e-06 
3.0 2.25 0 3.0 1e-06 
0.05 2.251 0 3.0 1e-06 
3.0 2.251 0 3.0 1e-06 
0.05 2.252 0 3.0 1e-06 
3.0 2.252 0 3.0 1e-06 
0.05 2.253 0 3.0 1e-06 
3.0 2.253 0 3.0 1e-06 
0.05 2.254 0 3.0 1e-06 
3.0 2.254 0 3.0 1e-06 
0.05 2.255 0 3.0 1e-06 
3.0 2.255 0 3.0 1e-06 
0.05 2.256 0 3.0 1e-06 
3.0 2.256 0 3.0 1e-06 
0.05 2.257 0 3.0 1e-06 
3.0 2.257 0 3.0 1e-06 
0.05 2.258 0 3.0 1e-06 
3.0 2.258 0 3.0 1e-06 
0.05 2.259 0 3.0 1e-06 
3.0 2.259 0 3.0 1e-06 
0.05 2.26 0 3.0 1e-06 
3.0 2.26 0 3.0 1e-06 
0.05 2.261 0 3.0 1e-06 
3.0 2.261 0 3.0 1e-06 
0.05 2.262 0 3.0 1e-06 
3.0 2.262 0 3.0 1e-06 
0.05 2.263 0 3.0 1e-06 
3.0 2.263 0 3.0 1e-06 
0.05 2.264 0 3.0 1e-06 
3.0 2.264 0 3.0 1e-06 
0.05 2.265 0 3.0 1e-06 
3.0 2.265 0 3.0 1e-06 
0.05 2.266 0 3.0 1e-06 
3.0 2.266 0 3.0 1e-06 
0.05 2.267 0 3.0 1e-06 
3.0 2.267 0 3.0 1e-06 
0.05 2.268 0 3.0 1e-06 
3.0 2.268 0 3.0 1e-06 
0.05 2.269 0 3.0 1e-06 
3.0 2.269 0 3.0 1e-06 
0.05 2.27 0 3.0 1e-06 
3.0 2.27 0 3.0 1e-06 
0.05 2.271 0 3.0 1e-06 
3.0 2.271 0 3.0 1e-06 
0.05 2.272 0 3.0 1e-06 
3.0 2.272 0 3.0 1e-06 
0.05 2.273 0 3.0 1e-06 
3.0 2.273 0 3.0 1e-06 
0.05 2.274 0 3.0 1e-06 
3.0 2.274 0 3.0 1e-06 
0.05 2.275 0 3.0 1e-06 
3.0 2.275 0 3.0 1e-06 
0.05 2.276 0 3.0 1e-06 
3.0 2.276 0 3.0 1e-06 
0.05 2.277 0 3.0 1e-06 
3.0 2.277 0 3.0 1e-06 
0.05 2.278 0 3.0 1e-06 
3.0 2.278 0 3.0 1e-06 
0.05 2.279 0 3.0 1e-06 
3.0 2.279 0 3.0 1e-06 
0.05 2.28 0 3.0 1e-06 
3.0 2.28 0 3.0 1e-06 
0.05 2.281 0 3.0 1e-06 
3.0 2.281 0 3.0 1e-06 
0.05 2.282 0 3.0 1e-06 
3.0 2.282 0 3.0 1e-06 
0.05 2.283 0 3.0 1e-06 
3.0 2.283 0 3.0 1e-06 
0.05 2.284 0 3.0 1e-06 
3.0 2.284 0 3.0 1e-06 
0.05 2.285 0 3.0 1e-06 
3.0 2.285 0 3.0 1e-06 
0.05 2.286 0 3.0 1e-06 
3.0 2.286 0 3.0 1e-06 
0.05 2.287 0 3.0 1e-06 
3.0 2.287 0 3.0 1e-06 
0.05 2.288 0 3.0 1e-06 
3.0 2.288 0 3.0 1e-06 
0.05 2.289 0 3.0 1e-06 
3.0 2.289 0 3.0 1e-06 
0.05 2.29 0 3.0 1e-06 
3.0 2.29 0 3.0 1e-06 
0.05 2.291 0 3.0 1e-06 
3.0 2.291 0 3.0 1e-06 
0.05 2.292 0 3.0 1e-06 
3.0 2.292 0 3.0 1e-06 
0.05 2.293 0 3.0 1e-06 
3.0 2.293 0 3.0 1e-06 
0.05 2.294 0 3.0 1e-06 
3.0 2.294 0 3.0 1e-06 
0.05 2.295 0 3.0 1e-06 
3.0 2.295 0 3.0 1e-06 
0.05 2.296 0 3.0 1e-06 
3.0 2.296 0 3.0 1e-06 
0.05 2.297 0 3.0 1e-06 
3.0 2.297 0 3.0 1e-06 
0.05 2.298 0 3.0 1e-06 
3.0 2.298 0 3.0 1e-06 
0.05 2.299 0 3.0 1e-06 
3.0 2.299 0 3.0 1e-06 
0.05 2.3 0 3.0 1e-06 
3.0 2.3 0 3.0 1e-06 
0.05 2.301 0 3.0 1e-06 
3.0 2.301 0 3.0 1e-06 
0.05 2.302 0 3.0 1e-06 
3.0 2.302 0 3.0 1e-06 
0.05 2.303 0 3.0 1e-06 
3.0 2.303 0 3.0 1e-06 
0.05 2.304 0 3.0 1e-06 
3.0 2.304 0 3.0 1e-06 
0.05 2.305 0 3.0 1e-06 
3.0 2.305 0 3.0 1e-06 
0.05 2.306 0 3.0 1e-06 
3.0 2.306 0 3.0 1e-06 
0.05 2.307 0 3.0 1e-06 
3.0 2.307 0 3.0 1e-06 
0.05 2.308 0 3.0 1e-06 
3.0 2.308 0 3.0 1e-06 
0.05 2.309 0 3.0 1e-06 
3.0 2.309 0 3.0 1e-06 
0.05 2.31 0 3.0 1e-06 
3.0 2.31 0 3.0 1e-06 
0.05 2.311 0 3.0 1e-06 
3.0 2.311 0 3.0 1e-06 
0.05 2.312 0 3.0 1e-06 
3.0 2.312 0 3.0 1e-06 
0.05 2.313 0 3.0 1e-06 
3.0 2.313 0 3.0 1e-06 
0.05 2.314 0 3.0 1e-06 
3.0 2.314 0 3.0 1e-06 
0.05 2.315 0 3.0 1e-06 
3.0 2.315 0 3.0 1e-06 
0.05 2.316 0 3.0 1e-06 
3.0 2.316 0 3.0 1e-06 
0.05 2.317 0 3.0 1e-06 
3.0 2.317 0 3.0 1e-06 
0.05 2.318 0 3.0 1e-06 
3.0 2.318 0 3.0 1e-06 
0.05 2.319 0 3.0 1e-06 
3.0 2.319 0 3.0 1e-06 
0.05 2.32 0 3.0 1e-06 
3.0 2.32 0 3.0 1e-06 
0.05 2.321 0 3.0 1e-06 
3.0 2.321 0 3.0 1e-06 
0.05 2.322 0 3.0 1e-06 
3.0 2.322 0 3.0 1e-06 
0.05 2.323 0 3.0 1e-06 
3.0 2.323 0 3.0 1e-06 
0.05 2.324 0 3.0 1e-06 
3.0 2.324 0 3.0 1e-06 
0.05 2.325 0 3.0 1e-06 
3.0 2.325 0 3.0 1e-06 
0.05 2.326 0 3.0 1e-06 
3.0 2.326 0 3.0 1e-06 
0.05 2.327 0 3.0 1e-06 
3.0 2.327 0 3.0 1e-06 
0.05 2.328 0 3.0 1e-06 
3.0 2.328 0 3.0 1e-06 
0.05 2.329 0 3.0 1e-06 
3.0 2.329 0 3.0 1e-06 
0.05 2.33 0 3.0 1e-06 
3.0 2.33 0 3.0 1e-06 
0.05 2.331 0 3.0 1e-06 
3.0 2.331 0 3.0 1e-06 
0.05 2.332 0 3.0 1e-06 
3.0 2.332 0 3.0 1e-06 
0.05 2.333 0 3.0 1e-06 
3.0 2.333 0 3.0 1e-06 
0.05 2.334 0 3.0 1e-06 
3.0 2.334 0 3.0 1e-06 
0.05 2.335 0 3.0 1e-06 
3.0 2.335 0 3.0 1e-06 
0.05 2.336 0 3.0 1e-06 
3.0 2.336 0 3.0 1e-06 
0.05 2.337 0 3.0 1e-06 
3.0 2.337 0 3.0 1e-06 
0.05 2.338 0 3.0 1e-06 
3.0 2.338 0 3.0 1e-06 
0.05 2.339 0 3.0 1e-06 
3.0 2.339 0 3.0 1e-06 
0.05 2.34 0 3.0 1e-06 
3.0 2.34 0 3.0 1e-06 
0.05 2.341 0 3.0 1e-06 
3.0 2.341 0 3.0 1e-06 
0.05 2.342 0 3.0 1e-06 
3.0 2.342 0 3.0 1e-06 
0.05 2.343 0 3.0 1e-06 
3.0 2.343 0 3.0 1e-06 
0.05 2.344 0 3.0 1e-06 
3.0 2.344 0 3.0 1e-06 
0.05 2.345 0 3.0 1e-06 
3.0 2.345 0 3.0 1e-06 
0.05 2.346 0 3.0 1e-06 
3.0 2.346 0 3.0 1e-06 
0.05 2.347 0 3.0 1e-06 
3.0 2.347 0 3.0 1e-06 
0.05 2.348 0 3.0 1e-06 
3.0 2.348 0 3.0 1e-06 
0.05 2.349 0 3.0 1e-06 
3.0 2.349 0 3.0 1e-06 
0.05 2.35 0 3.0 1e-06 
3.0 2.35 0 3.0 1e-06 
0.05 2.351 0 3.0 1e-06 
3.0 2.351 0 3.0 1e-06 
0.05 2.352 0 3.0 1e-06 
3.0 2.352 0 3.0 1e-06 
0.05 2.353 0 3.0 1e-06 
3.0 2.353 0 3.0 1e-06 
0.05 2.354 0 3.0 1e-06 
3.0 2.354 0 3.0 1e-06 
0.05 2.355 0 3.0 1e-06 
3.0 2.355 0 3.0 1e-06 
0.05 2.356 0 3.0 1e-06 
3.0 2.356 0 3.0 1e-06 
0.05 2.357 0 3.0 1e-06 
3.0 2.357 0 3.0 1e-06 
0.05 2.358 0 3.0 1e-06 
3.0 2.358 0 3.0 1e-06 
0.05 2.359 0 3.0 1e-06 
3.0 2.359 0 3.0 1e-06 
0.05 2.36 0 3.0 1e-06 
3.0 2.36 0 3.0 1e-06 
0.05 2.361 0 3.0 1e-06 
3.0 2.361 0 3.0 1e-06 
0.05 2.362 0 3.0 1e-06 
3.0 2.362 0 3.0 1e-06 
0.05 2.363 0 3.0 1e-06 
3.0 2.363 0 3.0 1e-06 
0.05 2.364 0 3.0 1e-06 
3.0 2.364 0 3.0 1e-06 
0.05 2.365 0 3.0 1e-06 
3.0 2.365 0 3.0 1e-06 
0.05 2.366 0 3.0 1e-06 
3.0 2.366 0 3.0 1e-06 
0.05 2.367 0 3.0 1e-06 
3.0 2.367 0 3.0 1e-06 
0.05 2.368 0 3.0 1e-06 
3.0 2.368 0 3.0 1e-06 
0.05 2.369 0 3.0 1e-06 
3.0 2.369 0 3.0 1e-06 
0.05 2.37 0 3.0 1e-06 
3.0 2.37 0 3.0 1e-06 
0.05 2.371 0 3.0 1e-06 
3.0 2.371 0 3.0 1e-06 
0.05 2.372 0 3.0 1e-06 
3.0 2.372 0 3.0 1e-06 
0.05 2.373 0 3.0 1e-06 
3.0 2.373 0 3.0 1e-06 
0.05 2.374 0 3.0 1e-06 
3.0 2.374 0 3.0 1e-06 
0.05 2.375 0 3.0 1e-06 
3.0 2.375 0 3.0 1e-06 
0.05 2.376 0 3.0 1e-06 
3.0 2.376 0 3.0 1e-06 
0.05 2.377 0 3.0 1e-06 
3.0 2.377 0 3.0 1e-06 
0.05 2.378 0 3.0 1e-06 
3.0 2.378 0 3.0 1e-06 
0.05 2.379 0 3.0 1e-06 
3.0 2.379 0 3.0 1e-06 
0.05 2.38 0 3.0 1e-06 
3.0 2.38 0 3.0 1e-06 
0.05 2.381 0 3.0 1e-06 
3.0 2.381 0 3.0 1e-06 
0.05 2.382 0 3.0 1e-06 
3.0 2.382 0 3.0 1e-06 
0.05 2.383 0 3.0 1e-06 
3.0 2.383 0 3.0 1e-06 
0.05 2.384 0 3.0 1e-06 
3.0 2.384 0 3.0 1e-06 
0.05 2.385 0 3.0 1e-06 
3.0 2.385 0 3.0 1e-06 
0.05 2.386 0 3.0 1e-06 
3.0 2.386 0 3.0 1e-06 
0.05 2.387 0 3.0 1e-06 
3.0 2.387 0 3.0 1e-06 
0.05 2.388 0 3.0 1e-06 
3.0 2.388 0 3.0 1e-06 
0.05 2.389 0 3.0 1e-06 
3.0 2.389 0 3.0 1e-06 
0.05 2.39 0 3.0 1e-06 
3.0 2.39 0 3.0 1e-06 
0.05 2.391 0 3.0 1e-06 
3.0 2.391 0 3.0 1e-06 
0.05 2.392 0 3.0 1e-06 
3.0 2.392 0 3.0 1e-06 
0.05 2.393 0 3.0 1e-06 
3.0 2.393 0 3.0 1e-06 
0.05 2.394 0 3.0 1e-06 
3.0 2.394 0 3.0 1e-06 
0.05 2.395 0 3.0 1e-06 
3.0 2.395 0 3.0 1e-06 
0.05 2.396 0 3.0 1e-06 
3.0 2.396 0 3.0 1e-06 
0.05 2.397 0 3.0 1e-06 
3.0 2.397 0 3.0 1e-06 
0.05 2.398 0 3.0 1e-06 
3.0 2.398 0 3.0 1e-06 
0.05 2.399 0 3.0 1e-06 
3.0 2.399 0 3.0 1e-06 
0.05 2.4 0 3.0 1e-06 
3.0 2.4 0 3.0 1e-06 
0.05 2.401 0 3.0 1e-06 
3.0 2.401 0 3.0 1e-06 
0.05 2.402 0 3.0 1e-06 
3.0 2.402 0 3.0 1e-06 
0.05 2.403 0 3.0 1e-06 
3.0 2.403 0 3.0 1e-06 
0.05 2.404 0 3.0 1e-06 
3.0 2.404 0 3.0 1e-06 
0.05 2.405 0 3.0 1e-06 
3.0 2.405 0 3.0 1e-06 
0.05 2.406 0 3.0 1e-06 
3.0 2.406 0 3.0 1e-06 
0.05 2.407 0 3.0 1e-06 
3.0 2.407 0 3.0 1e-06 
0.05 2.408 0 3.0 1e-06 
3.0 2.408 0 3.0 1e-06 
0.05 2.409 0 3.0 1e-06 
3.0 2.409 0 3.0 1e-06 
0.05 2.41 0 3.0 1e-06 
3.0 2.41 0 3.0 1e-06 
0.05 2.411 0 3.0 1e-06 
3.0 2.411 0 3.0 1e-06 
0.05 2.412 0 3.0 1e-06 
3.0 2.412 0 3.0 1e-06 
0.05 2.413 0 3.0 1e-06 
3.0 2.413 0 3.0 1e-06 
0.05 2.414 0 3.0 1e-06 
3.0 2.414 0 3.0 1e-06 
0.05 2.415 0 3.0 1e-06 
3.0 2.415 0 3.0 1e-06 
0.05 2.416 0 3.0 1e-06 
3.0 2.416 0 3.0 1e-06 
0.05 2.417 0 3.0 1e-06 
3.0 2.417 0 3.0 1e-06 
0.05 2.418 0 3.0 1e-06 
3.0 2.418 0 3.0 1e-06 
0.05 2.419 0 3.0 1e-06 
3.0 2.419 0 3.0 1e-06 
0.05 2.42 0 3.0 1e-06 
3.0 2.42 0 3.0 1e-06 
0.05 2.421 0 3.0 1e-06 
3.0 2.421 0 3.0 1e-06 
0.05 2.422 0 3.0 1e-06 
3.0 2.422 0 3.0 1e-06 
0.05 2.423 0 3.0 1e-06 
3.0 2.423 0 3.0 1e-06 
0.05 2.424 0 3.0 1e-06 
3.0 2.424 0 3.0 1e-06 
0.05 2.425 0 3.0 1e-06 
3.0 2.425 0 3.0 1e-06 
0.05 2.426 0 3.0 1e-06 
3.0 2.426 0 3.0 1e-06 
0.05 2.427 0 3.0 1e-06 
3.0 2.427 0 3.0 1e-06 
0.05 2.428 0 3.0 1e-06 
3.0 2.428 0 3.0 1e-06 
0.05 2.429 0 3.0 1e-06 
3.0 2.429 0 3.0 1e-06 
0.05 2.43 0 3.0 1e-06 
3.0 2.43 0 3.0 1e-06 
0.05 2.431 0 3.0 1e-06 
3.0 2.431 0 3.0 1e-06 
0.05 2.432 0 3.0 1e-06 
3.0 2.432 0 3.0 1e-06 
0.05 2.433 0 3.0 1e-06 
3.0 2.433 0 3.0 1e-06 
0.05 2.434 0 3.0 1e-06 
3.0 2.434 0 3.0 1e-06 
0.05 2.435 0 3.0 1e-06 
3.0 2.435 0 3.0 1e-06 
0.05 2.436 0 3.0 1e-06 
3.0 2.436 0 3.0 1e-06 
0.05 2.437 0 3.0 1e-06 
3.0 2.437 0 3.0 1e-06 
0.05 2.438 0 3.0 1e-06 
3.0 2.438 0 3.0 1e-06 
0.05 2.439 0 3.0 1e-06 
3.0 2.439 0 3.0 1e-06 
0.05 2.44 0 3.0 1e-06 
3.0 2.44 0 3.0 1e-06 
0.05 2.441 0 3.0 1e-06 
3.0 2.441 0 3.0 1e-06 
0.05 2.442 0 3.0 1e-06 
3.0 2.442 0 3.0 1e-06 
0.05 2.443 0 3.0 1e-06 
3.0 2.443 0 3.0 1e-06 
0.05 2.444 0 3.0 1e-06 
3.0 2.444 0 3.0 1e-06 
0.05 2.445 0 3.0 1e-06 
3.0 2.445 0 3.0 1e-06 
0.05 2.446 0 3.0 1e-06 
3.0 2.446 0 3.0 1e-06 
0.05 2.447 0 3.0 1e-06 
3.0 2.447 0 3.0 1e-06 
0.05 2.448 0 3.0 1e-06 
3.0 2.448 0 3.0 1e-06 
0.05 2.449 0 3.0 1e-06 
3.0 2.449 0 3.0 1e-06 
0.05 2.45 0 3.0 1e-06 
3.0 2.45 0 3.0 1e-06 
0.05 2.451 0 3.0 1e-06 
3.0 2.451 0 3.0 1e-06 
0.05 2.452 0 3.0 1e-06 
3.0 2.452 0 3.0 1e-06 
0.05 2.453 0 3.0 1e-06 
3.0 2.453 0 3.0 1e-06 
0.05 2.454 0 3.0 1e-06 
3.0 2.454 0 3.0 1e-06 
0.05 2.455 0 3.0 1e-06 
3.0 2.455 0 3.0 1e-06 
0.05 2.456 0 3.0 1e-06 
3.0 2.456 0 3.0 1e-06 
0.05 2.457 0 3.0 1e-06 
3.0 2.457 0 3.0 1e-06 
0.05 2.458 0 3.0 1e-06 
3.0 2.458 0 3.0 1e-06 
0.05 2.459 0 3.0 1e-06 
3.0 2.459 0 3.0 1e-06 
0.05 2.46 0 3.0 1e-06 
3.0 2.46 0 3.0 1e-06 
0.05 2.461 0 3.0 1e-06 
3.0 2.461 0 3.0 1e-06 
0.05 2.462 0 3.0 1e-06 
3.0 2.462 0 3.0 1e-06 
0.05 2.463 0 3.0 1e-06 
3.0 2.463 0 3.0 1e-06 
0.05 2.464 0 3.0 1e-06 
3.0 2.464 0 3.0 1e-06 
0.05 2.465 0 3.0 1e-06 
3.0 2.465 0 3.0 1e-06 
0.05 2.466 0 3.0 1e-06 
3.0 2.466 0 3.0 1e-06 
0.05 2.467 0 3.0 1e-06 
3.0 2.467 0 3.0 1e-06 
0.05 2.468 0 3.0 1e-06 
3.0 2.468 0 3.0 1e-06 
0.05 2.469 0 3.0 1e-06 
3.0 2.469 0 3.0 1e-06 
0.05 2.47 0 3.0 1e-06 
3.0 2.47 0 3.0 1e-06 
0.05 2.471 0 3.0 1e-06 
3.0 2.471 0 3.0 1e-06 
0.05 2.472 0 3.0 1e-06 
3.0 2.472 0 3.0 1e-06 
0.05 2.473 0 3.0 1e-06 
3.0 2.473 0 3.0 1e-06 
0.05 2.474 0 3.0 1e-06 
3.0 2.474 0 3.0 1e-06 
0.05 2.475 0 3.0 1e-06 
3.0 2.475 0 3.0 1e-06 
0.05 2.476 0 3.0 1e-06 
3.0 2.476 0 3.0 1e-06 
0.05 2.477 0 3.0 1e-06 
3.0 2.477 0 3.0 1e-06 
0.05 2.478 0 3.0 1e-06 
3.0 2.478 0 3.0 1e-06 
0.05 2.479 0 3.0 1e-06 
3.0 2.479 0 3.0 1e-06 
0.05 2.48 0 3.0 1e-06 
3.0 2.48 0 3.0 1e-06 
0.05 2.481 0 3.0 1e-06 
3.0 2.481 0 3.0 1e-06 
0.05 2.482 0 3.0 1e-06 
3.0 2.482 0 3.0 1e-06 
0.05 2.483 0 3.0 1e-06 
3.0 2.483 0 3.0 1e-06 
0.05 2.484 0 3.0 1e-06 
3.0 2.484 0 3.0 1e-06 
0.05 2.485 0 3.0 1e-06 
3.0 2.485 0 3.0 1e-06 
0.05 2.486 0 3.0 1e-06 
3.0 2.486 0 3.0 1e-06 
0.05 2.487 0 3.0 1e-06 
3.0 2.487 0 3.0 1e-06 
0.05 2.488 0 3.0 1e-06 
3.0 2.488 0 3.0 1e-06 
0.05 2.489 0 3.0 1e-06 
3.0 2.489 0 3.0 1e-06 
0.05 2.49 0 3.0 1e-06 
3.0 2.49 0 3.0 1e-06 
0.05 2.491 0 3.0 1e-06 
3.0 2.491 0 3.0 1e-06 
0.05 2.492 0 3.0 1e-06 
3.0 2.492 0 3.0 1e-06 
0.05 2.493 0 3.0 1e-06 
3.0 2.493 0 3.0 1e-06 
0.05 2.494 0 3.0 1e-06 
3.0 2.494 0 3.0 1e-06 
0.05 2.495 0 3.0 1e-06 
3.0 2.495 0 3.0 1e-06 
0.05 2.496 0 3.0 1e-06 
3.0 2.496 0 3.0 1e-06 
0.05 2.497 0 3.0 1e-06 
3.0 2.497 0 3.0 1e-06 
0.05 2.498 0 3.0 1e-06 
3.0 2.498 0 3.0 1e-06 
0.05 2.499 0 3.0 1e-06 
3.0 2.499 0 3.0 1e-06 
0.05 2.5 0 3.0 1e-06 
3.0 2.5 0 3.0 1e-06 
0.05 2.501 0 3.0 1e-06 
3.0 2.501 0 3.0 1e-06 
0.05 2.502 0 3.0 1e-06 
3.0 2.502 0 3.0 1e-06 
0.05 2.503 0 3.0 1e-06 
3.0 2.503 0 3.0 1e-06 
0.05 2.504 0 3.0 1e-06 
3.0 2.504 0 3.0 1e-06 
0.05 2.505 0 3.0 1e-06 
3.0 2.505 0 3.0 1e-06 
0.05 2.506 0 3.0 1e-06 
3.0 2.506 0 3.0 1e-06 
0.05 2.507 0 3.0 1e-06 
3.0 2.507 0 3.0 1e-06 
0.05 2.508 0 3.0 1e-06 
3.0 2.508 0 3.0 1e-06 
0.05 2.509 0 3.0 1e-06 
3.0 2.509 0 3.0 1e-06 
0.05 2.51 0 3.0 1e-06 
3.0 2.51 0 3.0 1e-06 
0.05 2.511 0 3.0 1e-06 
3.0 2.511 0 3.0 1e-06 
0.05 2.512 0 3.0 1e-06 
3.0 2.512 0 3.0 1e-06 
0.05 2.513 0 3.0 1e-06 
3.0 2.513 0 3.0 1e-06 
0.05 2.514 0 3.0 1e-06 
3.0 2.514 0 3.0 1e-06 
0.05 2.515 0 3.0 1e-06 
3.0 2.515 0 3.0 1e-06 
0.05 2.516 0 3.0 1e-06 
3.0 2.516 0 3.0 1e-06 
0.05 2.517 0 3.0 1e-06 
3.0 2.517 0 3.0 1e-06 
0.05 2.518 0 3.0 1e-06 
3.0 2.518 0 3.0 1e-06 
0.05 2.519 0 3.0 1e-06 
3.0 2.519 0 3.0 1e-06 
0.05 2.52 0 3.0 1e-06 
3.0 2.52 0 3.0 1e-06 
0.05 2.521 0 3.0 1e-06 
3.0 2.521 0 3.0 1e-06 
0.05 2.522 0 3.0 1e-06 
3.0 2.522 0 3.0 1e-06 
0.05 2.523 0 3.0 1e-06 
3.0 2.523 0 3.0 1e-06 
0.05 2.524 0 3.0 1e-06 
3.0 2.524 0 3.0 1e-06 
0.05 2.525 0 3.0 1e-06 
3.0 2.525 0 3.0 1e-06 
0.05 2.526 0 3.0 1e-06 
3.0 2.526 0 3.0 1e-06 
0.05 2.527 0 3.0 1e-06 
3.0 2.527 0 3.0 1e-06 
0.05 2.528 0 3.0 1e-06 
3.0 2.528 0 3.0 1e-06 
0.05 2.529 0 3.0 1e-06 
3.0 2.529 0 3.0 1e-06 
0.05 2.53 0 3.0 1e-06 
3.0 2.53 0 3.0 1e-06 
0.05 2.531 0 3.0 1e-06 
3.0 2.531 0 3.0 1e-06 
0.05 2.532 0 3.0 1e-06 
3.0 2.532 0 3.0 1e-06 
0.05 2.533 0 3.0 1e-06 
3.0 2.533 0 3.0 1e-06 
0.05 2.534 0 3.0 1e-06 
3.0 2.534 0 3.0 1e-06 
0.05 2.535 0 3.0 1e-06 
3.0 2.535 0 3.0 1e-06 
0.05 2.536 0 3.0 1e-06 
3.0 2.536 0 3.0 1e-06 
0.05 2.537 0 3.0 1e-06 
3.0 2.537 0 3.0 1e-06 
0.05 2.538 0 3.0 1e-06 
3.0 2.538 0 3.0 1e-06 
0.05 2.539 0 3.0 1e-06 
3.0 2.539 0 3.0 1e-06 
0.05 2.54 0 3.0 1e-06 
3.0 2.54 0 3.0 1e-06 
0.05 2.541 0 3.0 1e-06 
3.0 2.541 0 3.0 1e-06 
0.05 2.542 0 3.0 1e-06 
3.0 2.542 0 3.0 1e-06 
0.05 2.543 0 3.0 1e-06 
3.0 2.543 0 3.0 1e-06 
0.05 2.544 0 3.0 1e-06 
3.0 2.544 0 3.0 1e-06 
0.05 2.545 0 3.0 1e-06 
3.0 2.545 0 3.0 1e-06 
0.05 2.546 0 3.0 1e-06 
3.0 2.546 0 3.0 1e-06 
0.05 2.547 0 3.0 1e-06 
3.0 2.547 0 3.0 1e-06 
0.05 2.548 0 3.0 1e-06 
3.0 2.548 0 3.0 1e-06 
0.05 2.549 0 3.0 1e-06 
3.0 2.549 0 3.0 1e-06 
0.05 2.55 0 3.0 1e-06 
3.0 2.55 0 3.0 1e-06 
0.05 2.551 0 3.0 1e-06 
3.0 2.551 0 3.0 1e-06 
0.05 2.552 0 3.0 1e-06 
3.0 2.552 0 3.0 1e-06 
0.05 2.553 0 3.0 1e-06 
3.0 2.553 0 3.0 1e-06 
0.05 2.554 0 3.0 1e-06 
3.0 2.554 0 3.0 1e-06 
0.05 2.555 0 3.0 1e-06 
3.0 2.555 0 3.0 1e-06 
0.05 2.556 0 3.0 1e-06 
3.0 2.556 0 3.0 1e-06 
0.05 2.557 0 3.0 1e-06 
3.0 2.557 0 3.0 1e-06 
0.05 2.558 0 3.0 1e-06 
3.0 2.558 0 3.0 1e-06 
0.05 2.559 0 3.0 1e-06 
3.0 2.559 0 3.0 1e-06 
0.05 2.56 0 3.0 1e-06 
3.0 2.56 0 3.0 1e-06 
0.05 2.561 0 3.0 1e-06 
3.0 2.561 0 3.0 1e-06 
0.05 2.562 0 3.0 1e-06 
3.0 2.562 0 3.0 1e-06 
0.05 2.563 0 3.0 1e-06 
3.0 2.563 0 3.0 1e-06 
0.05 2.564 0 3.0 1e-06 
3.0 2.564 0 3.0 1e-06 
0.05 2.565 0 3.0 1e-06 
3.0 2.565 0 3.0 1e-06 
0.05 2.566 0 3.0 1e-06 
3.0 2.566 0 3.0 1e-06 
0.05 2.567 0 3.0 1e-06 
3.0 2.567 0 3.0 1e-06 
0.05 2.568 0 3.0 1e-06 
3.0 2.568 0 3.0 1e-06 
0.05 2.569 0 3.0 1e-06 
3.0 2.569 0 3.0 1e-06 
0.05 2.57 0 3.0 1e-06 
3.0 2.57 0 3.0 1e-06 
0.05 2.571 0 3.0 1e-06 
3.0 2.571 0 3.0 1e-06 
0.05 2.572 0 3.0 1e-06 
3.0 2.572 0 3.0 1e-06 
0.05 2.573 0 3.0 1e-06 
3.0 2.573 0 3.0 1e-06 
0.05 2.574 0 3.0 1e-06 
3.0 2.574 0 3.0 1e-06 
0.05 2.575 0 3.0 1e-06 
3.0 2.575 0 3.0 1e-06 
0.05 2.576 0 3.0 1e-06 
3.0 2.576 0 3.0 1e-06 
0.05 2.577 0 3.0 1e-06 
3.0 2.577 0 3.0 1e-06 
0.05 2.578 0 3.0 1e-06 
3.0 2.578 0 3.0 1e-06 
0.05 2.579 0 3.0 1e-06 
3.0 2.579 0 3.0 1e-06 
0.05 2.58 0 3.0 1e-06 
3.0 2.58 0 3.0 1e-06 
0.05 2.581 0 3.0 1e-06 
3.0 2.581 0 3.0 1e-06 
0.05 2.582 0 3.0 1e-06 
3.0 2.582 0 3.0 1e-06 
0.05 2.583 0 3.0 1e-06 
3.0 2.583 0 3.0 1e-06 
0.05 2.584 0 3.0 1e-06 
3.0 2.584 0 3.0 1e-06 
0.05 2.585 0 3.0 1e-06 
3.0 2.585 0 3.0 1e-06 
0.05 2.586 0 3.0 1e-06 
3.0 2.586 0 3.0 1e-06 
0.05 2.587 0 3.0 1e-06 
3.0 2.587 0 3.0 1e-06 
0.05 2.588 0 3.0 1e-06 
3.0 2.588 0 3.0 1e-06 
0.05 2.589 0 3.0 1e-06 
3.0 2.589 0 3.0 1e-06 
0.05 2.59 0 3.0 1e-06 
3.0 2.59 0 3.0 1e-06 
0.05 2.591 0 3.0 1e-06 
3.0 2.591 0 3.0 1e-06 
0.05 2.592 0 3.0 1e-06 
3.0 2.592 0 3.0 1e-06 
0.05 2.593 0 3.0 1e-06 
3.0 2.593 0 3.0 1e-06 
0.05 2.594 0 3.0 1e-06 
3.0 2.594 0 3.0 1e-06 
0.05 2.595 0 3.0 1e-06 
3.0 2.595 0 3.0 1e-06 
0.05 2.596 0 3.0 1e-06 
3.0 2.596 0 3.0 1e-06 
0.05 2.597 0 3.0 1e-06 
3.0 2.597 0 3.0 1e-06 
0.05 2.598 0 3.0 1e-06 
3.0 2.598 0 3.0 1e-06 
0.05 2.599 0 3.0 1e-06 
3.0 2.599 0 3.0 1e-06 
0.05 2.6 0 3.0 1e-06 
3.0 2.6 0 3.0 1e-06 
0.05 2.601 0 3.0 1e-06 
3.0 2.601 0 3.0 1e-06 
0.05 2.602 0 3.0 1e-06 
3.0 2.602 0 3.0 1e-06 
0.05 2.603 0 3.0 1e-06 
3.0 2.603 0 3.0 1e-06 
0.05 2.604 0 3.0 1e-06 
3.0 2.604 0 3.0 1e-06 
0.05 2.605 0 3.0 1e-06 
3.0 2.605 0 3.0 1e-06 
0.05 2.606 0 3.0 1e-06 
3.0 2.606 0 3.0 1e-06 
0.05 2.607 0 3.0 1e-06 
3.0 2.607 0 3.0 1e-06 
0.05 2.608 0 3.0 1e-06 
3.0 2.608 0 3.0 1e-06 
0.05 2.609 0 3.0 1e-06 
3.0 2.609 0 3.0 1e-06 
0.05 2.61 0 3.0 1e-06 
3.0 2.61 0 3.0 1e-06 
0.05 2.611 0 3.0 1e-06 
3.0 2.611 0 3.0 1e-06 
0.05 2.612 0 3.0 1e-06 
3.0 2.612 0 3.0 1e-06 
0.05 2.613 0 3.0 1e-06 
3.0 2.613 0 3.0 1e-06 
0.05 2.614 0 3.0 1e-06 
3.0 2.614 0 3.0 1e-06 
0.05 2.615 0 3.0 1e-06 
3.0 2.615 0 3.0 1e-06 
0.05 2.616 0 3.0 1e-06 
3.0 2.616 0 3.0 1e-06 
0.05 2.617 0 3.0 1e-06 
3.0 2.617 0 3.0 1e-06 
0.05 2.618 0 3.0 1e-06 
3.0 2.618 0 3.0 1e-06 
0.05 2.619 0 3.0 1e-06 
3.0 2.619 0 3.0 1e-06 
0.05 2.62 0 3.0 1e-06 
3.0 2.62 0 3.0 1e-06 
0.05 2.621 0 3.0 1e-06 
3.0 2.621 0 3.0 1e-06 
0.05 2.622 0 3.0 1e-06 
3.0 2.622 0 3.0 1e-06 
0.05 2.623 0 3.0 1e-06 
3.0 2.623 0 3.0 1e-06 
0.05 2.624 0 3.0 1e-06 
3.0 2.624 0 3.0 1e-06 
0.05 2.625 0 3.0 1e-06 
3.0 2.625 0 3.0 1e-06 
0.05 2.626 0 3.0 1e-06 
3.0 2.626 0 3.0 1e-06 
0.05 2.627 0 3.0 1e-06 
3.0 2.627 0 3.0 1e-06 
0.05 2.628 0 3.0 1e-06 
3.0 2.628 0 3.0 1e-06 
0.05 2.629 0 3.0 1e-06 
3.0 2.629 0 3.0 1e-06 
0.05 2.63 0 3.0 1e-06 
3.0 2.63 0 3.0 1e-06 
0.05 2.631 0 3.0 1e-06 
3.0 2.631 0 3.0 1e-06 
0.05 2.632 0 3.0 1e-06 
3.0 2.632 0 3.0 1e-06 
0.05 2.633 0 3.0 1e-06 
3.0 2.633 0 3.0 1e-06 
0.05 2.634 0 3.0 1e-06 
3.0 2.634 0 3.0 1e-06 
0.05 2.635 0 3.0 1e-06 
3.0 2.635 0 3.0 1e-06 
0.05 2.636 0 3.0 1e-06 
3.0 2.636 0 3.0 1e-06 
0.05 2.637 0 3.0 1e-06 
3.0 2.637 0 3.0 1e-06 
0.05 2.638 0 3.0 1e-06 
3.0 2.638 0 3.0 1e-06 
0.05 2.639 0 3.0 1e-06 
3.0 2.639 0 3.0 1e-06 
0.05 2.64 0 3.0 1e-06 
3.0 2.64 0 3.0 1e-06 
0.05 2.641 0 3.0 1e-06 
3.0 2.641 0 3.0 1e-06 
0.05 2.642 0 3.0 1e-06 
3.0 2.642 0 3.0 1e-06 
0.05 2.643 0 3.0 1e-06 
3.0 2.643 0 3.0 1e-06 
0.05 2.644 0 3.0 1e-06 
3.0 2.644 0 3.0 1e-06 
0.05 2.645 0 3.0 1e-06 
3.0 2.645 0 3.0 1e-06 
0.05 2.646 0 3.0 1e-06 
3.0 2.646 0 3.0 1e-06 
0.05 2.647 0 3.0 1e-06 
3.0 2.647 0 3.0 1e-06 
0.05 2.648 0 3.0 1e-06 
3.0 2.648 0 3.0 1e-06 
0.05 2.649 0 3.0 1e-06 
3.0 2.649 0 3.0 1e-06 
0.05 2.65 0 3.0 1e-06 
3.0 2.65 0 3.0 1e-06 
0.05 2.651 0 3.0 1e-06 
3.0 2.651 0 3.0 1e-06 
0.05 2.652 0 3.0 1e-06 
3.0 2.652 0 3.0 1e-06 
0.05 2.653 0 3.0 1e-06 
3.0 2.653 0 3.0 1e-06 
0.05 2.654 0 3.0 1e-06 
3.0 2.654 0 3.0 1e-06 
0.05 2.655 0 3.0 1e-06 
3.0 2.655 0 3.0 1e-06 
0.05 2.656 0 3.0 1e-06 
3.0 2.656 0 3.0 1e-06 
0.05 2.657 0 3.0 1e-06 
3.0 2.657 0 3.0 1e-06 
0.05 2.658 0 3.0 1e-06 
3.0 2.658 0 3.0 1e-06 
0.05 2.659 0 3.0 1e-06 
3.0 2.659 0 3.0 1e-06 
0.05 2.66 0 3.0 1e-06 
3.0 2.66 0 3.0 1e-06 
0.05 2.661 0 3.0 1e-06 
3.0 2.661 0 3.0 1e-06 
0.05 2.662 0 3.0 1e-06 
3.0 2.662 0 3.0 1e-06 
0.05 2.663 0 3.0 1e-06 
3.0 2.663 0 3.0 1e-06 
0.05 2.664 0 3.0 1e-06 
3.0 2.664 0 3.0 1e-06 
0.05 2.665 0 3.0 1e-06 
3.0 2.665 0 3.0 1e-06 
0.05 2.666 0 3.0 1e-06 
3.0 2.666 0 3.0 1e-06 
0.05 2.667 0 3.0 1e-06 
3.0 2.667 0 3.0 1e-06 
0.05 2.668 0 3.0 1e-06 
3.0 2.668 0 3.0 1e-06 
0.05 2.669 0 3.0 1e-06 
3.0 2.669 0 3.0 1e-06 
0.05 2.67 0 3.0 1e-06 
3.0 2.67 0 3.0 1e-06 
0.05 2.671 0 3.0 1e-06 
3.0 2.671 0 3.0 1e-06 
0.05 2.672 0 3.0 1e-06 
3.0 2.672 0 3.0 1e-06 
0.05 2.673 0 3.0 1e-06 
3.0 2.673 0 3.0 1e-06 
0.05 2.674 0 3.0 1e-06 
3.0 2.674 0 3.0 1e-06 
0.05 2.675 0 3.0 1e-06 
3.0 2.675 0 3.0 1e-06 
0.05 2.676 0 3.0 1e-06 
3.0 2.676 0 3.0 1e-06 
0.05 2.677 0 3.0 1e-06 
3.0 2.677 0 3.0 1e-06 
0.05 2.678 0 3.0 1e-06 
3.0 2.678 0 3.0 1e-06 
0.05 2.679 0 3.0 1e-06 
3.0 2.679 0 3.0 1e-06 
0.05 2.68 0 3.0 1e-06 
3.0 2.68 0 3.0 1e-06 
0.05 2.681 0 3.0 1e-06 
3.0 2.681 0 3.0 1e-06 
0.05 2.682 0 3.0 1e-06 
3.0 2.682 0 3.0 1e-06 
0.05 2.683 0 3.0 1e-06 
3.0 2.683 0 3.0 1e-06 
0.05 2.684 0 3.0 1e-06 
3.0 2.684 0 3.0 1e-06 
0.05 2.685 0 3.0 1e-06 
3.0 2.685 0 3.0 1e-06 
0.05 2.686 0 3.0 1e-06 
3.0 2.686 0 3.0 1e-06 
0.05 2.687 0 3.0 1e-06 
3.0 2.687 0 3.0 1e-06 
0.05 2.688 0 3.0 1e-06 
3.0 2.688 0 3.0 1e-06 
0.05 2.689 0 3.0 1e-06 
3.0 2.689 0 3.0 1e-06 
0.05 2.69 0 3.0 1e-06 
3.0 2.69 0 3.0 1e-06 
0.05 2.691 0 3.0 1e-06 
3.0 2.691 0 3.0 1e-06 
0.05 2.692 0 3.0 1e-06 
3.0 2.692 0 3.0 1e-06 
0.05 2.693 0 3.0 1e-06 
3.0 2.693 0 3.0 1e-06 
0.05 2.694 0 3.0 1e-06 
3.0 2.694 0 3.0 1e-06 
0.05 2.695 0 3.0 1e-06 
3.0 2.695 0 3.0 1e-06 
0.05 2.696 0 3.0 1e-06 
3.0 2.696 0 3.0 1e-06 
0.05 2.697 0 3.0 1e-06 
3.0 2.697 0 3.0 1e-06 
0.05 2.698 0 3.0 1e-06 
3.0 2.698 0 3.0 1e-06 
0.05 2.699 0 3.0 1e-06 
3.0 2.699 0 3.0 1e-06 
0.05 2.7 0 3.0 1e-06 
3.0 2.7 0 3.0 1e-06 
0.05 2.701 0 3.0 1e-06 
3.0 2.701 0 3.0 1e-06 
0.05 2.702 0 3.0 1e-06 
3.0 2.702 0 3.0 1e-06 
0.05 2.703 0 3.0 1e-06 
3.0 2.703 0 3.0 1e-06 
0.05 2.704 0 3.0 1e-06 
3.0 2.704 0 3.0 1e-06 
0.05 2.705 0 3.0 1e-06 
3.0 2.705 0 3.0 1e-06 
0.05 2.706 0 3.0 1e-06 
3.0 2.706 0 3.0 1e-06 
0.05 2.707 0 3.0 1e-06 
3.0 2.707 0 3.0 1e-06 
0.05 2.708 0 3.0 1e-06 
3.0 2.708 0 3.0 1e-06 
0.05 2.709 0 3.0 1e-06 
3.0 2.709 0 3.0 1e-06 
0.05 2.71 0 3.0 1e-06 
3.0 2.71 0 3.0 1e-06 
0.05 2.711 0 3.0 1e-06 
3.0 2.711 0 3.0 1e-06 
0.05 2.712 0 3.0 1e-06 
3.0 2.712 0 3.0 1e-06 
0.05 2.713 0 3.0 1e-06 
3.0 2.713 0 3.0 1e-06 
0.05 2.714 0 3.0 1e-06 
3.0 2.714 0 3.0 1e-06 
0.05 2.715 0 3.0 1e-06 
3.0 2.715 0 3.0 1e-06 
0.05 2.716 0 3.0 1e-06 
3.0 2.716 0 3.0 1e-06 
0.05 2.717 0 3.0 1e-06 
3.0 2.717 0 3.0 1e-06 
0.05 2.718 0 3.0 1e-06 
3.0 2.718 0 3.0 1e-06 
0.05 2.719 0 3.0 1e-06 
3.0 2.719 0 3.0 1e-06 
0.05 2.72 0 3.0 1e-06 
3.0 2.72 0 3.0 1e-06 
0.05 2.721 0 3.0 1e-06 
3.0 2.721 0 3.0 1e-06 
0.05 2.722 0 3.0 1e-06 
3.0 2.722 0 3.0 1e-06 
0.05 2.723 0 3.0 1e-06 
3.0 2.723 0 3.0 1e-06 
0.05 2.724 0 3.0 1e-06 
3.0 2.724 0 3.0 1e-06 
0.05 2.725 0 3.0 1e-06 
3.0 2.725 0 3.0 1e-06 
0.05 2.726 0 3.0 1e-06 
3.0 2.726 0 3.0 1e-06 
0.05 2.727 0 3.0 1e-06 
3.0 2.727 0 3.0 1e-06 
0.05 2.728 0 3.0 1e-06 
3.0 2.728 0 3.0 1e-06 
0.05 2.729 0 3.0 1e-06 
3.0 2.729 0 3.0 1e-06 
0.05 2.73 0 3.0 1e-06 
3.0 2.73 0 3.0 1e-06 
0.05 2.731 0 3.0 1e-06 
3.0 2.731 0 3.0 1e-06 
0.05 2.732 0 3.0 1e-06 
3.0 2.732 0 3.0 1e-06 
0.05 2.733 0 3.0 1e-06 
3.0 2.733 0 3.0 1e-06 
0.05 2.734 0 3.0 1e-06 
3.0 2.734 0 3.0 1e-06 
0.05 2.735 0 3.0 1e-06 
3.0 2.735 0 3.0 1e-06 
0.05 2.736 0 3.0 1e-06 
3.0 2.736 0 3.0 1e-06 
0.05 2.737 0 3.0 1e-06 
3.0 2.737 0 3.0 1e-06 
0.05 2.738 0 3.0 1e-06 
3.0 2.738 0 3.0 1e-06 
0.05 2.739 0 3.0 1e-06 
3.0 2.739 0 3.0 1e-06 
0.05 2.74 0 3.0 1e-06 
3.0 2.74 0 3.0 1e-06 
0.05 2.741 0 3.0 1e-06 
3.0 2.741 0 3.0 1e-06 
0.05 2.742 0 3.0 1e-06 
3.0 2.742 0 3.0 1e-06 
0.05 2.743 0 3.0 1e-06 
3.0 2.743 0 3.0 1e-06 
0.05 2.744 0 3.0 1e-06 
3.0 2.744 0 3.0 1e-06 
0.05 2.745 0 3.0 1e-06 
3.0 2.745 0 3.0 1e-06 
0.05 2.746 0 3.0 1e-06 
3.0 2.746 0 3.0 1e-06 
0.05 2.747 0 3.0 1e-06 
3.0 2.747 0 3.0 1e-06 
0.05 2.748 0 3.0 1e-06 
3.0 2.748 0 3.0 1e-06 
0.05 2.749 0 3.0 1e-06 
3.0 2.749 0 3.0 1e-06 
0.05 2.75 0 3.0 1e-06 
3.0 2.75 0 3.0 1e-06 
0.05 2.751 0 3.0 1e-06 
3.0 2.751 0 3.0 1e-06 
0.05 2.752 0 3.0 1e-06 
3.0 2.752 0 3.0 1e-06 
0.05 2.753 0 3.0 1e-06 
3.0 2.753 0 3.0 1e-06 
0.05 2.754 0 3.0 1e-06 
3.0 2.754 0 3.0 1e-06 
0.05 2.755 0 3.0 1e-06 
3.0 2.755 0 3.0 1e-06 
0.05 2.756 0 3.0 1e-06 
3.0 2.756 0 3.0 1e-06 
0.05 2.757 0 3.0 1e-06 
3.0 2.757 0 3.0 1e-06 
0.05 2.758 0 3.0 1e-06 
3.0 2.758 0 3.0 1e-06 
0.05 2.759 0 3.0 1e-06 
3.0 2.759 0 3.0 1e-06 
0.05 2.76 0 3.0 1e-06 
3.0 2.76 0 3.0 1e-06 
0.05 2.761 0 3.0 1e-06 
3.0 2.761 0 3.0 1e-06 
0.05 2.762 0 3.0 1e-06 
3.0 2.762 0 3.0 1e-06 
0.05 2.763 0 3.0 1e-06 
3.0 2.763 0 3.0 1e-06 
0.05 2.764 0 3.0 1e-06 
3.0 2.764 0 3.0 1e-06 
0.05 2.765 0 3.0 1e-06 
3.0 2.765 0 3.0 1e-06 
0.05 2.766 0 3.0 1e-06 
3.0 2.766 0 3.0 1e-06 
0.05 2.767 0 3.0 1e-06 
3.0 2.767 0 3.0 1e-06 
0.05 2.768 0 3.0 1e-06 
3.0 2.768 0 3.0 1e-06 
0.05 2.769 0 3.0 1e-06 
3.0 2.769 0 3.0 1e-06 
0.05 2.77 0 3.0 1e-06 
3.0 2.77 0 3.0 1e-06 
0.05 2.771 0 3.0 1e-06 
3.0 2.771 0 3.0 1e-06 
0.05 2.772 0 3.0 1e-06 
3.0 2.772 0 3.0 1e-06 
0.05 2.773 0 3.0 1e-06 
3.0 2.773 0 3.0 1e-06 
0.05 2.774 0 3.0 1e-06 
3.0 2.774 0 3.0 1e-06 
0.05 2.775 0 3.0 1e-06 
3.0 2.775 0 3.0 1e-06 
0.05 2.776 0 3.0 1e-06 
3.0 2.776 0 3.0 1e-06 
0.05 2.777 0 3.0 1e-06 
3.0 2.777 0 3.0 1e-06 
0.05 2.778 0 3.0 1e-06 
3.0 2.778 0 3.0 1e-06 
0.05 2.779 0 3.0 1e-06 
3.0 2.779 0 3.0 1e-06 
0.05 2.78 0 3.0 1e-06 
3.0 2.78 0 3.0 1e-06 
0.05 2.781 0 3.0 1e-06 
3.0 2.781 0 3.0 1e-06 
0.05 2.782 0 3.0 1e-06 
3.0 2.782 0 3.0 1e-06 
0.05 2.783 0 3.0 1e-06 
3.0 2.783 0 3.0 1e-06 
0.05 2.784 0 3.0 1e-06 
3.0 2.784 0 3.0 1e-06 
0.05 2.785 0 3.0 1e-06 
3.0 2.785 0 3.0 1e-06 
0.05 2.786 0 3.0 1e-06 
3.0 2.786 0 3.0 1e-06 
0.05 2.787 0 3.0 1e-06 
3.0 2.787 0 3.0 1e-06 
0.05 2.788 0 3.0 1e-06 
3.0 2.788 0 3.0 1e-06 
0.05 2.789 0 3.0 1e-06 
3.0 2.789 0 3.0 1e-06 
0.05 2.79 0 3.0 1e-06 
3.0 2.79 0 3.0 1e-06 
0.05 2.791 0 3.0 1e-06 
3.0 2.791 0 3.0 1e-06 
0.05 2.792 0 3.0 1e-06 
3.0 2.792 0 3.0 1e-06 
0.05 2.793 0 3.0 1e-06 
3.0 2.793 0 3.0 1e-06 
0.05 2.794 0 3.0 1e-06 
3.0 2.794 0 3.0 1e-06 
0.05 2.795 0 3.0 1e-06 
3.0 2.795 0 3.0 1e-06 
0.05 2.796 0 3.0 1e-06 
3.0 2.796 0 3.0 1e-06 
0.05 2.797 0 3.0 1e-06 
3.0 2.797 0 3.0 1e-06 
0.05 2.798 0 3.0 1e-06 
3.0 2.798 0 3.0 1e-06 
0.05 2.799 0 3.0 1e-06 
3.0 2.799 0 3.0 1e-06 
0.05 2.8 0 3.0 1e-06 
3.0 2.8 0 3.0 1e-06 
0.05 2.801 0 3.0 1e-06 
3.0 2.801 0 3.0 1e-06 
0.05 2.802 0 3.0 1e-06 
3.0 2.802 0 3.0 1e-06 
0.05 2.803 0 3.0 1e-06 
3.0 2.803 0 3.0 1e-06 
0.05 2.804 0 3.0 1e-06 
3.0 2.804 0 3.0 1e-06 
0.05 2.805 0 3.0 1e-06 
3.0 2.805 0 3.0 1e-06 
0.05 2.806 0 3.0 1e-06 
3.0 2.806 0 3.0 1e-06 
0.05 2.807 0 3.0 1e-06 
3.0 2.807 0 3.0 1e-06 
0.05 2.808 0 3.0 1e-06 
3.0 2.808 0 3.0 1e-06 
0.05 2.809 0 3.0 1e-06 
3.0 2.809 0 3.0 1e-06 
0.05 2.81 0 3.0 1e-06 
3.0 2.81 0 3.0 1e-06 
0.05 2.811 0 3.0 1e-06 
3.0 2.811 0 3.0 1e-06 
0.05 2.812 0 3.0 1e-06 
3.0 2.812 0 3.0 1e-06 
0.05 2.813 0 3.0 1e-06 
3.0 2.813 0 3.0 1e-06 
0.05 2.814 0 3.0 1e-06 
3.0 2.814 0 3.0 1e-06 
0.05 2.815 0 3.0 1e-06 
3.0 2.815 0 3.0 1e-06 
0.05 2.816 0 3.0 1e-06 
3.0 2.816 0 3.0 1e-06 
0.05 2.817 0 3.0 1e-06 
3.0 2.817 0 3.0 1e-06 
0.05 2.818 0 3.0 1e-06 
3.0 2.818 0 3.0 1e-06 
0.05 2.819 0 3.0 1e-06 
3.0 2.819 0 3.0 1e-06 
0.05 2.82 0 3.0 1e-06 
3.0 2.82 0 3.0 1e-06 
0.05 2.821 0 3.0 1e-06 
3.0 2.821 0 3.0 1e-06 
0.05 2.822 0 3.0 1e-06 
3.0 2.822 0 3.0 1e-06 
0.05 2.823 0 3.0 1e-06 
3.0 2.823 0 3.0 1e-06 
0.05 2.824 0 3.0 1e-06 
3.0 2.824 0 3.0 1e-06 
0.05 2.825 0 3.0 1e-06 
3.0 2.825 0 3.0 1e-06 
0.05 2.826 0 3.0 1e-06 
3.0 2.826 0 3.0 1e-06 
0.05 2.827 0 3.0 1e-06 
3.0 2.827 0 3.0 1e-06 
0.05 2.828 0 3.0 1e-06 
3.0 2.828 0 3.0 1e-06 
0.05 2.829 0 3.0 1e-06 
3.0 2.829 0 3.0 1e-06 
0.05 2.83 0 3.0 1e-06 
3.0 2.83 0 3.0 1e-06 
0.05 2.831 0 3.0 1e-06 
3.0 2.831 0 3.0 1e-06 
0.05 2.832 0 3.0 1e-06 
3.0 2.832 0 3.0 1e-06 
0.05 2.833 0 3.0 1e-06 
3.0 2.833 0 3.0 1e-06 
0.05 2.834 0 3.0 1e-06 
3.0 2.834 0 3.0 1e-06 
0.05 2.835 0 3.0 1e-06 
3.0 2.835 0 3.0 1e-06 
0.05 2.836 0 3.0 1e-06 
3.0 2.836 0 3.0 1e-06 
0.05 2.837 0 3.0 1e-06 
3.0 2.837 0 3.0 1e-06 
0.05 2.838 0 3.0 1e-06 
3.0 2.838 0 3.0 1e-06 
0.05 2.839 0 3.0 1e-06 
3.0 2.839 0 3.0 1e-06 
0.05 2.84 0 3.0 1e-06 
3.0 2.84 0 3.0 1e-06 
0.05 2.841 0 3.0 1e-06 
3.0 2.841 0 3.0 1e-06 
0.05 2.842 0 3.0 1e-06 
3.0 2.842 0 3.0 1e-06 
0.05 2.843 0 3.0 1e-06 
3.0 2.843 0 3.0 1e-06 
0.05 2.844 0 3.0 1e-06 
3.0 2.844 0 3.0 1e-06 
0.05 2.845 0 3.0 1e-06 
3.0 2.845 0 3.0 1e-06 
0.05 2.846 0 3.0 1e-06 
3.0 2.846 0 3.0 1e-06 
0.05 2.847 0 3.0 1e-06 
3.0 2.847 0 3.0 1e-06 
0.05 2.848 0 3.0 1e-06 
3.0 2.848 0 3.0 1e-06 
0.05 2.849 0 3.0 1e-06 
3.0 2.849 0 3.0 1e-06 
0.05 2.85 0 3.0 1e-06 
3.0 2.85 0 3.0 1e-06 
0.05 2.851 0 3.0 1e-06 
3.0 2.851 0 3.0 1e-06 
0.05 2.852 0 3.0 1e-06 
3.0 2.852 0 3.0 1e-06 
0.05 2.853 0 3.0 1e-06 
3.0 2.853 0 3.0 1e-06 
0.05 2.854 0 3.0 1e-06 
3.0 2.854 0 3.0 1e-06 
0.05 2.855 0 3.0 1e-06 
3.0 2.855 0 3.0 1e-06 
0.05 2.856 0 3.0 1e-06 
3.0 2.856 0 3.0 1e-06 
0.05 2.857 0 3.0 1e-06 
3.0 2.857 0 3.0 1e-06 
0.05 2.858 0 3.0 1e-06 
3.0 2.858 0 3.0 1e-06 
0.05 2.859 0 3.0 1e-06 
3.0 2.859 0 3.0 1e-06 
0.05 2.86 0 3.0 1e-06 
3.0 2.86 0 3.0 1e-06 
0.05 2.861 0 3.0 1e-06 
3.0 2.861 0 3.0 1e-06 
0.05 2.862 0 3.0 1e-06 
3.0 2.862 0 3.0 1e-06 
0.05 2.863 0 3.0 1e-06 
3.0 2.863 0 3.0 1e-06 
0.05 2.864 0 3.0 1e-06 
3.0 2.864 0 3.0 1e-06 
0.05 2.865 0 3.0 1e-06 
3.0 2.865 0 3.0 1e-06 
0.05 2.866 0 3.0 1e-06 
3.0 2.866 0 3.0 1e-06 
0.05 2.867 0 3.0 1e-06 
3.0 2.867 0 3.0 1e-06 
0.05 2.868 0 3.0 1e-06 
3.0 2.868 0 3.0 1e-06 
0.05 2.869 0 3.0 1e-06 
3.0 2.869 0 3.0 1e-06 
0.05 2.87 0 3.0 1e-06 
3.0 2.87 0 3.0 1e-06 
0.05 2.871 0 3.0 1e-06 
3.0 2.871 0 3.0 1e-06 
0.05 2.872 0 3.0 1e-06 
3.0 2.872 0 3.0 1e-06 
0.05 2.873 0 3.0 1e-06 
3.0 2.873 0 3.0 1e-06 
0.05 2.874 0 3.0 1e-06 
3.0 2.874 0 3.0 1e-06 
0.05 2.875 0 3.0 1e-06 
3.0 2.875 0 3.0 1e-06 
0.05 2.876 0 3.0 1e-06 
3.0 2.876 0 3.0 1e-06 
0.05 2.877 0 3.0 1e-06 
3.0 2.877 0 3.0 1e-06 
0.05 2.878 0 3.0 1e-06 
3.0 2.878 0 3.0 1e-06 
0.05 2.879 0 3.0 1e-06 
3.0 2.879 0 3.0 1e-06 
0.05 2.88 0 3.0 1e-06 
3.0 2.88 0 3.0 1e-06 
0.05 2.881 0 3.0 1e-06 
3.0 2.881 0 3.0 1e-06 
0.05 2.882 0 3.0 1e-06 
3.0 2.882 0 3.0 1e-06 
0.05 2.883 0 3.0 1e-06 
3.0 2.883 0 3.0 1e-06 
0.05 2.884 0 3.0 1e-06 
3.0 2.884 0 3.0 1e-06 
0.05 2.885 0 3.0 1e-06 
3.0 2.885 0 3.0 1e-06 
0.05 2.886 0 3.0 1e-06 
3.0 2.886 0 3.0 1e-06 
0.05 2.887 0 3.0 1e-06 
3.0 2.887 0 3.0 1e-06 
0.05 2.888 0 3.0 1e-06 
3.0 2.888 0 3.0 1e-06 
0.05 2.889 0 3.0 1e-06 
3.0 2.889 0 3.0 1e-06 
0.05 2.89 0 3.0 1e-06 
3.0 2.89 0 3.0 1e-06 
0.05 2.891 0 3.0 1e-06 
3.0 2.891 0 3.0 1e-06 
0.05 2.892 0 3.0 1e-06 
3.0 2.892 0 3.0 1e-06 
0.05 2.893 0 3.0 1e-06 
3.0 2.893 0 3.0 1e-06 
0.05 2.894 0 3.0 1e-06 
3.0 2.894 0 3.0 1e-06 
0.05 2.895 0 3.0 1e-06 
3.0 2.895 0 3.0 1e-06 
0.05 2.896 0 3.0 1e-06 
3.0 2.896 0 3.0 1e-06 
0.05 2.897 0 3.0 1e-06 
3.0 2.897 0 3.0 1e-06 
0.05 2.898 0 3.0 1e-06 
3.0 2.898 0 3.0 1e-06 
0.05 2.899 0 3.0 1e-06 
3.0 2.899 0 3.0 1e-06 
0.05 2.9 0 3.0 1e-06 
3.0 2.9 0 3.0 1e-06 
0.05 2.901 0 3.0 1e-06 
3.0 2.901 0 3.0 1e-06 
0.05 2.902 0 3.0 1e-06 
3.0 2.902 0 3.0 1e-06 
0.05 2.903 0 3.0 1e-06 
3.0 2.903 0 3.0 1e-06 
0.05 2.904 0 3.0 1e-06 
3.0 2.904 0 3.0 1e-06 
0.05 2.905 0 3.0 1e-06 
3.0 2.905 0 3.0 1e-06 
0.05 2.906 0 3.0 1e-06 
3.0 2.906 0 3.0 1e-06 
0.05 2.907 0 3.0 1e-06 
3.0 2.907 0 3.0 1e-06 
0.05 2.908 0 3.0 1e-06 
3.0 2.908 0 3.0 1e-06 
0.05 2.909 0 3.0 1e-06 
3.0 2.909 0 3.0 1e-06 
0.05 2.91 0 3.0 1e-06 
3.0 2.91 0 3.0 1e-06 
0.05 2.911 0 3.0 1e-06 
3.0 2.911 0 3.0 1e-06 
0.05 2.912 0 3.0 1e-06 
3.0 2.912 0 3.0 1e-06 
0.05 2.913 0 3.0 1e-06 
3.0 2.913 0 3.0 1e-06 
0.05 2.914 0 3.0 1e-06 
3.0 2.914 0 3.0 1e-06 
0.05 2.915 0 3.0 1e-06 
3.0 2.915 0 3.0 1e-06 
0.05 2.916 0 3.0 1e-06 
3.0 2.916 0 3.0 1e-06 
0.05 2.917 0 3.0 1e-06 
3.0 2.917 0 3.0 1e-06 
0.05 2.918 0 3.0 1e-06 
3.0 2.918 0 3.0 1e-06 
0.05 2.919 0 3.0 1e-06 
3.0 2.919 0 3.0 1e-06 
0.05 2.92 0 3.0 1e-06 
3.0 2.92 0 3.0 1e-06 
0.05 2.921 0 3.0 1e-06 
3.0 2.921 0 3.0 1e-06 
0.05 2.922 0 3.0 1e-06 
3.0 2.922 0 3.0 1e-06 
0.05 2.923 0 3.0 1e-06 
3.0 2.923 0 3.0 1e-06 
0.05 2.924 0 3.0 1e-06 
3.0 2.924 0 3.0 1e-06 
0.05 2.925 0 3.0 1e-06 
3.0 2.925 0 3.0 1e-06 
0.05 2.926 0 3.0 1e-06 
3.0 2.926 0 3.0 1e-06 
0.05 2.927 0 3.0 1e-06 
3.0 2.927 0 3.0 1e-06 
0.05 2.928 0 3.0 1e-06 
3.0 2.928 0 3.0 1e-06 
0.05 2.929 0 3.0 1e-06 
3.0 2.929 0 3.0 1e-06 
0.05 2.93 0 3.0 1e-06 
3.0 2.93 0 3.0 1e-06 
0.05 2.931 0 3.0 1e-06 
3.0 2.931 0 3.0 1e-06 
0.05 2.932 0 3.0 1e-06 
3.0 2.932 0 3.0 1e-06 
0.05 2.933 0 3.0 1e-06 
3.0 2.933 0 3.0 1e-06 
0.05 2.934 0 3.0 1e-06 
3.0 2.934 0 3.0 1e-06 
0.05 2.935 0 3.0 1e-06 
3.0 2.935 0 3.0 1e-06 
0.05 2.936 0 3.0 1e-06 
3.0 2.936 0 3.0 1e-06 
0.05 2.937 0 3.0 1e-06 
3.0 2.937 0 3.0 1e-06 
0.05 2.938 0 3.0 1e-06 
3.0 2.938 0 3.0 1e-06 
0.05 2.939 0 3.0 1e-06 
3.0 2.939 0 3.0 1e-06 
0.05 2.94 0 3.0 1e-06 
3.0 2.94 0 3.0 1e-06 
0.05 2.941 0 3.0 1e-06 
3.0 2.941 0 3.0 1e-06 
0.05 2.942 0 3.0 1e-06 
3.0 2.942 0 3.0 1e-06 
0.05 2.943 0 3.0 1e-06 
3.0 2.943 0 3.0 1e-06 
0.05 2.944 0 3.0 1e-06 
3.0 2.944 0 3.0 1e-06 
0.05 2.945 0 3.0 1e-06 
3.0 2.945 0 3.0 1e-06 
0.05 2.946 0 3.0 1e-06 
3.0 2.946 0 3.0 1e-06 
0.05 2.947 0 3.0 1e-06 
3.0 2.947 0 3.0 1e-06 
0.05 2.948 0 3.0 1e-06 
3.0 2.948 0 3.0 1e-06 
0.05 2.949 0 3.0 1e-06 
3.0 2.949 0 3.0 1e-06 
0.05 2.95 0 3.0 1e-06 
3.0 2.95 0 3.0 1e-06 
0.05 2.951 0 3.0 1e-06 
3.0 2.951 0 3.0 1e-06 
0.05 2.952 0 3.0 1e-06 
3.0 2.952 0 3.0 1e-06 
0.05 2.953 0 3.0 1e-06 
3.0 2.953 0 3.0 1e-06 
0.05 2.954 0 3.0 1e-06 
3.0 2.954 0 3.0 1e-06 
0.05 2.955 0 3.0 1e-06 
3.0 2.955 0 3.0 1e-06 
0.05 2.956 0 3.0 1e-06 
3.0 2.956 0 3.0 1e-06 
0.05 2.957 0 3.0 1e-06 
3.0 2.957 0 3.0 1e-06 
0.05 2.958 0 3.0 1e-06 
3.0 2.958 0 3.0 1e-06 
0.05 2.959 0 3.0 1e-06 
3.0 2.959 0 3.0 1e-06 
0.05 2.96 0 3.0 1e-06 
3.0 2.96 0 3.0 1e-06 
0.05 2.961 0 3.0 1e-06 
3.0 2.961 0 3.0 1e-06 
0.05 2.962 0 3.0 1e-06 
3.0 2.962 0 3.0 1e-06 
0.05 2.963 0 3.0 1e-06 
3.0 2.963 0 3.0 1e-06 
0.05 2.964 0 3.0 1e-06 
3.0 2.964 0 3.0 1e-06 
0.05 2.965 0 3.0 1e-06 
3.0 2.965 0 3.0 1e-06 
0.05 2.966 0 3.0 1e-06 
3.0 2.966 0 3.0 1e-06 
0.05 2.967 0 3.0 1e-06 
3.0 2.967 0 3.0 1e-06 
0.05 2.968 0 3.0 1e-06 
3.0 2.968 0 3.0 1e-06 
0.05 2.969 0 3.0 1e-06 
3.0 2.969 0 3.0 1e-06 
0.05 2.97 0 3.0 1e-06 
3.0 2.97 0 3.0 1e-06 
0.05 2.971 0 3.0 1e-06 
3.0 2.971 0 3.0 1e-06 
0.05 2.972 0 3.0 1e-06 
3.0 2.972 0 3.0 1e-06 
0.05 2.973 0 3.0 1e-06 
3.0 2.973 0 3.0 1e-06 
0.05 2.974 0 3.0 1e-06 
3.0 2.974 0 3.0 1e-06 
0.05 2.975 0 3.0 1e-06 
3.0 2.975 0 3.0 1e-06 
0.05 2.976 0 3.0 1e-06 
3.0 2.976 0 3.0 1e-06 
0.05 2.977 0 3.0 1e-06 
3.0 2.977 0 3.0 1e-06 
0.05 2.978 0 3.0 1e-06 
3.0 2.978 0 3.0 1e-06 
0.05 2.979 0 3.0 1e-06 
3.0 2.979 0 3.0 1e-06 
0.05 2.98 0 3.0 1e-06 
3.0 2.98 0 3.0 1e-06 
0.05 2.981 0 3.0 1e-06 
3.0 2.981 0 3.0 1e-06 
0.05 2.982 0 3.0 1e-06 
3.0 2.982 0 3.0 1e-06 
0.05 2.983 0 3.0 1e-06 
3.0 2.983 0 3.0 1e-06 
0.05 2.984 0 3.0 1e-06 
3.0 2.984 0 3.0 1e-06 
0.05 2.985 0 3.0 1e-06 
3.0 2.985 0 3.0 1e-06 
0.05 2.986 0 3.0 1e-06 
3.0 2.986 0 3.0 1e-06 
0.05 2.987 0 3.0 1e-06 
3.0 2.987 0 3.0 1e-06 
0.05 2.988 0 3.0 1e-06 
3.0 2.988 0 3.0 1e-06 
0.05 2.989 0 3.0 1e-06 
3.0 2.989 0 3.0 1e-06 
0.05 2.99 0 3.0 1e-06 
3.0 2.99 0 3.0 1e-06 
0.05 2.991 0 3.0 1e-06 
3.0 2.991 0 3.0 1e-06 
0.05 2.992 0 3.0 1e-06 
3.0 2.992 0 3.0 1e-06 
0.05 2.993 0 3.0 1e-06 
3.0 2.993 0 3.0 1e-06 
0.05 2.994 0 3.0 1e-06 
3.0 2.994 0 3.0 1e-06 
0.05 2.995 0 3.0 1e-06 
3.0 2.995 0 3.0 1e-06 
0.05 2.996 0 3.0 1e-06 
3.0 2.996 0 3.0 1e-06 
0.05 2.997 0 3.0 1e-06 
3.0 2.997 0 3.0 1e-06 
0.05 2.998 0 3.0 1e-06 
3.0 2.998 0 3.0 1e-06 
0.05 2.999 0 3.0 1e-06 
3.0 2.999 0 3.0 1e-06 
0.05 3.0 0 3.0 1e-06 
3.0 3.0 0 3.0 1e-06 
0.05 3.001 0 3.0 1e-06 
3.0 3.001 0 3.0 1e-06 
0.05 3.002 0 3.0 1e-06 
3.0 3.002 0 3.0 1e-06 
0.05 3.003 0 3.0 1e-06 
3.0 3.003 0 3.0 1e-06 
0.05 3.004 0 3.0 1e-06 
3.0 3.004 0 3.0 1e-06 
0.05 3.005 0 3.0 1e-06 
3.0 3.005 0 3.0 1e-06 
0.05 3.006 0 3.0 1e-06 
3.0 3.006 0 3.0 1e-06 
0.05 3.007 0 3.0 1e-06 
3.0 3.007 0 3.0 1e-06 
0.05 3.008 0 3.0 1e-06 
3.0 3.008 0 3.0 1e-06 
0.05 3.009 0 3.0 1e-06 
3.0 3.009 0 3.0 1e-06 
0.05 3.01 0 3.0 1e-06 
3.0 3.01 0 3.0 1e-06 
0.05 3.011 0 3.0 1e-06 
3.0 3.011 0 3.0 1e-06 
0.05 3.012 0 3.0 1e-06 
3.0 3.012 0 3.0 1e-06 
0.05 3.013 0 3.0 1e-06 
3.0 3.013 0 3.0 1e-06 
0.05 3.014 0 3.0 1e-06 
3.0 3.014 0 3.0 1e-06 
0.05 3.015 0 3.0 1e-06 
3.0 3.015 0 3.0 1e-06 
0.05 3.016 0 3.0 1e-06 
3.0 3.016 0 3.0 1e-06 
0.05 3.017 0 3.0 1e-06 
3.0 3.017 0 3.0 1e-06 
0.05 3.018 0 3.0 1e-06 
3.0 3.018 0 3.0 1e-06 
0.05 3.019 0 3.0 1e-06 
3.0 3.019 0 3.0 1e-06 
0.05 3.02 0 3.0 1e-06 
3.0 3.02 0 3.0 1e-06 
0.05 3.021 0 3.0 1e-06 
3.0 3.021 0 3.0 1e-06 
0.05 3.022 0 3.0 1e-06 
3.0 3.022 0 3.0 1e-06 
0.05 3.023 0 3.0 1e-06 
3.0 3.023 0 3.0 1e-06 
0.05 3.024 0 3.0 1e-06 
3.0 3.024 0 3.0 1e-06 
0.05 3.025 0 3.0 1e-06 
3.0 3.025 0 3.0 1e-06 
0.05 3.026 0 3.0 1e-06 
3.0 3.026 0 3.0 1e-06 
0.05 3.027 0 3.0 1e-06 
3.0 3.027 0 3.0 1e-06 
0.05 3.028 0 3.0 1e-06 
3.0 3.028 0 3.0 1e-06 
0.05 3.029 0 3.0 1e-06 
3.0 3.029 0 3.0 1e-06 
0.05 3.03 0 3.0 1e-06 
3.0 3.03 0 3.0 1e-06 
0.05 3.031 0 3.0 1e-06 
3.0 3.031 0 3.0 1e-06 
0.05 3.032 0 3.0 1e-06 
3.0 3.032 0 3.0 1e-06 
0.05 3.033 0 3.0 1e-06 
3.0 3.033 0 3.0 1e-06 
0.05 3.034 0 3.0 1e-06 
3.0 3.034 0 3.0 1e-06 
0.05 3.035 0 3.0 1e-06 
3.0 3.035 0 3.0 1e-06 
0.05 3.036 0 3.0 1e-06 
3.0 3.036 0 3.0 1e-06 
0.05 3.037 0 3.0 1e-06 
3.0 3.037 0 3.0 1e-06 
0.05 3.038 0 3.0 1e-06 
3.0 3.038 0 3.0 1e-06 
0.05 3.039 0 3.0 1e-06 
3.0 3.039 0 3.0 1e-06 
0.05 3.04 0 3.0 1e-06 
3.0 3.04 0 3.0 1e-06 
0.05 3.041 0 3.0 1e-06 
3.0 3.041 0 3.0 1e-06 
0.05 3.042 0 3.0 1e-06 
3.0 3.042 0 3.0 1e-06 
0.05 3.043 0 3.0 1e-06 
3.0 3.043 0 3.0 1e-06 
0.05 3.044 0 3.0 1e-06 
3.0 3.044 0 3.0 1e-06 
0.05 3.045 0 3.0 1e-06 
3.0 3.045 0 3.0 1e-06 
0.05 3.046 0 3.0 1e-06 
3.0 3.046 0 3.0 1e-06 
0.05 3.047 0 3.0 1e-06 
3.0 3.047 0 3.0 1e-06 
0.05 3.048 0 3.0 1e-06 
3.0 3.048 0 3.0 1e-06 
0.05 3.049 0 3.0 1e-06 
3.0 3.049 0 3.0 1e-06 
0.05 3.05 0 3.0 1e-06 
3.0 3.05 0 3.0 1e-06 
0.05 3.051 0 3.0 1e-06 
3.0 3.051 0 3.0 1e-06 
0.05 3.052 0 3.0 1e-06 
3.0 3.052 0 3.0 1e-06 
0.05 3.053 0 3.0 1e-06 
3.0 3.053 0 3.0 1e-06 
0.05 3.054 0 3.0 1e-06 
3.0 3.054 0 3.0 1e-06 
0.05 3.055 0 3.0 1e-06 
3.0 3.055 0 3.0 1e-06 
0.05 3.056 0 3.0 1e-06 
3.0 3.056 0 3.0 1e-06 
0.05 3.057 0 3.0 1e-06 
3.0 3.057 0 3.0 1e-06 
0.05 3.058 0 3.0 1e-06 
3.0 3.058 0 3.0 1e-06 
0.05 3.059 0 3.0 1e-06 
3.0 3.059 0 3.0 1e-06 
0.05 3.06 0 3.0 1e-06 
3.0 3.06 0 3.0 1e-06 
0.05 3.061 0 3.0 1e-06 
3.0 3.061 0 3.0 1e-06 
0.05 3.062 0 3.0 1e-06 
3.0 3.062 0 3.0 1e-06 
0.05 3.063 0 3.0 1e-06 
3.0 3.063 0 3.0 1e-06 
0.05 3.064 0 3.0 1e-06 
3.0 3.064 0 3.0 1e-06 
0.05 3.065 0 3.0 1e-06 
3.0 3.065 0 3.0 1e-06 
0.05 3.066 0 3.0 1e-06 
3.0 3.066 0 3.0 1e-06 
0.05 3.067 0 3.0 1e-06 
3.0 3.067 0 3.0 1e-06 
0.05 3.068 0 3.0 1e-06 
3.0 3.068 0 3.0 1e-06 
0.05 3.069 0 3.0 1e-06 
3.0 3.069 0 3.0 1e-06 
0.05 3.07 0 3.0 1e-06 
3.0 3.07 0 3.0 1e-06 
0.05 3.071 0 3.0 1e-06 
3.0 3.071 0 3.0 1e-06 
0.05 3.072 0 3.0 1e-06 
3.0 3.072 0 3.0 1e-06 
0.05 3.073 0 3.0 1e-06 
3.0 3.073 0 3.0 1e-06 
0.05 3.074 0 3.0 1e-06 
3.0 3.074 0 3.0 1e-06 
0.05 3.075 0 3.0 1e-06 
3.0 3.075 0 3.0 1e-06 
0.05 3.076 0 3.0 1e-06 
3.0 3.076 0 3.0 1e-06 
0.05 3.077 0 3.0 1e-06 
3.0 3.077 0 3.0 1e-06 
0.05 3.078 0 3.0 1e-06 
3.0 3.078 0 3.0 1e-06 
0.05 3.079 0 3.0 1e-06 
3.0 3.079 0 3.0 1e-06 
0.05 3.08 0 3.0 1e-06 
3.0 3.08 0 3.0 1e-06 
0.05 3.081 0 3.0 1e-06 
3.0 3.081 0 3.0 1e-06 
0.05 3.082 0 3.0 1e-06 
3.0 3.082 0 3.0 1e-06 
0.05 3.083 0 3.0 1e-06 
3.0 3.083 0 3.0 1e-06 
0.05 3.084 0 3.0 1e-06 
3.0 3.084 0 3.0 1e-06 
0.05 3.085 0 3.0 1e-06 
3.0 3.085 0 3.0 1e-06 
0.05 3.086 0 3.0 1e-06 
3.0 3.086 0 3.0 1e-06 
0.05 3.087 0 3.0 1e-06 
3.0 3.087 0 3.0 1e-06 
0.05 3.088 0 3.0 1e-06 
3.0 3.088 0 3.0 1e-06 
0.05 3.089 0 3.0 1e-06 
3.0 3.089 0 3.0 1e-06 
0.05 3.09 0 3.0 1e-06 
3.0 3.09 0 3.0 1e-06 
0.05 3.091 0 3.0 1e-06 
3.0 3.091 0 3.0 1e-06 
0.05 3.092 0 3.0 1e-06 
3.0 3.092 0 3.0 1e-06 
0.05 3.093 0 3.0 1e-06 
3.0 3.093 0 3.0 1e-06 
0.05 3.094 0 3.0 1e-06 
3.0 3.094 0 3.0 1e-06 
0.05 3.095 0 3.0 1e-06 
3.0 3.095 0 3.0 1e-06 
0.05 3.096 0 3.0 1e-06 
3.0 3.096 0 3.0 1e-06 
0.05 3.097 0 3.0 1e-06 
3.0 3.097 0 3.0 1e-06 
0.05 3.098 0 3.0 1e-06 
3.0 3.098 0 3.0 1e-06 
0.05 3.099 0 3.0 1e-06 
3.0 3.099 0 3.0 1e-06 
0.05 3.1 0 3.0 1e-06 
3.0 3.1 0 3.0 1e-06 
0.05 3.101 0 3.0 1e-06 
3.0 3.101 0 3.0 1e-06 
0.05 3.102 0 3.0 1e-06 
3.0 3.102 0 3.0 1e-06 
0.05 3.103 0 3.0 1e-06 
3.0 3.103 0 3.0 1e-06 
0.05 3.104 0 3.0 1e-06 
3.0 3.104 0 3.0 1e-06 
0.05 3.105 0 3.0 1e-06 
3.0 3.105 0 3.0 1e-06 
0.05 3.106 0 3.0 1e-06 
3.0 3.106 0 3.0 1e-06 
0.05 3.107 0 3.0 1e-06 
3.0 3.107 0 3.0 1e-06 
0.05 3.108 0 3.0 1e-06 
3.0 3.108 0 3.0 1e-06 
0.05 3.109 0 3.0 1e-06 
3.0 3.109 0 3.0 1e-06 
0.05 3.11 0 3.0 1e-06 
3.0 3.11 0 3.0 1e-06 
0.05 3.111 0 3.0 1e-06 
3.0 3.111 0 3.0 1e-06 
0.05 3.112 0 3.0 1e-06 
3.0 3.112 0 3.0 1e-06 
0.05 3.113 0 3.0 1e-06 
3.0 3.113 0 3.0 1e-06 
0.05 3.114 0 3.0 1e-06 
3.0 3.114 0 3.0 1e-06 
0.05 3.115 0 3.0 1e-06 
3.0 3.115 0 3.0 1e-06 
0.05 3.116 0 3.0 1e-06 
3.0 3.116 0 3.0 1e-06 
0.05 3.117 0 3.0 1e-06 
3.0 3.117 0 3.0 1e-06 
0.05 3.118 0 3.0 1e-06 
3.0 3.118 0 3.0 1e-06 
0.05 3.119 0 3.0 1e-06 
3.0 3.119 0 3.0 1e-06 
0.05 3.12 0 3.0 1e-06 
3.0 3.12 0 3.0 1e-06 
0.05 3.121 0 3.0 1e-06 
3.0 3.121 0 3.0 1e-06 
0.05 3.122 0 3.0 1e-06 
3.0 3.122 0 3.0 1e-06 
0.05 3.123 0 3.0 1e-06 
3.0 3.123 0 3.0 1e-06 
0.05 3.124 0 3.0 1e-06 
3.0 3.124 0 3.0 1e-06 
0.05 3.125 0 3.0 1e-06 
3.0 3.125 0 3.0 1e-06 
0.05 3.126 0 3.0 1e-06 
3.0 3.126 0 3.0 1e-06 
0.05 3.127 0 3.0 1e-06 
3.0 3.127 0 3.0 1e-06 
0.05 3.128 0 3.0 1e-06 
3.0 3.128 0 3.0 1e-06 
0.05 3.129 0 3.0 1e-06 
3.0 3.129 0 3.0 1e-06 
0.05 3.13 0 3.0 1e-06 
3.0 3.13 0 3.0 1e-06 
0.05 3.131 0 3.0 1e-06 
3.0 3.131 0 3.0 1e-06 
0.05 3.132 0 3.0 1e-06 
3.0 3.132 0 3.0 1e-06 
0.05 3.133 0 3.0 1e-06 
3.0 3.133 0 3.0 1e-06 
0.05 3.134 0 3.0 1e-06 
3.0 3.134 0 3.0 1e-06 
0.05 3.135 0 3.0 1e-06 
3.0 3.135 0 3.0 1e-06 
0.05 3.136 0 3.0 1e-06 
3.0 3.136 0 3.0 1e-06 
0.05 3.137 0 3.0 1e-06 
3.0 3.137 0 3.0 1e-06 
0.05 3.138 0 3.0 1e-06 
3.0 3.138 0 3.0 1e-06 
0.05 3.139 0 3.0 1e-06 
3.0 3.139 0 3.0 1e-06 
0.05 3.14 0 3.0 1e-06 
3.0 3.14 0 3.0 1e-06 
0.05 3.141 0 3.0 1e-06 
3.0 3.141 0 3.0 1e-06 
0.05 3.142 0 3.0 1e-06 
3.0 3.142 0 3.0 1e-06 
0.05 3.143 0 3.0 1e-06 
3.0 3.143 0 3.0 1e-06 
0.05 3.144 0 3.0 1e-06 
3.0 3.144 0 3.0 1e-06 
0.05 3.145 0 3.0 1e-06 
3.0 3.145 0 3.0 1e-06 
0.05 3.146 0 3.0 1e-06 
3.0 3.146 0 3.0 1e-06 
0.05 3.147 0 3.0 1e-06 
3.0 3.147 0 3.0 1e-06 
0.05 3.148 0 3.0 1e-06 
3.0 3.148 0 3.0 1e-06 
0.05 3.149 0 3.0 1e-06 
3.0 3.149 0 3.0 1e-06 
0.05 3.15 0 3.0 1e-06 
3.0 3.15 0 3.0 1e-06 
0.05 3.151 0 3.0 1e-06 
3.0 3.151 0 3.0 1e-06 
0.05 3.152 0 3.0 1e-06 
3.0 3.152 0 3.0 1e-06 
0.05 3.153 0 3.0 1e-06 
3.0 3.153 0 3.0 1e-06 
0.05 3.154 0 3.0 1e-06 
3.0 3.154 0 3.0 1e-06 
0.05 3.155 0 3.0 1e-06 
3.0 3.155 0 3.0 1e-06 
0.05 3.156 0 3.0 1e-06 
3.0 3.156 0 3.0 1e-06 
0.05 3.157 0 3.0 1e-06 
3.0 3.157 0 3.0 1e-06 
0.05 3.158 0 3.0 1e-06 
3.0 3.158 0 3.0 1e-06 
0.05 3.159 0 3.0 1e-06 
3.0 3.159 0 3.0 1e-06 
0.05 3.16 0 3.0 1e-06 
3.0 3.16 0 3.0 1e-06 
0.05 3.161 0 3.0 1e-06 
3.0 3.161 0 3.0 1e-06 
0.05 3.162 0 3.0 1e-06 
3.0 3.162 0 3.0 1e-06 
0.05 3.163 0 3.0 1e-06 
3.0 3.163 0 3.0 1e-06 
0.05 3.164 0 3.0 1e-06 
3.0 3.164 0 3.0 1e-06 
0.05 3.165 0 3.0 1e-06 
3.0 3.165 0 3.0 1e-06 
0.05 3.166 0 3.0 1e-06 
3.0 3.166 0 3.0 1e-06 
0.05 3.167 0 3.0 1e-06 
3.0 3.167 0 3.0 1e-06 
0.05 3.168 0 3.0 1e-06 
3.0 3.168 0 3.0 1e-06 
0.05 3.169 0 3.0 1e-06 
3.0 3.169 0 3.0 1e-06 
0.05 3.17 0 3.0 1e-06 
3.0 3.17 0 3.0 1e-06 
0.05 3.171 0 3.0 1e-06 
3.0 3.171 0 3.0 1e-06 
0.05 3.172 0 3.0 1e-06 
3.0 3.172 0 3.0 1e-06 
0.05 3.173 0 3.0 1e-06 
3.0 3.173 0 3.0 1e-06 
0.05 3.174 0 3.0 1e-06 
3.0 3.174 0 3.0 1e-06 
0.05 3.175 0 3.0 1e-06 
3.0 3.175 0 3.0 1e-06 
0.05 3.176 0 3.0 1e-06 
3.0 3.176 0 3.0 1e-06 
0.05 3.177 0 3.0 1e-06 
3.0 3.177 0 3.0 1e-06 
0.05 3.178 0 3.0 1e-06 
3.0 3.178 0 3.0 1e-06 
0.05 3.179 0 3.0 1e-06 
3.0 3.179 0 3.0 1e-06 
0.05 3.18 0 3.0 1e-06 
3.0 3.18 0 3.0 1e-06 
0.05 3.181 0 3.0 1e-06 
3.0 3.181 0 3.0 1e-06 
0.05 3.182 0 3.0 1e-06 
3.0 3.182 0 3.0 1e-06 
0.05 3.183 0 3.0 1e-06 
3.0 3.183 0 3.0 1e-06 
0.05 3.184 0 3.0 1e-06 
3.0 3.184 0 3.0 1e-06 
0.05 3.185 0 3.0 1e-06 
3.0 3.185 0 3.0 1e-06 
0.05 3.186 0 3.0 1e-06 
3.0 3.186 0 3.0 1e-06 
0.05 3.187 0 3.0 1e-06 
3.0 3.187 0 3.0 1e-06 
0.05 3.188 0 3.0 1e-06 
3.0 3.188 0 3.0 1e-06 
0.05 3.189 0 3.0 1e-06 
3.0 3.189 0 3.0 1e-06 
0.05 3.19 0 3.0 1e-06 
3.0 3.19 0 3.0 1e-06 
0.05 3.191 0 3.0 1e-06 
3.0 3.191 0 3.0 1e-06 
0.05 3.192 0 3.0 1e-06 
3.0 3.192 0 3.0 1e-06 
0.05 3.193 0 3.0 1e-06 
3.0 3.193 0 3.0 1e-06 
0.05 3.194 0 3.0 1e-06 
3.0 3.194 0 3.0 1e-06 
0.05 3.195 0 3.0 1e-06 
3.0 3.195 0 3.0 1e-06 
0.05 3.196 0 3.0 1e-06 
3.0 3.196 0 3.0 1e-06 
0.05 3.197 0 3.0 1e-06 
3.0 3.197 0 3.0 1e-06 
0.05 3.198 0 3.0 1e-06 
3.0 3.198 0 3.0 1e-06 
0.05 3.199 0 3.0 1e-06 
3.0 3.199 0 3.0 1e-06 
0.05 3.2 0 3.0 1e-06 
3.0 3.2 0 3.0 1e-06 
0.05 3.201 0 3.0 1e-06 
3.0 3.201 0 3.0 1e-06 
0.05 3.202 0 3.0 1e-06 
3.0 3.202 0 3.0 1e-06 
0.05 3.203 0 3.0 1e-06 
3.0 3.203 0 3.0 1e-06 
0.05 3.204 0 3.0 1e-06 
3.0 3.204 0 3.0 1e-06 
0.05 3.205 0 3.0 1e-06 
3.0 3.205 0 3.0 1e-06 
0.05 3.206 0 3.0 1e-06 
3.0 3.206 0 3.0 1e-06 
0.05 3.207 0 3.0 1e-06 
3.0 3.207 0 3.0 1e-06 
0.05 3.208 0 3.0 1e-06 
3.0 3.208 0 3.0 1e-06 
0.05 3.209 0 3.0 1e-06 
3.0 3.209 0 3.0 1e-06 
0.05 3.21 0 3.0 1e-06 
3.0 3.21 0 3.0 1e-06 
0.05 3.211 0 3.0 1e-06 
3.0 3.211 0 3.0 1e-06 
0.05 3.212 0 3.0 1e-06 
3.0 3.212 0 3.0 1e-06 
0.05 3.213 0 3.0 1e-06 
3.0 3.213 0 3.0 1e-06 
0.05 3.214 0 3.0 1e-06 
3.0 3.214 0 3.0 1e-06 
0.05 3.215 0 3.0 1e-06 
3.0 3.215 0 3.0 1e-06 
0.05 3.216 0 3.0 1e-06 
3.0 3.216 0 3.0 1e-06 
0.05 3.217 0 3.0 1e-06 
3.0 3.217 0 3.0 1e-06 
0.05 3.218 0 3.0 1e-06 
3.0 3.218 0 3.0 1e-06 
0.05 3.219 0 3.0 1e-06 
3.0 3.219 0 3.0 1e-06 
0.05 3.22 0 3.0 1e-06 
3.0 3.22 0 3.0 1e-06 
0.05 3.221 0 3.0 1e-06 
3.0 3.221 0 3.0 1e-06 
0.05 3.222 0 3.0 1e-06 
3.0 3.222 0 3.0 1e-06 
0.05 3.223 0 3.0 1e-06 
3.0 3.223 0 3.0 1e-06 
0.05 3.224 0 3.0 1e-06 
3.0 3.224 0 3.0 1e-06 
0.05 3.225 0 3.0 1e-06 
3.0 3.225 0 3.0 1e-06 
0.05 3.226 0 3.0 1e-06 
3.0 3.226 0 3.0 1e-06 
0.05 3.227 0 3.0 1e-06 
3.0 3.227 0 3.0 1e-06 
0.05 3.228 0 3.0 1e-06 
3.0 3.228 0 3.0 1e-06 
0.05 3.229 0 3.0 1e-06 
3.0 3.229 0 3.0 1e-06 
0.05 3.23 0 3.0 1e-06 
3.0 3.23 0 3.0 1e-06 
0.05 3.231 0 3.0 1e-06 
3.0 3.231 0 3.0 1e-06 
0.05 3.232 0 3.0 1e-06 
3.0 3.232 0 3.0 1e-06 
0.05 3.233 0 3.0 1e-06 
3.0 3.233 0 3.0 1e-06 
0.05 3.234 0 3.0 1e-06 
3.0 3.234 0 3.0 1e-06 
0.05 3.235 0 3.0 1e-06 
3.0 3.235 0 3.0 1e-06 
0.05 3.236 0 3.0 1e-06 
3.0 3.236 0 3.0 1e-06 
0.05 3.237 0 3.0 1e-06 
3.0 3.237 0 3.0 1e-06 
0.05 3.238 0 3.0 1e-06 
3.0 3.238 0 3.0 1e-06 
0.05 3.239 0 3.0 1e-06 
3.0 3.239 0 3.0 1e-06 
0.05 3.24 0 3.0 1e-06 
3.0 3.24 0 3.0 1e-06 
0.05 3.241 0 3.0 1e-06 
3.0 3.241 0 3.0 1e-06 
0.05 3.242 0 3.0 1e-06 
3.0 3.242 0 3.0 1e-06 
0.05 3.243 0 3.0 1e-06 
3.0 3.243 0 3.0 1e-06 
0.05 3.244 0 3.0 1e-06 
3.0 3.244 0 3.0 1e-06 
0.05 3.245 0 3.0 1e-06 
3.0 3.245 0 3.0 1e-06 
0.05 3.246 0 3.0 1e-06 
3.0 3.246 0 3.0 1e-06 
0.05 3.247 0 3.0 1e-06 
3.0 3.247 0 3.0 1e-06 
0.05 3.248 0 3.0 1e-06 
3.0 3.248 0 3.0 1e-06 
0.05 3.249 0 3.0 1e-06 
3.0 3.249 0 3.0 1e-06 
0.05 3.25 0 3.0 1e-06 
3.0 3.25 0 3.0 1e-06 
0.05 3.251 0 3.0 1e-06 
3.0 3.251 0 3.0 1e-06 
0.05 3.252 0 3.0 1e-06 
3.0 3.252 0 3.0 1e-06 
0.05 3.253 0 3.0 1e-06 
3.0 3.253 0 3.0 1e-06 
0.05 3.254 0 3.0 1e-06 
3.0 3.254 0 3.0 1e-06 
0.05 3.255 0 3.0 1e-06 
3.0 3.255 0 3.0 1e-06 
0.05 3.256 0 3.0 1e-06 
3.0 3.256 0 3.0 1e-06 
0.05 3.257 0 3.0 1e-06 
3.0 3.257 0 3.0 1e-06 
0.05 3.258 0 3.0 1e-06 
3.0 3.258 0 3.0 1e-06 
0.05 3.259 0 3.0 1e-06 
3.0 3.259 0 3.0 1e-06 
0.05 3.26 0 3.0 1e-06 
3.0 3.26 0 3.0 1e-06 
0.05 3.261 0 3.0 1e-06 
3.0 3.261 0 3.0 1e-06 
0.05 3.262 0 3.0 1e-06 
3.0 3.262 0 3.0 1e-06 
0.05 3.263 0 3.0 1e-06 
3.0 3.263 0 3.0 1e-06 
0.05 3.264 0 3.0 1e-06 
3.0 3.264 0 3.0 1e-06 
0.05 3.265 0 3.0 1e-06 
3.0 3.265 0 3.0 1e-06 
0.05 3.266 0 3.0 1e-06 
3.0 3.266 0 3.0 1e-06 
0.05 3.267 0 3.0 1e-06 
3.0 3.267 0 3.0 1e-06 
0.05 3.268 0 3.0 1e-06 
3.0 3.268 0 3.0 1e-06 
0.05 3.269 0 3.0 1e-06 
3.0 3.269 0 3.0 1e-06 
0.05 3.27 0 3.0 1e-06 
3.0 3.27 0 3.0 1e-06 
0.05 3.271 0 3.0 1e-06 
3.0 3.271 0 3.0 1e-06 
0.05 3.272 0 3.0 1e-06 
3.0 3.272 0 3.0 1e-06 
0.05 3.273 0 3.0 1e-06 
3.0 3.273 0 3.0 1e-06 
0.05 3.274 0 3.0 1e-06 
3.0 3.274 0 3.0 1e-06 
0.05 3.275 0 3.0 1e-06 
3.0 3.275 0 3.0 1e-06 
0.05 3.276 0 3.0 1e-06 
3.0 3.276 0 3.0 1e-06 
0.05 3.277 0 3.0 1e-06 
3.0 3.277 0 3.0 1e-06 
0.05 3.278 0 3.0 1e-06 
3.0 3.278 0 3.0 1e-06 
0.05 3.279 0 3.0 1e-06 
3.0 3.279 0 3.0 1e-06 
0.05 3.28 0 3.0 1e-06 
3.0 3.28 0 3.0 1e-06 
0.05 3.281 0 3.0 1e-06 
3.0 3.281 0 3.0 1e-06 
0.05 3.282 0 3.0 1e-06 
3.0 3.282 0 3.0 1e-06 
0.05 3.283 0 3.0 1e-06 
3.0 3.283 0 3.0 1e-06 
0.05 3.284 0 3.0 1e-06 
3.0 3.284 0 3.0 1e-06 
0.05 3.285 0 3.0 1e-06 
3.0 3.285 0 3.0 1e-06 
0.05 3.286 0 3.0 1e-06 
3.0 3.286 0 3.0 1e-06 
0.05 3.287 0 3.0 1e-06 
3.0 3.287 0 3.0 1e-06 
0.05 3.288 0 3.0 1e-06 
3.0 3.288 0 3.0 1e-06 
0.05 3.289 0 3.0 1e-06 
3.0 3.289 0 3.0 1e-06 
0.05 3.29 0 3.0 1e-06 
3.0 3.29 0 3.0 1e-06 
0.05 3.291 0 3.0 1e-06 
3.0 3.291 0 3.0 1e-06 
0.05 3.292 0 3.0 1e-06 
3.0 3.292 0 3.0 1e-06 
0.05 3.293 0 3.0 1e-06 
3.0 3.293 0 3.0 1e-06 
0.05 3.294 0 3.0 1e-06 
3.0 3.294 0 3.0 1e-06 
0.05 3.295 0 3.0 1e-06 
3.0 3.295 0 3.0 1e-06 
0.05 3.296 0 3.0 1e-06 
3.0 3.296 0 3.0 1e-06 
0.05 3.297 0 3.0 1e-06 
3.0 3.297 0 3.0 1e-06 
0.05 3.298 0 3.0 1e-06 
3.0 3.298 0 3.0 1e-06 
0.05 3.299 0 3.0 1e-06 
3.0 3.299 0 3.0 1e-06 
0.05 3.3 0 3.0 1e-06 
3.0 3.3 0 3.0 1e-06 
0.05 3.301 0 3.0 1e-06 
3.0 3.301 0 3.0 1e-06 
0.05 3.302 0 3.0 1e-06 
3.0 3.302 0 3.0 1e-06 
0.05 3.303 0 3.0 1e-06 
3.0 3.303 0 3.0 1e-06 
0.05 3.304 0 3.0 1e-06 
3.0 3.304 0 3.0 1e-06 
0.05 3.305 0 3.0 1e-06 
3.0 3.305 0 3.0 1e-06 
0.05 3.306 0 3.0 1e-06 
3.0 3.306 0 3.0 1e-06 
0.05 3.307 0 3.0 1e-06 
3.0 3.307 0 3.0 1e-06 
0.05 3.308 0 3.0 1e-06 
3.0 3.308 0 3.0 1e-06 
0.05 3.309 0 3.0 1e-06 
3.0 3.309 0 3.0 1e-06 
0.05 3.31 0 3.0 1e-06 
3.0 3.31 0 3.0 1e-06 
0.05 3.311 0 3.0 1e-06 
3.0 3.311 0 3.0 1e-06 
0.05 3.312 0 3.0 1e-06 
3.0 3.312 0 3.0 1e-06 
0.05 3.313 0 3.0 1e-06 
3.0 3.313 0 3.0 1e-06 
0.05 3.314 0 3.0 1e-06 
3.0 3.314 0 3.0 1e-06 
0.05 3.315 0 3.0 1e-06 
3.0 3.315 0 3.0 1e-06 
0.05 3.316 0 3.0 1e-06 
3.0 3.316 0 3.0 1e-06 
0.05 3.317 0 3.0 1e-06 
3.0 3.317 0 3.0 1e-06 
0.05 3.318 0 3.0 1e-06 
3.0 3.318 0 3.0 1e-06 
0.05 3.319 0 3.0 1e-06 
3.0 3.319 0 3.0 1e-06 
0.05 3.32 0 3.0 1e-06 
3.0 3.32 0 3.0 1e-06 
0.05 3.321 0 3.0 1e-06 
3.0 3.321 0 3.0 1e-06 
0.05 3.322 0 3.0 1e-06 
3.0 3.322 0 3.0 1e-06 
0.05 3.323 0 3.0 1e-06 
3.0 3.323 0 3.0 1e-06 
0.05 3.324 0 3.0 1e-06 
3.0 3.324 0 3.0 1e-06 
0.05 3.325 0 3.0 1e-06 
3.0 3.325 0 3.0 1e-06 
0.05 3.326 0 3.0 1e-06 
3.0 3.326 0 3.0 1e-06 
0.05 3.327 0 3.0 1e-06 
3.0 3.327 0 3.0 1e-06 
0.05 3.328 0 3.0 1e-06 
3.0 3.328 0 3.0 1e-06 
0.05 3.329 0 3.0 1e-06 
3.0 3.329 0 3.0 1e-06 
0.05 3.33 0 3.0 1e-06 
3.0 3.33 0 3.0 1e-06 
0.05 3.331 0 3.0 1e-06 
3.0 3.331 0 3.0 1e-06 
0.05 3.332 0 3.0 1e-06 
3.0 3.332 0 3.0 1e-06 
0.05 3.333 0 3.0 1e-06 
3.0 3.333 0 3.0 1e-06 
0.05 3.334 0 3.0 1e-06 
3.0 3.334 0 3.0 1e-06 
0.05 3.335 0 3.0 1e-06 
3.0 3.335 0 3.0 1e-06 
0.05 3.336 0 3.0 1e-06 
3.0 3.336 0 3.0 1e-06 
0.05 3.337 0 3.0 1e-06 
3.0 3.337 0 3.0 1e-06 
0.05 3.338 0 3.0 1e-06 
3.0 3.338 0 3.0 1e-06 
0.05 3.339 0 3.0 1e-06 
3.0 3.339 0 3.0 1e-06 
0.05 3.34 0 3.0 1e-06 
3.0 3.34 0 3.0 1e-06 
0.05 3.341 0 3.0 1e-06 
3.0 3.341 0 3.0 1e-06 
0.05 3.342 0 3.0 1e-06 
3.0 3.342 0 3.0 1e-06 
0.05 3.343 0 3.0 1e-06 
3.0 3.343 0 3.0 1e-06 
0.05 3.344 0 3.0 1e-06 
3.0 3.344 0 3.0 1e-06 
0.05 3.345 0 3.0 1e-06 
3.0 3.345 0 3.0 1e-06 
0.05 3.346 0 3.0 1e-06 
3.0 3.346 0 3.0 1e-06 
0.05 3.347 0 3.0 1e-06 
3.0 3.347 0 3.0 1e-06 
0.05 3.348 0 3.0 1e-06 
3.0 3.348 0 3.0 1e-06 
0.05 3.349 0 3.0 1e-06 
3.0 3.349 0 3.0 1e-06 
0.05 3.35 0 3.0 1e-06 
3.0 3.35 0 3.0 1e-06 
0.05 3.351 0 3.0 1e-06 
3.0 3.351 0 3.0 1e-06 
0.05 3.352 0 3.0 1e-06 
3.0 3.352 0 3.0 1e-06 
0.05 3.353 0 3.0 1e-06 
3.0 3.353 0 3.0 1e-06 
0.05 3.354 0 3.0 1e-06 
3.0 3.354 0 3.0 1e-06 
0.05 3.355 0 3.0 1e-06 
3.0 3.355 0 3.0 1e-06 
0.05 3.356 0 3.0 1e-06 
3.0 3.356 0 3.0 1e-06 
0.05 3.357 0 3.0 1e-06 
3.0 3.357 0 3.0 1e-06 
0.05 3.358 0 3.0 1e-06 
3.0 3.358 0 3.0 1e-06 
0.05 3.359 0 3.0 1e-06 
3.0 3.359 0 3.0 1e-06 
0.05 3.36 0 3.0 1e-06 
3.0 3.36 0 3.0 1e-06 
0.05 3.361 0 3.0 1e-06 
3.0 3.361 0 3.0 1e-06 
0.05 3.362 0 3.0 1e-06 
3.0 3.362 0 3.0 1e-06 
0.05 3.363 0 3.0 1e-06 
3.0 3.363 0 3.0 1e-06 
0.05 3.364 0 3.0 1e-06 
3.0 3.364 0 3.0 1e-06 
0.05 3.365 0 3.0 1e-06 
3.0 3.365 0 3.0 1e-06 
0.05 3.366 0 3.0 1e-06 
3.0 3.366 0 3.0 1e-06 
0.05 3.367 0 3.0 1e-06 
3.0 3.367 0 3.0 1e-06 
0.05 3.368 0 3.0 1e-06 
3.0 3.368 0 3.0 1e-06 
0.05 3.369 0 3.0 1e-06 
3.0 3.369 0 3.0 1e-06 
0.05 3.37 0 3.0 1e-06 
3.0 3.37 0 3.0 1e-06 
0.05 3.371 0 3.0 1e-06 
3.0 3.371 0 3.0 1e-06 
0.05 3.372 0 3.0 1e-06 
3.0 3.372 0 3.0 1e-06 
0.05 3.373 0 3.0 1e-06 
3.0 3.373 0 3.0 1e-06 
0.05 3.374 0 3.0 1e-06 
3.0 3.374 0 3.0 1e-06 
0.05 3.375 0 3.0 1e-06 
3.0 3.375 0 3.0 1e-06 
0.05 3.376 0 3.0 1e-06 
3.0 3.376 0 3.0 1e-06 
0.05 3.377 0 3.0 1e-06 
3.0 3.377 0 3.0 1e-06 
0.05 3.378 0 3.0 1e-06 
3.0 3.378 0 3.0 1e-06 
0.05 3.379 0 3.0 1e-06 
3.0 3.379 0 3.0 1e-06 
0.05 3.38 0 3.0 1e-06 
3.0 3.38 0 3.0 1e-06 
0.05 3.381 0 3.0 1e-06 
3.0 3.381 0 3.0 1e-06 
0.05 3.382 0 3.0 1e-06 
3.0 3.382 0 3.0 1e-06 
0.05 3.383 0 3.0 1e-06 
3.0 3.383 0 3.0 1e-06 
0.05 3.384 0 3.0 1e-06 
3.0 3.384 0 3.0 1e-06 
0.05 3.385 0 3.0 1e-06 
3.0 3.385 0 3.0 1e-06 
0.05 3.386 0 3.0 1e-06 
3.0 3.386 0 3.0 1e-06 
0.05 3.387 0 3.0 1e-06 
3.0 3.387 0 3.0 1e-06 
0.05 3.388 0 3.0 1e-06 
3.0 3.388 0 3.0 1e-06 
0.05 3.389 0 3.0 1e-06 
3.0 3.389 0 3.0 1e-06 
0.05 3.39 0 3.0 1e-06 
3.0 3.39 0 3.0 1e-06 
0.05 3.391 0 3.0 1e-06 
3.0 3.391 0 3.0 1e-06 
0.05 3.392 0 3.0 1e-06 
3.0 3.392 0 3.0 1e-06 
0.05 3.393 0 3.0 1e-06 
3.0 3.393 0 3.0 1e-06 
0.05 3.394 0 3.0 1e-06 
3.0 3.394 0 3.0 1e-06 
0.05 3.395 0 3.0 1e-06 
3.0 3.395 0 3.0 1e-06 
0.05 3.396 0 3.0 1e-06 
3.0 3.396 0 3.0 1e-06 
0.05 3.397 0 3.0 1e-06 
3.0 3.397 0 3.0 1e-06 
0.05 3.398 0 3.0 1e-06 
3.0 3.398 0 3.0 1e-06 
0.05 3.399 0 3.0 1e-06 
3.0 3.399 0 3.0 1e-06 
0.05 3.4 0 3.0 1e-06 
3.0 3.4 0 3.0 1e-06 
0.05 3.401 0 3.0 1e-06 
3.0 3.401 0 3.0 1e-06 
0.05 3.402 0 3.0 1e-06 
3.0 3.402 0 3.0 1e-06 
0.05 3.403 0 3.0 1e-06 
3.0 3.403 0 3.0 1e-06 
0.05 3.404 0 3.0 1e-06 
3.0 3.404 0 3.0 1e-06 
0.05 3.405 0 3.0 1e-06 
3.0 3.405 0 3.0 1e-06 
0.05 3.406 0 3.0 1e-06 
3.0 3.406 0 3.0 1e-06 
0.05 3.407 0 3.0 1e-06 
3.0 3.407 0 3.0 1e-06 
0.05 3.408 0 3.0 1e-06 
3.0 3.408 0 3.0 1e-06 
0.05 3.409 0 3.0 1e-06 
3.0 3.409 0 3.0 1e-06 
0.05 3.41 0 3.0 1e-06 
3.0 3.41 0 3.0 1e-06 
0.05 3.411 0 3.0 1e-06 
3.0 3.411 0 3.0 1e-06 
0.05 3.412 0 3.0 1e-06 
3.0 3.412 0 3.0 1e-06 
0.05 3.413 0 3.0 1e-06 
3.0 3.413 0 3.0 1e-06 
0.05 3.414 0 3.0 1e-06 
3.0 3.414 0 3.0 1e-06 
0.05 3.415 0 3.0 1e-06 
3.0 3.415 0 3.0 1e-06 
0.05 3.416 0 3.0 1e-06 
3.0 3.416 0 3.0 1e-06 
0.05 3.417 0 3.0 1e-06 
3.0 3.417 0 3.0 1e-06 
0.05 3.418 0 3.0 1e-06 
3.0 3.418 0 3.0 1e-06 
0.05 3.419 0 3.0 1e-06 
3.0 3.419 0 3.0 1e-06 
0.05 3.42 0 3.0 1e-06 
3.0 3.42 0 3.0 1e-06 
0.05 3.421 0 3.0 1e-06 
3.0 3.421 0 3.0 1e-06 
0.05 3.422 0 3.0 1e-06 
3.0 3.422 0 3.0 1e-06 
0.05 3.423 0 3.0 1e-06 
3.0 3.423 0 3.0 1e-06 
0.05 3.424 0 3.0 1e-06 
3.0 3.424 0 3.0 1e-06 
0.05 3.425 0 3.0 1e-06 
3.0 3.425 0 3.0 1e-06 
0.05 3.426 0 3.0 1e-06 
3.0 3.426 0 3.0 1e-06 
0.05 3.427 0 3.0 1e-06 
3.0 3.427 0 3.0 1e-06 
0.05 3.428 0 3.0 1e-06 
3.0 3.428 0 3.0 1e-06 
0.05 3.429 0 3.0 1e-06 
3.0 3.429 0 3.0 1e-06 
0.05 3.43 0 3.0 1e-06 
3.0 3.43 0 3.0 1e-06 
0.05 3.431 0 3.0 1e-06 
3.0 3.431 0 3.0 1e-06 
0.05 3.432 0 3.0 1e-06 
3.0 3.432 0 3.0 1e-06 
0.05 3.433 0 3.0 1e-06 
3.0 3.433 0 3.0 1e-06 
0.05 3.434 0 3.0 1e-06 
3.0 3.434 0 3.0 1e-06 
0.05 3.435 0 3.0 1e-06 
3.0 3.435 0 3.0 1e-06 
0.05 3.436 0 3.0 1e-06 
3.0 3.436 0 3.0 1e-06 
0.05 3.437 0 3.0 1e-06 
3.0 3.437 0 3.0 1e-06 
0.05 3.438 0 3.0 1e-06 
3.0 3.438 0 3.0 1e-06 
0.05 3.439 0 3.0 1e-06 
3.0 3.439 0 3.0 1e-06 
0.05 3.44 0 3.0 1e-06 
3.0 3.44 0 3.0 1e-06 
0.05 3.441 0 3.0 1e-06 
3.0 3.441 0 3.0 1e-06 
0.05 3.442 0 3.0 1e-06 
3.0 3.442 0 3.0 1e-06 
0.05 3.443 0 3.0 1e-06 
3.0 3.443 0 3.0 1e-06 
0.05 3.444 0 3.0 1e-06 
3.0 3.444 0 3.0 1e-06 
0.05 3.445 0 3.0 1e-06 
3.0 3.445 0 3.0 1e-06 
0.05 3.446 0 3.0 1e-06 
3.0 3.446 0 3.0 1e-06 
0.05 3.447 0 3.0 1e-06 
3.0 3.447 0 3.0 1e-06 
0.05 3.448 0 3.0 1e-06 
3.0 3.448 0 3.0 1e-06 
0.05 3.449 0 3.0 1e-06 
3.0 3.449 0 3.0 1e-06 
0.05 3.45 0 3.0 1e-06 
3.0 3.45 0 3.0 1e-06 
0.05 3.451 0 3.0 1e-06 
3.0 3.451 0 3.0 1e-06 
0.05 3.452 0 3.0 1e-06 
3.0 3.452 0 3.0 1e-06 
0.05 3.453 0 3.0 1e-06 
3.0 3.453 0 3.0 1e-06 
0.05 3.454 0 3.0 1e-06 
3.0 3.454 0 3.0 1e-06 
0.05 3.455 0 3.0 1e-06 
3.0 3.455 0 3.0 1e-06 
0.05 3.456 0 3.0 1e-06 
3.0 3.456 0 3.0 1e-06 
0.05 3.457 0 3.0 1e-06 
3.0 3.457 0 3.0 1e-06 
0.05 3.458 0 3.0 1e-06 
3.0 3.458 0 3.0 1e-06 
0.05 3.459 0 3.0 1e-06 
3.0 3.459 0 3.0 1e-06 
0.05 3.46 0 3.0 1e-06 
3.0 3.46 0 3.0 1e-06 
0.05 3.461 0 3.0 1e-06 
3.0 3.461 0 3.0 1e-06 
0.05 3.462 0 3.0 1e-06 
3.0 3.462 0 3.0 1e-06 
0.05 3.463 0 3.0 1e-06 
3.0 3.463 0 3.0 1e-06 
0.05 3.464 0 3.0 1e-06 
3.0 3.464 0 3.0 1e-06 
0.05 3.465 0 3.0 1e-06 
3.0 3.465 0 3.0 1e-06 
0.05 3.466 0 3.0 1e-06 
3.0 3.466 0 3.0 1e-06 
0.05 3.467 0 3.0 1e-06 
3.0 3.467 0 3.0 1e-06 
0.05 3.468 0 3.0 1e-06 
3.0 3.468 0 3.0 1e-06 
0.05 3.469 0 3.0 1e-06 
3.0 3.469 0 3.0 1e-06 
0.05 3.47 0 3.0 1e-06 
3.0 3.47 0 3.0 1e-06 
0.05 3.471 0 3.0 1e-06 
3.0 3.471 0 3.0 1e-06 
0.05 3.472 0 3.0 1e-06 
3.0 3.472 0 3.0 1e-06 
0.05 3.473 0 3.0 1e-06 
3.0 3.473 0 3.0 1e-06 
0.05 3.474 0 3.0 1e-06 
3.0 3.474 0 3.0 1e-06 
0.05 3.475 0 3.0 1e-06 
3.0 3.475 0 3.0 1e-06 
0.05 3.476 0 3.0 1e-06 
3.0 3.476 0 3.0 1e-06 
0.05 3.477 0 3.0 1e-06 
3.0 3.477 0 3.0 1e-06 
0.05 3.478 0 3.0 1e-06 
3.0 3.478 0 3.0 1e-06 
0.05 3.479 0 3.0 1e-06 
3.0 3.479 0 3.0 1e-06 
0.05 3.48 0 3.0 1e-06 
3.0 3.48 0 3.0 1e-06 
0.05 3.481 0 3.0 1e-06 
3.0 3.481 0 3.0 1e-06 
0.05 3.482 0 3.0 1e-06 
3.0 3.482 0 3.0 1e-06 
0.05 3.483 0 3.0 1e-06 
3.0 3.483 0 3.0 1e-06 
0.05 3.484 0 3.0 1e-06 
3.0 3.484 0 3.0 1e-06 
0.05 3.485 0 3.0 1e-06 
3.0 3.485 0 3.0 1e-06 
0.05 3.486 0 3.0 1e-06 
3.0 3.486 0 3.0 1e-06 
0.05 3.487 0 3.0 1e-06 
3.0 3.487 0 3.0 1e-06 
0.05 3.488 0 3.0 1e-06 
3.0 3.488 0 3.0 1e-06 
0.05 3.489 0 3.0 1e-06 
3.0 3.489 0 3.0 1e-06 
0.05 3.49 0 3.0 1e-06 
3.0 3.49 0 3.0 1e-06 
0.05 3.491 0 3.0 1e-06 
3.0 3.491 0 3.0 1e-06 
0.05 3.492 0 3.0 1e-06 
3.0 3.492 0 3.0 1e-06 
0.05 3.493 0 3.0 1e-06 
3.0 3.493 0 3.0 1e-06 
0.05 3.494 0 3.0 1e-06 
3.0 3.494 0 3.0 1e-06 
0.05 3.495 0 3.0 1e-06 
3.0 3.495 0 3.0 1e-06 
0.05 3.496 0 3.0 1e-06 
3.0 3.496 0 3.0 1e-06 
0.05 3.497 0 3.0 1e-06 
3.0 3.497 0 3.0 1e-06 
0.05 3.498 0 3.0 1e-06 
3.0 3.498 0 3.0 1e-06 
0.05 3.499 0 3.0 1e-06 
3.0 3.499 0 3.0 1e-06 
0.05 3.5 0 3.0 1e-06 
3.0 3.5 0 3.0 1e-06 
0.05 3.501 0 3.0 1e-06 
3.0 3.501 0 3.0 1e-06 
0.05 3.502 0 3.0 1e-06 
3.0 3.502 0 3.0 1e-06 
0.05 3.503 0 3.0 1e-06 
3.0 3.503 0 3.0 1e-06 
0.05 3.504 0 3.0 1e-06 
3.0 3.504 0 3.0 1e-06 
0.05 3.505 0 3.0 1e-06 
3.0 3.505 0 3.0 1e-06 
0.05 3.506 0 3.0 1e-06 
3.0 3.506 0 3.0 1e-06 
0.05 3.507 0 3.0 1e-06 
3.0 3.507 0 3.0 1e-06 
0.05 3.508 0 3.0 1e-06 
3.0 3.508 0 3.0 1e-06 
0.05 3.509 0 3.0 1e-06 
3.0 3.509 0 3.0 1e-06 
0.05 3.51 0 3.0 1e-06 
3.0 3.51 0 3.0 1e-06 
0.05 3.511 0 3.0 1e-06 
3.0 3.511 0 3.0 1e-06 
0.05 3.512 0 3.0 1e-06 
3.0 3.512 0 3.0 1e-06 
0.05 3.513 0 3.0 1e-06 
3.0 3.513 0 3.0 1e-06 
0.05 3.514 0 3.0 1e-06 
3.0 3.514 0 3.0 1e-06 
0.05 3.515 0 3.0 1e-06 
3.0 3.515 0 3.0 1e-06 
0.05 3.516 0 3.0 1e-06 
3.0 3.516 0 3.0 1e-06 
0.05 3.517 0 3.0 1e-06 
3.0 3.517 0 3.0 1e-06 
0.05 3.518 0 3.0 1e-06 
3.0 3.518 0 3.0 1e-06 
0.05 3.519 0 3.0 1e-06 
3.0 3.519 0 3.0 1e-06 
0.05 3.52 0 3.0 1e-06 
3.0 3.52 0 3.0 1e-06 
0.05 3.521 0 3.0 1e-06 
3.0 3.521 0 3.0 1e-06 
0.05 3.522 0 3.0 1e-06 
3.0 3.522 0 3.0 1e-06 
0.05 3.523 0 3.0 1e-06 
3.0 3.523 0 3.0 1e-06 
0.05 3.524 0 3.0 1e-06 
3.0 3.524 0 3.0 1e-06 
0.05 3.525 0 3.0 1e-06 
3.0 3.525 0 3.0 1e-06 
0.05 3.526 0 3.0 1e-06 
3.0 3.526 0 3.0 1e-06 
0.05 3.527 0 3.0 1e-06 
3.0 3.527 0 3.0 1e-06 
0.05 3.528 0 3.0 1e-06 
3.0 3.528 0 3.0 1e-06 
0.05 3.529 0 3.0 1e-06 
3.0 3.529 0 3.0 1e-06 
0.05 3.53 0 3.0 1e-06 
3.0 3.53 0 3.0 1e-06 
0.05 3.531 0 3.0 1e-06 
3.0 3.531 0 3.0 1e-06 
0.05 3.532 0 3.0 1e-06 
3.0 3.532 0 3.0 1e-06 
0.05 3.533 0 3.0 1e-06 
3.0 3.533 0 3.0 1e-06 
0.05 3.534 0 3.0 1e-06 
3.0 3.534 0 3.0 1e-06 
0.05 3.535 0 3.0 1e-06 
3.0 3.535 0 3.0 1e-06 
0.05 3.536 0 3.0 1e-06 
3.0 3.536 0 3.0 1e-06 
0.05 3.537 0 3.0 1e-06 
3.0 3.537 0 3.0 1e-06 
0.05 3.538 0 3.0 1e-06 
3.0 3.538 0 3.0 1e-06 
0.05 3.539 0 3.0 1e-06 
3.0 3.539 0 3.0 1e-06 
0.05 3.54 0 3.0 1e-06 
3.0 3.54 0 3.0 1e-06 
0.05 3.541 0 3.0 1e-06 
3.0 3.541 0 3.0 1e-06 
0.05 3.542 0 3.0 1e-06 
3.0 3.542 0 3.0 1e-06 
0.05 3.543 0 3.0 1e-06 
3.0 3.543 0 3.0 1e-06 
0.05 3.544 0 3.0 1e-06 
3.0 3.544 0 3.0 1e-06 
0.05 3.545 0 3.0 1e-06 
3.0 3.545 0 3.0 1e-06 
0.05 3.546 0 3.0 1e-06 
3.0 3.546 0 3.0 1e-06 
0.05 3.547 0 3.0 1e-06 
3.0 3.547 0 3.0 1e-06 
0.05 3.548 0 3.0 1e-06 
3.0 3.548 0 3.0 1e-06 
0.05 3.549 0 3.0 1e-06 
3.0 3.549 0 3.0 1e-06 
0.05 3.55 0 3.0 1e-06 
3.0 3.55 0 3.0 1e-06 
0.05 3.551 0 3.0 1e-06 
3.0 3.551 0 3.0 1e-06 
0.05 3.552 0 3.0 1e-06 
3.0 3.552 0 3.0 1e-06 
0.05 3.553 0 3.0 1e-06 
3.0 3.553 0 3.0 1e-06 
0.05 3.554 0 3.0 1e-06 
3.0 3.554 0 3.0 1e-06 
0.05 3.555 0 3.0 1e-06 
3.0 3.555 0 3.0 1e-06 
0.05 3.556 0 3.0 1e-06 
3.0 3.556 0 3.0 1e-06 
0.05 3.557 0 3.0 1e-06 
3.0 3.557 0 3.0 1e-06 
0.05 3.558 0 3.0 1e-06 
3.0 3.558 0 3.0 1e-06 
0.05 3.559 0 3.0 1e-06 
3.0 3.559 0 3.0 1e-06 
0.05 3.56 0 3.0 1e-06 
3.0 3.56 0 3.0 1e-06 
0.05 3.561 0 3.0 1e-06 
3.0 3.561 0 3.0 1e-06 
0.05 3.562 0 3.0 1e-06 
3.0 3.562 0 3.0 1e-06 
0.05 3.563 0 3.0 1e-06 
3.0 3.563 0 3.0 1e-06 
0.05 3.564 0 3.0 1e-06 
3.0 3.564 0 3.0 1e-06 
0.05 3.565 0 3.0 1e-06 
3.0 3.565 0 3.0 1e-06 
0.05 3.566 0 3.0 1e-06 
3.0 3.566 0 3.0 1e-06 
0.05 3.567 0 3.0 1e-06 
3.0 3.567 0 3.0 1e-06 
0.05 3.568 0 3.0 1e-06 
3.0 3.568 0 3.0 1e-06 
0.05 3.569 0 3.0 1e-06 
3.0 3.569 0 3.0 1e-06 
0.05 3.57 0 3.0 1e-06 
3.0 3.57 0 3.0 1e-06 
0.05 3.571 0 3.0 1e-06 
3.0 3.571 0 3.0 1e-06 
0.05 3.572 0 3.0 1e-06 
3.0 3.572 0 3.0 1e-06 
0.05 3.573 0 3.0 1e-06 
3.0 3.573 0 3.0 1e-06 
0.05 3.574 0 3.0 1e-06 
3.0 3.574 0 3.0 1e-06 
0.05 3.575 0 3.0 1e-06 
3.0 3.575 0 3.0 1e-06 
0.05 3.576 0 3.0 1e-06 
3.0 3.576 0 3.0 1e-06 
0.05 3.577 0 3.0 1e-06 
3.0 3.577 0 3.0 1e-06 
0.05 3.578 0 3.0 1e-06 
3.0 3.578 0 3.0 1e-06 
0.05 3.579 0 3.0 1e-06 
3.0 3.579 0 3.0 1e-06 
0.05 3.58 0 3.0 1e-06 
3.0 3.58 0 3.0 1e-06 
0.05 3.581 0 3.0 1e-06 
3.0 3.581 0 3.0 1e-06 
0.05 3.582 0 3.0 1e-06 
3.0 3.582 0 3.0 1e-06 
0.05 3.583 0 3.0 1e-06 
3.0 3.583 0 3.0 1e-06 
0.05 3.584 0 3.0 1e-06 
3.0 3.584 0 3.0 1e-06 
0.05 3.585 0 3.0 1e-06 
3.0 3.585 0 3.0 1e-06 
0.05 3.586 0 3.0 1e-06 
3.0 3.586 0 3.0 1e-06 
0.05 3.587 0 3.0 1e-06 
3.0 3.587 0 3.0 1e-06 
0.05 3.588 0 3.0 1e-06 
3.0 3.588 0 3.0 1e-06 
0.05 3.589 0 3.0 1e-06 
3.0 3.589 0 3.0 1e-06 
0.05 3.59 0 3.0 1e-06 
3.0 3.59 0 3.0 1e-06 
0.05 3.591 0 3.0 1e-06 
3.0 3.591 0 3.0 1e-06 
0.05 3.592 0 3.0 1e-06 
3.0 3.592 0 3.0 1e-06 
0.05 3.593 0 3.0 1e-06 
3.0 3.593 0 3.0 1e-06 
0.05 3.594 0 3.0 1e-06 
3.0 3.594 0 3.0 1e-06 
0.05 3.595 0 3.0 1e-06 
3.0 3.595 0 3.0 1e-06 
0.05 3.596 0 3.0 1e-06 
3.0 3.596 0 3.0 1e-06 
0.05 3.597 0 3.0 1e-06 
3.0 3.597 0 3.0 1e-06 
0.05 3.598 0 3.0 1e-06 
3.0 3.598 0 3.0 1e-06 
0.05 3.599 0 3.0 1e-06 
3.0 3.599 0 3.0 1e-06 
0.05 3.6 0 3.0 1e-06 
3.0 3.6 0 3.0 1e-06 
0.05 3.601 0 3.0 1e-06 
3.0 3.601 0 3.0 1e-06 
0.05 3.602 0 3.0 1e-06 
3.0 3.602 0 3.0 1e-06 
0.05 3.603 0 3.0 1e-06 
3.0 3.603 0 3.0 1e-06 
0.05 3.604 0 3.0 1e-06 
3.0 3.604 0 3.0 1e-06 
0.05 3.605 0 3.0 1e-06 
3.0 3.605 0 3.0 1e-06 
0.05 3.606 0 3.0 1e-06 
3.0 3.606 0 3.0 1e-06 
0.05 3.607 0 3.0 1e-06 
3.0 3.607 0 3.0 1e-06 
0.05 3.608 0 3.0 1e-06 
3.0 3.608 0 3.0 1e-06 
0.05 3.609 0 3.0 1e-06 
3.0 3.609 0 3.0 1e-06 
0.05 3.61 0 3.0 1e-06 
3.0 3.61 0 3.0 1e-06 
0.05 3.611 0 3.0 1e-06 
3.0 3.611 0 3.0 1e-06 
0.05 3.612 0 3.0 1e-06 
3.0 3.612 0 3.0 1e-06 
0.05 3.613 0 3.0 1e-06 
3.0 3.613 0 3.0 1e-06 
0.05 3.614 0 3.0 1e-06 
3.0 3.614 0 3.0 1e-06 
0.05 3.615 0 3.0 1e-06 
3.0 3.615 0 3.0 1e-06 
0.05 3.616 0 3.0 1e-06 
3.0 3.616 0 3.0 1e-06 
0.05 3.617 0 3.0 1e-06 
3.0 3.617 0 3.0 1e-06 
0.05 3.618 0 3.0 1e-06 
3.0 3.618 0 3.0 1e-06 
0.05 3.619 0 3.0 1e-06 
3.0 3.619 0 3.0 1e-06 
0.05 3.62 0 3.0 1e-06 
3.0 3.62 0 3.0 1e-06 
0.05 3.621 0 3.0 1e-06 
3.0 3.621 0 3.0 1e-06 
0.05 3.622 0 3.0 1e-06 
3.0 3.622 0 3.0 1e-06 
0.05 3.623 0 3.0 1e-06 
3.0 3.623 0 3.0 1e-06 
0.05 3.624 0 3.0 1e-06 
3.0 3.624 0 3.0 1e-06 
0.05 3.625 0 3.0 1e-06 
3.0 3.625 0 3.0 1e-06 
0.05 3.626 0 3.0 1e-06 
3.0 3.626 0 3.0 1e-06 
0.05 3.627 0 3.0 1e-06 
3.0 3.627 0 3.0 1e-06 
0.05 3.628 0 3.0 1e-06 
3.0 3.628 0 3.0 1e-06 
0.05 3.629 0 3.0 1e-06 
3.0 3.629 0 3.0 1e-06 
0.05 3.63 0 3.0 1e-06 
3.0 3.63 0 3.0 1e-06 
0.05 3.631 0 3.0 1e-06 
3.0 3.631 0 3.0 1e-06 
0.05 3.632 0 3.0 1e-06 
3.0 3.632 0 3.0 1e-06 
0.05 3.633 0 3.0 1e-06 
3.0 3.633 0 3.0 1e-06 
0.05 3.634 0 3.0 1e-06 
3.0 3.634 0 3.0 1e-06 
0.05 3.635 0 3.0 1e-06 
3.0 3.635 0 3.0 1e-06 
0.05 3.636 0 3.0 1e-06 
3.0 3.636 0 3.0 1e-06 
0.05 3.637 0 3.0 1e-06 
3.0 3.637 0 3.0 1e-06 
0.05 3.638 0 3.0 1e-06 
3.0 3.638 0 3.0 1e-06 
0.05 3.639 0 3.0 1e-06 
3.0 3.639 0 3.0 1e-06 
0.05 3.64 0 3.0 1e-06 
3.0 3.64 0 3.0 1e-06 
0.05 3.641 0 3.0 1e-06 
3.0 3.641 0 3.0 1e-06 
0.05 3.642 0 3.0 1e-06 
3.0 3.642 0 3.0 1e-06 
0.05 3.643 0 3.0 1e-06 
3.0 3.643 0 3.0 1e-06 
0.05 3.644 0 3.0 1e-06 
3.0 3.644 0 3.0 1e-06 
0.05 3.645 0 3.0 1e-06 
3.0 3.645 0 3.0 1e-06 
0.05 3.646 0 3.0 1e-06 
3.0 3.646 0 3.0 1e-06 
0.05 3.647 0 3.0 1e-06 
3.0 3.647 0 3.0 1e-06 
0.05 3.648 0 3.0 1e-06 
3.0 3.648 0 3.0 1e-06 
0.05 3.649 0 3.0 1e-06 
3.0 3.649 0 3.0 1e-06 
0.05 3.65 0 3.0 1e-06 
3.0 3.65 0 3.0 1e-06 
0.05 3.651 0 3.0 1e-06 
3.0 3.651 0 3.0 1e-06 
0.05 3.652 0 3.0 1e-06 
3.0 3.652 0 3.0 1e-06 
0.05 3.653 0 3.0 1e-06 
3.0 3.653 0 3.0 1e-06 
0.05 3.654 0 3.0 1e-06 
3.0 3.654 0 3.0 1e-06 
0.05 3.655 0 3.0 1e-06 
3.0 3.655 0 3.0 1e-06 
0.05 3.656 0 3.0 1e-06 
3.0 3.656 0 3.0 1e-06 
0.05 3.657 0 3.0 1e-06 
3.0 3.657 0 3.0 1e-06 
0.05 3.658 0 3.0 1e-06 
3.0 3.658 0 3.0 1e-06 
0.05 3.659 0 3.0 1e-06 
3.0 3.659 0 3.0 1e-06 
0.05 3.66 0 3.0 1e-06 
3.0 3.66 0 3.0 1e-06 
0.05 3.661 0 3.0 1e-06 
3.0 3.661 0 3.0 1e-06 
0.05 3.662 0 3.0 1e-06 
3.0 3.662 0 3.0 1e-06 
0.05 3.663 0 3.0 1e-06 
3.0 3.663 0 3.0 1e-06 
0.05 3.664 0 3.0 1e-06 
3.0 3.664 0 3.0 1e-06 
0.05 3.665 0 3.0 1e-06 
3.0 3.665 0 3.0 1e-06 
0.05 3.666 0 3.0 1e-06 
3.0 3.666 0 3.0 1e-06 
0.05 3.667 0 3.0 1e-06 
3.0 3.667 0 3.0 1e-06 
0.05 3.668 0 3.0 1e-06 
3.0 3.668 0 3.0 1e-06 
0.05 3.669 0 3.0 1e-06 
3.0 3.669 0 3.0 1e-06 
0.05 3.67 0 3.0 1e-06 
3.0 3.67 0 3.0 1e-06 
0.05 3.671 0 3.0 1e-06 
3.0 3.671 0 3.0 1e-06 
0.05 3.672 0 3.0 1e-06 
3.0 3.672 0 3.0 1e-06 
0.05 3.673 0 3.0 1e-06 
3.0 3.673 0 3.0 1e-06 
0.05 3.674 0 3.0 1e-06 
3.0 3.674 0 3.0 1e-06 
0.05 3.675 0 3.0 1e-06 
3.0 3.675 0 3.0 1e-06 
0.05 3.676 0 3.0 1e-06 
3.0 3.676 0 3.0 1e-06 
0.05 3.677 0 3.0 1e-06 
3.0 3.677 0 3.0 1e-06 
0.05 3.678 0 3.0 1e-06 
3.0 3.678 0 3.0 1e-06 
0.05 3.679 0 3.0 1e-06 
3.0 3.679 0 3.0 1e-06 
0.05 3.68 0 3.0 1e-06 
3.0 3.68 0 3.0 1e-06 
0.05 3.681 0 3.0 1e-06 
3.0 3.681 0 3.0 1e-06 
0.05 3.682 0 3.0 1e-06 
3.0 3.682 0 3.0 1e-06 
0.05 3.683 0 3.0 1e-06 
3.0 3.683 0 3.0 1e-06 
0.05 3.684 0 3.0 1e-06 
3.0 3.684 0 3.0 1e-06 
0.05 3.685 0 3.0 1e-06 
3.0 3.685 0 3.0 1e-06 
0.05 3.686 0 3.0 1e-06 
3.0 3.686 0 3.0 1e-06 
0.05 3.687 0 3.0 1e-06 
3.0 3.687 0 3.0 1e-06 
0.05 3.688 0 3.0 1e-06 
3.0 3.688 0 3.0 1e-06 
0.05 3.689 0 3.0 1e-06 
3.0 3.689 0 3.0 1e-06 
0.05 3.69 0 3.0 1e-06 
3.0 3.69 0 3.0 1e-06 
0.05 3.691 0 3.0 1e-06 
3.0 3.691 0 3.0 1e-06 
0.05 3.692 0 3.0 1e-06 
3.0 3.692 0 3.0 1e-06 
0.05 3.693 0 3.0 1e-06 
3.0 3.693 0 3.0 1e-06 
0.05 3.694 0 3.0 1e-06 
3.0 3.694 0 3.0 1e-06 
0.05 3.695 0 3.0 1e-06 
3.0 3.695 0 3.0 1e-06 
0.05 3.696 0 3.0 1e-06 
3.0 3.696 0 3.0 1e-06 
0.05 3.697 0 3.0 1e-06 
3.0 3.697 0 3.0 1e-06 
0.05 3.698 0 3.0 1e-06 
3.0 3.698 0 3.0 1e-06 
0.05 3.699 0 3.0 1e-06 
3.0 3.699 0 3.0 1e-06 
0.05 3.7 0 3.0 1e-06 
3.0 3.7 0 3.0 1e-06 
0.05 3.701 0 3.0 1e-06 
3.0 3.701 0 3.0 1e-06 
0.05 3.702 0 3.0 1e-06 
3.0 3.702 0 3.0 1e-06 
0.05 3.703 0 3.0 1e-06 
3.0 3.703 0 3.0 1e-06 
0.05 3.704 0 3.0 1e-06 
3.0 3.704 0 3.0 1e-06 
0.05 3.705 0 3.0 1e-06 
3.0 3.705 0 3.0 1e-06 
0.05 3.706 0 3.0 1e-06 
3.0 3.706 0 3.0 1e-06 
0.05 3.707 0 3.0 1e-06 
3.0 3.707 0 3.0 1e-06 
0.05 3.708 0 3.0 1e-06 
3.0 3.708 0 3.0 1e-06 
0.05 3.709 0 3.0 1e-06 
3.0 3.709 0 3.0 1e-06 
0.05 3.71 0 3.0 1e-06 
3.0 3.71 0 3.0 1e-06 
0.05 3.711 0 3.0 1e-06 
3.0 3.711 0 3.0 1e-06 
0.05 3.712 0 3.0 1e-06 
3.0 3.712 0 3.0 1e-06 
0.05 3.713 0 3.0 1e-06 
3.0 3.713 0 3.0 1e-06 
0.05 3.714 0 3.0 1e-06 
3.0 3.714 0 3.0 1e-06 
0.05 3.715 0 3.0 1e-06 
3.0 3.715 0 3.0 1e-06 
0.05 3.716 0 3.0 1e-06 
3.0 3.716 0 3.0 1e-06 
0.05 3.717 0 3.0 1e-06 
3.0 3.717 0 3.0 1e-06 
0.05 3.718 0 3.0 1e-06 
3.0 3.718 0 3.0 1e-06 
0.05 3.719 0 3.0 1e-06 
3.0 3.719 0 3.0 1e-06 
0.05 3.72 0 3.0 1e-06 
3.0 3.72 0 3.0 1e-06 
0.05 3.721 0 3.0 1e-06 
3.0 3.721 0 3.0 1e-06 
0.05 3.722 0 3.0 1e-06 
3.0 3.722 0 3.0 1e-06 
0.05 3.723 0 3.0 1e-06 
3.0 3.723 0 3.0 1e-06 
0.05 3.724 0 3.0 1e-06 
3.0 3.724 0 3.0 1e-06 
0.05 3.725 0 3.0 1e-06 
3.0 3.725 0 3.0 1e-06 
0.05 3.726 0 3.0 1e-06 
3.0 3.726 0 3.0 1e-06 
0.05 3.727 0 3.0 1e-06 
3.0 3.727 0 3.0 1e-06 
0.05 3.728 0 3.0 1e-06 
3.0 3.728 0 3.0 1e-06 
0.05 3.729 0 3.0 1e-06 
3.0 3.729 0 3.0 1e-06 
0.05 3.73 0 3.0 1e-06 
3.0 3.73 0 3.0 1e-06 
0.05 3.731 0 3.0 1e-06 
3.0 3.731 0 3.0 1e-06 
0.05 3.732 0 3.0 1e-06 
3.0 3.732 0 3.0 1e-06 
0.05 3.733 0 3.0 1e-06 
3.0 3.733 0 3.0 1e-06 
0.05 3.734 0 3.0 1e-06 
3.0 3.734 0 3.0 1e-06 
0.05 3.735 0 3.0 1e-06 
3.0 3.735 0 3.0 1e-06 
0.05 3.736 0 3.0 1e-06 
3.0 3.736 0 3.0 1e-06 
0.05 3.737 0 3.0 1e-06 
3.0 3.737 0 3.0 1e-06 
0.05 3.738 0 3.0 1e-06 
3.0 3.738 0 3.0 1e-06 
0.05 3.739 0 3.0 1e-06 
3.0 3.739 0 3.0 1e-06 
0.05 3.74 0 3.0 1e-06 
3.0 3.74 0 3.0 1e-06 
0.05 3.741 0 3.0 1e-06 
3.0 3.741 0 3.0 1e-06 
0.05 3.742 0 3.0 1e-06 
3.0 3.742 0 3.0 1e-06 
0.05 3.743 0 3.0 1e-06 
3.0 3.743 0 3.0 1e-06 
0.05 3.744 0 3.0 1e-06 
3.0 3.744 0 3.0 1e-06 
0.05 3.745 0 3.0 1e-06 
3.0 3.745 0 3.0 1e-06 
0.05 3.746 0 3.0 1e-06 
3.0 3.746 0 3.0 1e-06 
0.05 3.747 0 3.0 1e-06 
3.0 3.747 0 3.0 1e-06 
0.05 3.748 0 3.0 1e-06 
3.0 3.748 0 3.0 1e-06 
0.05 3.749 0 3.0 1e-06 
3.0 3.749 0 3.0 1e-06 
0.05 3.75 0 3.0 1e-06 
3.0 3.75 0 3.0 1e-06 
0.05 3.751 0 3.0 1e-06 
3.0 3.751 0 3.0 1e-06 
0.05 3.752 0 3.0 1e-06 
3.0 3.752 0 3.0 1e-06 
0.05 3.753 0 3.0 1e-06 
3.0 3.753 0 3.0 1e-06 
0.05 3.754 0 3.0 1e-06 
3.0 3.754 0 3.0 1e-06 
0.05 3.755 0 3.0 1e-06 
3.0 3.755 0 3.0 1e-06 
0.05 3.756 0 3.0 1e-06 
3.0 3.756 0 3.0 1e-06 
0.05 3.757 0 3.0 1e-06 
3.0 3.757 0 3.0 1e-06 
0.05 3.758 0 3.0 1e-06 
3.0 3.758 0 3.0 1e-06 
0.05 3.759 0 3.0 1e-06 
3.0 3.759 0 3.0 1e-06 
0.05 3.76 0 3.0 1e-06 
3.0 3.76 0 3.0 1e-06 
0.05 3.761 0 3.0 1e-06 
3.0 3.761 0 3.0 1e-06 
0.05 3.762 0 3.0 1e-06 
3.0 3.762 0 3.0 1e-06 
0.05 3.763 0 3.0 1e-06 
3.0 3.763 0 3.0 1e-06 
0.05 3.764 0 3.0 1e-06 
3.0 3.764 0 3.0 1e-06 
0.05 3.765 0 3.0 1e-06 
3.0 3.765 0 3.0 1e-06 
0.05 3.766 0 3.0 1e-06 
3.0 3.766 0 3.0 1e-06 
0.05 3.767 0 3.0 1e-06 
3.0 3.767 0 3.0 1e-06 
0.05 3.768 0 3.0 1e-06 
3.0 3.768 0 3.0 1e-06 
0.05 3.769 0 3.0 1e-06 
3.0 3.769 0 3.0 1e-06 
0.05 3.77 0 3.0 1e-06 
3.0 3.77 0 3.0 1e-06 
0.05 3.771 0 3.0 1e-06 
3.0 3.771 0 3.0 1e-06 
0.05 3.772 0 3.0 1e-06 
3.0 3.772 0 3.0 1e-06 
0.05 3.773 0 3.0 1e-06 
3.0 3.773 0 3.0 1e-06 
0.05 3.774 0 3.0 1e-06 
3.0 3.774 0 3.0 1e-06 
0.05 3.775 0 3.0 1e-06 
3.0 3.775 0 3.0 1e-06 
0.05 3.776 0 3.0 1e-06 
3.0 3.776 0 3.0 1e-06 
0.05 3.777 0 3.0 1e-06 
3.0 3.777 0 3.0 1e-06 
0.05 3.778 0 3.0 1e-06 
3.0 3.778 0 3.0 1e-06 
0.05 3.779 0 3.0 1e-06 
3.0 3.779 0 3.0 1e-06 
0.05 3.78 0 3.0 1e-06 
3.0 3.78 0 3.0 1e-06 
0.05 3.781 0 3.0 1e-06 
3.0 3.781 0 3.0 1e-06 
0.05 3.782 0 3.0 1e-06 
3.0 3.782 0 3.0 1e-06 
0.05 3.783 0 3.0 1e-06 
3.0 3.783 0 3.0 1e-06 
0.05 3.784 0 3.0 1e-06 
3.0 3.784 0 3.0 1e-06 
0.05 3.785 0 3.0 1e-06 
3.0 3.785 0 3.0 1e-06 
0.05 3.786 0 3.0 1e-06 
3.0 3.786 0 3.0 1e-06 
0.05 3.787 0 3.0 1e-06 
3.0 3.787 0 3.0 1e-06 
0.05 3.788 0 3.0 1e-06 
3.0 3.788 0 3.0 1e-06 
0.05 3.789 0 3.0 1e-06 
3.0 3.789 0 3.0 1e-06 
0.05 3.79 0 3.0 1e-06 
3.0 3.79 0 3.0 1e-06 
0.05 3.791 0 3.0 1e-06 
3.0 3.791 0 3.0 1e-06 
0.05 3.792 0 3.0 1e-06 
3.0 3.792 0 3.0 1e-06 
0.05 3.793 0 3.0 1e-06 
3.0 3.793 0 3.0 1e-06 
0.05 3.794 0 3.0 1e-06 
3.0 3.794 0 3.0 1e-06 
0.05 3.795 0 3.0 1e-06 
3.0 3.795 0 3.0 1e-06 
0.05 3.796 0 3.0 1e-06 
3.0 3.796 0 3.0 1e-06 
0.05 3.797 0 3.0 1e-06 
3.0 3.797 0 3.0 1e-06 
0.05 3.798 0 3.0 1e-06 
3.0 3.798 0 3.0 1e-06 
0.05 3.799 0 3.0 1e-06 
3.0 3.799 0 3.0 1e-06 
0.05 3.8 0 3.0 1e-06 
3.0 3.8 0 3.0 1e-06 
0.05 3.801 0 3.0 1e-06 
3.0 3.801 0 3.0 1e-06 
0.05 3.802 0 3.0 1e-06 
3.0 3.802 0 3.0 1e-06 
0.05 3.803 0 3.0 1e-06 
3.0 3.803 0 3.0 1e-06 
0.05 3.804 0 3.0 1e-06 
3.0 3.804 0 3.0 1e-06 
0.05 3.805 0 3.0 1e-06 
3.0 3.805 0 3.0 1e-06 
0.05 3.806 0 3.0 1e-06 
3.0 3.806 0 3.0 1e-06 
0.05 3.807 0 3.0 1e-06 
3.0 3.807 0 3.0 1e-06 
0.05 3.808 0 3.0 1e-06 
3.0 3.808 0 3.0 1e-06 
0.05 3.809 0 3.0 1e-06 
3.0 3.809 0 3.0 1e-06 
0.05 3.81 0 3.0 1e-06 
3.0 3.81 0 3.0 1e-06 
0.05 3.811 0 3.0 1e-06 
3.0 3.811 0 3.0 1e-06 
0.05 3.812 0 3.0 1e-06 
3.0 3.812 0 3.0 1e-06 
0.05 3.813 0 3.0 1e-06 
3.0 3.813 0 3.0 1e-06 
0.05 3.814 0 3.0 1e-06 
3.0 3.814 0 3.0 1e-06 
0.05 3.815 0 3.0 1e-06 
3.0 3.815 0 3.0 1e-06 
0.05 3.816 0 3.0 1e-06 
3.0 3.816 0 3.0 1e-06 
0.05 3.817 0 3.0 1e-06 
3.0 3.817 0 3.0 1e-06 
0.05 3.818 0 3.0 1e-06 
3.0 3.818 0 3.0 1e-06 
0.05 3.819 0 3.0 1e-06 
3.0 3.819 0 3.0 1e-06 
0.05 3.82 0 3.0 1e-06 
3.0 3.82 0 3.0 1e-06 
0.05 3.821 0 3.0 1e-06 
3.0 3.821 0 3.0 1e-06 
0.05 3.822 0 3.0 1e-06 
3.0 3.822 0 3.0 1e-06 
0.05 3.823 0 3.0 1e-06 
3.0 3.823 0 3.0 1e-06 
0.05 3.824 0 3.0 1e-06 
3.0 3.824 0 3.0 1e-06 
0.05 3.825 0 3.0 1e-06 
3.0 3.825 0 3.0 1e-06 
0.05 3.826 0 3.0 1e-06 
3.0 3.826 0 3.0 1e-06 
0.05 3.827 0 3.0 1e-06 
3.0 3.827 0 3.0 1e-06 
0.05 3.828 0 3.0 1e-06 
3.0 3.828 0 3.0 1e-06 
0.05 3.829 0 3.0 1e-06 
3.0 3.829 0 3.0 1e-06 
0.05 3.83 0 3.0 1e-06 
3.0 3.83 0 3.0 1e-06 
0.05 3.831 0 3.0 1e-06 
3.0 3.831 0 3.0 1e-06 
0.05 3.832 0 3.0 1e-06 
3.0 3.832 0 3.0 1e-06 
0.05 3.833 0 3.0 1e-06 
3.0 3.833 0 3.0 1e-06 
0.05 3.834 0 3.0 1e-06 
3.0 3.834 0 3.0 1e-06 
0.05 3.835 0 3.0 1e-06 
3.0 3.835 0 3.0 1e-06 
0.05 3.836 0 3.0 1e-06 
3.0 3.836 0 3.0 1e-06 
0.05 3.837 0 3.0 1e-06 
3.0 3.837 0 3.0 1e-06 
0.05 3.838 0 3.0 1e-06 
3.0 3.838 0 3.0 1e-06 
0.05 3.839 0 3.0 1e-06 
3.0 3.839 0 3.0 1e-06 
0.05 3.84 0 3.0 1e-06 
3.0 3.84 0 3.0 1e-06 
0.05 3.841 0 3.0 1e-06 
3.0 3.841 0 3.0 1e-06 
0.05 3.842 0 3.0 1e-06 
3.0 3.842 0 3.0 1e-06 
0.05 3.843 0 3.0 1e-06 
3.0 3.843 0 3.0 1e-06 
0.05 3.844 0 3.0 1e-06 
3.0 3.844 0 3.0 1e-06 
0.05 3.845 0 3.0 1e-06 
3.0 3.845 0 3.0 1e-06 
0.05 3.846 0 3.0 1e-06 
3.0 3.846 0 3.0 1e-06 
0.05 3.847 0 3.0 1e-06 
3.0 3.847 0 3.0 1e-06 
0.05 3.848 0 3.0 1e-06 
3.0 3.848 0 3.0 1e-06 
0.05 3.849 0 3.0 1e-06 
3.0 3.849 0 3.0 1e-06 
0.05 3.85 0 3.0 1e-06 
3.0 3.85 0 3.0 1e-06 
0.05 3.851 0 3.0 1e-06 
3.0 3.851 0 3.0 1e-06 
0.05 3.852 0 3.0 1e-06 
3.0 3.852 0 3.0 1e-06 
0.05 3.853 0 3.0 1e-06 
3.0 3.853 0 3.0 1e-06 
0.05 3.854 0 3.0 1e-06 
3.0 3.854 0 3.0 1e-06 
0.05 3.855 0 3.0 1e-06 
3.0 3.855 0 3.0 1e-06 
0.05 3.856 0 3.0 1e-06 
3.0 3.856 0 3.0 1e-06 
0.05 3.857 0 3.0 1e-06 
3.0 3.857 0 3.0 1e-06 
0.05 3.858 0 3.0 1e-06 
3.0 3.858 0 3.0 1e-06 
0.05 3.859 0 3.0 1e-06 
3.0 3.859 0 3.0 1e-06 
0.05 3.86 0 3.0 1e-06 
3.0 3.86 0 3.0 1e-06 
0.05 3.861 0 3.0 1e-06 
3.0 3.861 0 3.0 1e-06 
0.05 3.862 0 3.0 1e-06 
3.0 3.862 0 3.0 1e-06 
0.05 3.863 0 3.0 1e-06 
3.0 3.863 0 3.0 1e-06 
0.05 3.864 0 3.0 1e-06 
3.0 3.864 0 3.0 1e-06 
0.05 3.865 0 3.0 1e-06 
3.0 3.865 0 3.0 1e-06 
0.05 3.866 0 3.0 1e-06 
3.0 3.866 0 3.0 1e-06 
0.05 3.867 0 3.0 1e-06 
3.0 3.867 0 3.0 1e-06 
0.05 3.868 0 3.0 1e-06 
3.0 3.868 0 3.0 1e-06 
0.05 3.869 0 3.0 1e-06 
3.0 3.869 0 3.0 1e-06 
0.05 3.87 0 3.0 1e-06 
3.0 3.87 0 3.0 1e-06 
0.05 3.871 0 3.0 1e-06 
3.0 3.871 0 3.0 1e-06 
0.05 3.872 0 3.0 1e-06 
3.0 3.872 0 3.0 1e-06 
0.05 3.873 0 3.0 1e-06 
3.0 3.873 0 3.0 1e-06 
0.05 3.874 0 3.0 1e-06 
3.0 3.874 0 3.0 1e-06 
0.05 3.875 0 3.0 1e-06 
3.0 3.875 0 3.0 1e-06 
0.05 3.876 0 3.0 1e-06 
3.0 3.876 0 3.0 1e-06 
0.05 3.877 0 3.0 1e-06 
3.0 3.877 0 3.0 1e-06 
0.05 3.878 0 3.0 1e-06 
3.0 3.878 0 3.0 1e-06 
0.05 3.879 0 3.0 1e-06 
3.0 3.879 0 3.0 1e-06 
0.05 3.88 0 3.0 1e-06 
3.0 3.88 0 3.0 1e-06 
0.05 3.881 0 3.0 1e-06 
3.0 3.881 0 3.0 1e-06 
0.05 3.882 0 3.0 1e-06 
3.0 3.882 0 3.0 1e-06 
0.05 3.883 0 3.0 1e-06 
3.0 3.883 0 3.0 1e-06 
0.05 3.884 0 3.0 1e-06 
3.0 3.884 0 3.0 1e-06 
0.05 3.885 0 3.0 1e-06 
3.0 3.885 0 3.0 1e-06 
0.05 3.886 0 3.0 1e-06 
3.0 3.886 0 3.0 1e-06 
0.05 3.887 0 3.0 1e-06 
3.0 3.887 0 3.0 1e-06 
0.05 3.888 0 3.0 1e-06 
3.0 3.888 0 3.0 1e-06 
0.05 3.889 0 3.0 1e-06 
3.0 3.889 0 3.0 1e-06 
0.05 3.89 0 3.0 1e-06 
3.0 3.89 0 3.0 1e-06 
0.05 3.891 0 3.0 1e-06 
3.0 3.891 0 3.0 1e-06 
0.05 3.892 0 3.0 1e-06 
3.0 3.892 0 3.0 1e-06 
0.05 3.893 0 3.0 1e-06 
3.0 3.893 0 3.0 1e-06 
0.05 3.894 0 3.0 1e-06 
3.0 3.894 0 3.0 1e-06 
0.05 3.895 0 3.0 1e-06 
3.0 3.895 0 3.0 1e-06 
0.05 3.896 0 3.0 1e-06 
3.0 3.896 0 3.0 1e-06 
0.05 3.897 0 3.0 1e-06 
3.0 3.897 0 3.0 1e-06 
0.05 3.898 0 3.0 1e-06 
3.0 3.898 0 3.0 1e-06 
0.05 3.899 0 3.0 1e-06 
3.0 3.899 0 3.0 1e-06 
0.05 3.9 0 3.0 1e-06 
3.0 3.9 0 3.0 1e-06 
0.05 3.901 0 3.0 1e-06 
3.0 3.901 0 3.0 1e-06 
0.05 3.902 0 3.0 1e-06 
3.0 3.902 0 3.0 1e-06 
0.05 3.903 0 3.0 1e-06 
3.0 3.903 0 3.0 1e-06 
0.05 3.904 0 3.0 1e-06 
3.0 3.904 0 3.0 1e-06 
0.05 3.905 0 3.0 1e-06 
3.0 3.905 0 3.0 1e-06 
0.05 3.906 0 3.0 1e-06 
3.0 3.906 0 3.0 1e-06 
0.05 3.907 0 3.0 1e-06 
3.0 3.907 0 3.0 1e-06 
0.05 3.908 0 3.0 1e-06 
3.0 3.908 0 3.0 1e-06 
0.05 3.909 0 3.0 1e-06 
3.0 3.909 0 3.0 1e-06 
0.05 3.91 0 3.0 1e-06 
3.0 3.91 0 3.0 1e-06 
0.05 3.911 0 3.0 1e-06 
3.0 3.911 0 3.0 1e-06 
0.05 3.912 0 3.0 1e-06 
3.0 3.912 0 3.0 1e-06 
0.05 3.913 0 3.0 1e-06 
3.0 3.913 0 3.0 1e-06 
0.05 3.914 0 3.0 1e-06 
3.0 3.914 0 3.0 1e-06 
0.05 3.915 0 3.0 1e-06 
3.0 3.915 0 3.0 1e-06 
0.05 3.916 0 3.0 1e-06 
3.0 3.916 0 3.0 1e-06 
0.05 3.917 0 3.0 1e-06 
3.0 3.917 0 3.0 1e-06 
0.05 3.918 0 3.0 1e-06 
3.0 3.918 0 3.0 1e-06 
0.05 3.919 0 3.0 1e-06 
3.0 3.919 0 3.0 1e-06 
0.05 3.92 0 3.0 1e-06 
3.0 3.92 0 3.0 1e-06 
0.05 3.921 0 3.0 1e-06 
3.0 3.921 0 3.0 1e-06 
0.05 3.922 0 3.0 1e-06 
3.0 3.922 0 3.0 1e-06 
0.05 3.923 0 3.0 1e-06 
3.0 3.923 0 3.0 1e-06 
0.05 3.924 0 3.0 1e-06 
3.0 3.924 0 3.0 1e-06 
0.05 3.925 0 3.0 1e-06 
3.0 3.925 0 3.0 1e-06 
0.05 3.926 0 3.0 1e-06 
3.0 3.926 0 3.0 1e-06 
0.05 3.927 0 3.0 1e-06 
3.0 3.927 0 3.0 1e-06 
0.05 3.928 0 3.0 1e-06 
3.0 3.928 0 3.0 1e-06 
0.05 3.929 0 3.0 1e-06 
3.0 3.929 0 3.0 1e-06 
0.05 3.93 0 3.0 1e-06 
3.0 3.93 0 3.0 1e-06 
0.05 3.931 0 3.0 1e-06 
3.0 3.931 0 3.0 1e-06 
0.05 3.932 0 3.0 1e-06 
3.0 3.932 0 3.0 1e-06 
0.05 3.933 0 3.0 1e-06 
3.0 3.933 0 3.0 1e-06 
0.05 3.934 0 3.0 1e-06 
3.0 3.934 0 3.0 1e-06 
0.05 3.935 0 3.0 1e-06 
3.0 3.935 0 3.0 1e-06 
0.05 3.936 0 3.0 1e-06 
3.0 3.936 0 3.0 1e-06 
0.05 3.937 0 3.0 1e-06 
3.0 3.937 0 3.0 1e-06 
0.05 3.938 0 3.0 1e-06 
3.0 3.938 0 3.0 1e-06 
0.05 3.939 0 3.0 1e-06 
3.0 3.939 0 3.0 1e-06 
0.05 3.94 0 3.0 1e-06 
3.0 3.94 0 3.0 1e-06 
0.05 3.941 0 3.0 1e-06 
3.0 3.941 0 3.0 1e-06 
0.05 3.942 0 3.0 1e-06 
3.0 3.942 0 3.0 1e-06 
0.05 3.943 0 3.0 1e-06 
3.0 3.943 0 3.0 1e-06 
0.05 3.944 0 3.0 1e-06 
3.0 3.944 0 3.0 1e-06 
0.05 3.945 0 3.0 1e-06 
3.0 3.945 0 3.0 1e-06 
0.05 3.946 0 3.0 1e-06 
3.0 3.946 0 3.0 1e-06 
0.05 3.947 0 3.0 1e-06 
3.0 3.947 0 3.0 1e-06 
0.05 3.948 0 3.0 1e-06 
3.0 3.948 0 3.0 1e-06 
0.05 3.949 0 3.0 1e-06 
3.0 3.949 0 3.0 1e-06 
0.05 3.95 0 3.0 1e-06 
3.0 3.95 0 3.0 1e-06 
0.05 3.951 0 3.0 1e-06 
3.0 3.951 0 3.0 1e-06 
0.05 3.952 0 3.0 1e-06 
3.0 3.952 0 3.0 1e-06 
0.05 3.953 0 3.0 1e-06 
3.0 3.953 0 3.0 1e-06 
0.05 3.954 0 3.0 1e-06 
3.0 3.954 0 3.0 1e-06 
0.05 3.955 0 3.0 1e-06 
3.0 3.955 0 3.0 1e-06 
0.05 3.956 0 3.0 1e-06 
3.0 3.956 0 3.0 1e-06 
0.05 3.957 0 3.0 1e-06 
3.0 3.957 0 3.0 1e-06 
0.05 3.958 0 3.0 1e-06 
3.0 3.958 0 3.0 1e-06 
0.05 3.959 0 3.0 1e-06 
3.0 3.959 0 3.0 1e-06 
0.05 3.96 0 3.0 1e-06 
3.0 3.96 0 3.0 1e-06 
0.05 3.961 0 3.0 1e-06 
3.0 3.961 0 3.0 1e-06 
0.05 3.962 0 3.0 1e-06 
3.0 3.962 0 3.0 1e-06 
0.05 3.963 0 3.0 1e-06 
3.0 3.963 0 3.0 1e-06 
0.05 3.964 0 3.0 1e-06 
3.0 3.964 0 3.0 1e-06 
0.05 3.965 0 3.0 1e-06 
3.0 3.965 0 3.0 1e-06 
0.05 3.966 0 3.0 1e-06 
3.0 3.966 0 3.0 1e-06 
0.05 3.967 0 3.0 1e-06 
3.0 3.967 0 3.0 1e-06 
0.05 3.968 0 3.0 1e-06 
3.0 3.968 0 3.0 1e-06 
0.05 3.969 0 3.0 1e-06 
3.0 3.969 0 3.0 1e-06 
0.05 3.97 0 3.0 1e-06 
3.0 3.97 0 3.0 1e-06 
0.05 3.971 0 3.0 1e-06 
3.0 3.971 0 3.0 1e-06 
0.05 3.972 0 3.0 1e-06 
3.0 3.972 0 3.0 1e-06 
0.05 3.973 0 3.0 1e-06 
3.0 3.973 0 3.0 1e-06 
0.05 3.974 0 3.0 1e-06 
3.0 3.974 0 3.0 1e-06 
0.05 3.975 0 3.0 1e-06 
3.0 3.975 0 3.0 1e-06 
0.05 3.976 0 3.0 1e-06 
3.0 3.976 0 3.0 1e-06 
0.05 3.977 0 3.0 1e-06 
3.0 3.977 0 3.0 1e-06 
0.05 3.978 0 3.0 1e-06 
3.0 3.978 0 3.0 1e-06 
0.05 3.979 0 3.0 1e-06 
3.0 3.979 0 3.0 1e-06 
0.05 3.98 0 3.0 1e-06 
3.0 3.98 0 3.0 1e-06 
0.05 3.981 0 3.0 1e-06 
3.0 3.981 0 3.0 1e-06 
0.05 3.982 0 3.0 1e-06 
3.0 3.982 0 3.0 1e-06 
0.05 3.983 0 3.0 1e-06 
3.0 3.983 0 3.0 1e-06 
0.05 3.984 0 3.0 1e-06 
3.0 3.984 0 3.0 1e-06 
0.05 3.985 0 3.0 1e-06 
3.0 3.985 0 3.0 1e-06 
0.05 3.986 0 3.0 1e-06 
3.0 3.986 0 3.0 1e-06 
0.05 3.987 0 3.0 1e-06 
3.0 3.987 0 3.0 1e-06 
0.05 3.988 0 3.0 1e-06 
3.0 3.988 0 3.0 1e-06 
0.05 3.989 0 3.0 1e-06 
3.0 3.989 0 3.0 1e-06 
0.05 3.99 0 3.0 1e-06 
3.0 3.99 0 3.0 1e-06 
0.05 3.991 0 3.0 1e-06 
3.0 3.991 0 3.0 1e-06 
0.05 3.992 0 3.0 1e-06 
3.0 3.992 0 3.0 1e-06 
0.05 3.993 0 3.0 1e-06 
3.0 3.993 0 3.0 1e-06 
0.05 3.994 0 3.0 1e-06 
3.0 3.994 0 3.0 1e-06 
0.05 3.995 0 3.0 1e-06 
3.0 3.995 0 3.0 1e-06 
0.05 3.996 0 3.0 1e-06 
3.0 3.996 0 3.0 1e-06 
0.05 3.997 0 3.0 1e-06 
3.0 3.997 0 3.0 1e-06 
0.05 3.998 0 3.0 1e-06 
3.0 3.998 0 3.0 1e-06 
0.05 3.999 0 3.0 1e-06 
3.0 3.999 0 3.0 1e-06 
0.05 4.0 0 3.0 1e-06 
3.0 4.0 0 3.0 1e-06 
0.05 4.001 0 3.0 1e-06 
3.0 4.001 0 3.0 1e-06 
0.05 4.002 0 3.0 1e-06 
3.0 4.002 0 3.0 1e-06 
0.05 4.003 0 3.0 1e-06 
3.0 4.003 0 3.0 1e-06 
0.05 4.004 0 3.0 1e-06 
3.0 4.004 0 3.0 1e-06 
0.05 4.005 0 3.0 1e-06 
3.0 4.005 0 3.0 1e-06 
0.05 4.006 0 3.0 1e-06 
3.0 4.006 0 3.0 1e-06 
0.05 4.007 0 3.0 1e-06 
3.0 4.007 0 3.0 1e-06 
0.05 4.008 0 3.0 1e-06 
3.0 4.008 0 3.0 1e-06 
0.05 4.009 0 3.0 1e-06 
3.0 4.009 0 3.0 1e-06 
0.05 4.01 0 3.0 1e-06 
3.0 4.01 0 3.0 1e-06 
0.05 4.011 0 3.0 1e-06 
3.0 4.011 0 3.0 1e-06 
0.05 4.012 0 3.0 1e-06 
3.0 4.012 0 3.0 1e-06 
0.05 4.013 0 3.0 1e-06 
3.0 4.013 0 3.0 1e-06 
0.05 4.014 0 3.0 1e-06 
3.0 4.014 0 3.0 1e-06 
0.05 4.015 0 3.0 1e-06 
3.0 4.015 0 3.0 1e-06 
0.05 4.016 0 3.0 1e-06 
3.0 4.016 0 3.0 1e-06 
0.05 4.017 0 3.0 1e-06 
3.0 4.017 0 3.0 1e-06 
0.05 4.018 0 3.0 1e-06 
3.0 4.018 0 3.0 1e-06 
0.05 4.019 0 3.0 1e-06 
3.0 4.019 0 3.0 1e-06 
0.05 4.02 0 3.0 1e-06 
3.0 4.02 0 3.0 1e-06 
0.05 4.021 0 3.0 1e-06 
3.0 4.021 0 3.0 1e-06 
0.05 4.022 0 3.0 1e-06 
3.0 4.022 0 3.0 1e-06 
0.05 4.023 0 3.0 1e-06 
3.0 4.023 0 3.0 1e-06 
0.05 4.024 0 3.0 1e-06 
3.0 4.024 0 3.0 1e-06 
0.05 4.025 0 3.0 1e-06 
3.0 4.025 0 3.0 1e-06 
0.05 4.026 0 3.0 1e-06 
3.0 4.026 0 3.0 1e-06 
0.05 4.027 0 3.0 1e-06 
3.0 4.027 0 3.0 1e-06 
0.05 4.028 0 3.0 1e-06 
3.0 4.028 0 3.0 1e-06 
0.05 4.029 0 3.0 1e-06 
3.0 4.029 0 3.0 1e-06 
0.05 4.03 0 3.0 1e-06 
3.0 4.03 0 3.0 1e-06 
0.05 4.031 0 3.0 1e-06 
3.0 4.031 0 3.0 1e-06 
0.05 4.032 0 3.0 1e-06 
3.0 4.032 0 3.0 1e-06 
0.05 4.033 0 3.0 1e-06 
3.0 4.033 0 3.0 1e-06 
0.05 4.034 0 3.0 1e-06 
3.0 4.034 0 3.0 1e-06 
0.05 4.035 0 3.0 1e-06 
3.0 4.035 0 3.0 1e-06 
0.05 4.036 0 3.0 1e-06 
3.0 4.036 0 3.0 1e-06 
0.05 4.037 0 3.0 1e-06 
3.0 4.037 0 3.0 1e-06 
0.05 4.038 0 3.0 1e-06 
3.0 4.038 0 3.0 1e-06 
0.05 4.039 0 3.0 1e-06 
3.0 4.039 0 3.0 1e-06 
0.05 4.04 0 3.0 1e-06 
3.0 4.04 0 3.0 1e-06 
0.05 4.041 0 3.0 1e-06 
3.0 4.041 0 3.0 1e-06 
0.05 4.042 0 3.0 1e-06 
3.0 4.042 0 3.0 1e-06 
0.05 4.043 0 3.0 1e-06 
3.0 4.043 0 3.0 1e-06 
0.05 4.044 0 3.0 1e-06 
3.0 4.044 0 3.0 1e-06 
0.05 4.045 0 3.0 1e-06 
3.0 4.045 0 3.0 1e-06 
0.05 4.046 0 3.0 1e-06 
3.0 4.046 0 3.0 1e-06 
0.05 4.047 0 3.0 1e-06 
3.0 4.047 0 3.0 1e-06 
0.05 4.048 0 3.0 1e-06 
3.0 4.048 0 3.0 1e-06 
0.05 4.049 0 3.0 1e-06 
3.0 4.049 0 3.0 1e-06 
0.05 4.05 0 3.0 1e-06 
3.0 4.05 0 3.0 1e-06 
0.05 4.051 0 3.0 1e-06 
3.0 4.051 0 3.0 1e-06 
0.05 4.052 0 3.0 1e-06 
3.0 4.052 0 3.0 1e-06 
0.05 4.053 0 3.0 1e-06 
3.0 4.053 0 3.0 1e-06 
0.05 4.054 0 3.0 1e-06 
3.0 4.054 0 3.0 1e-06 
0.05 4.055 0 3.0 1e-06 
3.0 4.055 0 3.0 1e-06 
0.05 4.056 0 3.0 1e-06 
3.0 4.056 0 3.0 1e-06 
0.05 4.057 0 3.0 1e-06 
3.0 4.057 0 3.0 1e-06 
0.05 4.058 0 3.0 1e-06 
3.0 4.058 0 3.0 1e-06 
0.05 4.059 0 3.0 1e-06 
3.0 4.059 0 3.0 1e-06 
0.05 4.06 0 3.0 1e-06 
3.0 4.06 0 3.0 1e-06 
0.05 4.061 0 3.0 1e-06 
3.0 4.061 0 3.0 1e-06 
0.05 4.062 0 3.0 1e-06 
3.0 4.062 0 3.0 1e-06 
0.05 4.063 0 3.0 1e-06 
3.0 4.063 0 3.0 1e-06 
0.05 4.064 0 3.0 1e-06 
3.0 4.064 0 3.0 1e-06 
0.05 4.065 0 3.0 1e-06 
3.0 4.065 0 3.0 1e-06 
0.05 4.066 0 3.0 1e-06 
3.0 4.066 0 3.0 1e-06 
0.05 4.067 0 3.0 1e-06 
3.0 4.067 0 3.0 1e-06 
0.05 4.068 0 3.0 1e-06 
3.0 4.068 0 3.0 1e-06 
0.05 4.069 0 3.0 1e-06 
3.0 4.069 0 3.0 1e-06 
0.05 4.07 0 3.0 1e-06 
3.0 4.07 0 3.0 1e-06 
0.05 4.071 0 3.0 1e-06 
3.0 4.071 0 3.0 1e-06 
0.05 4.072 0 3.0 1e-06 
3.0 4.072 0 3.0 1e-06 
0.05 4.073 0 3.0 1e-06 
3.0 4.073 0 3.0 1e-06 
0.05 4.074 0 3.0 1e-06 
3.0 4.074 0 3.0 1e-06 
0.05 4.075 0 3.0 1e-06 
3.0 4.075 0 3.0 1e-06 
0.05 4.076 0 3.0 1e-06 
3.0 4.076 0 3.0 1e-06 
0.05 4.077 0 3.0 1e-06 
3.0 4.077 0 3.0 1e-06 
0.05 4.078 0 3.0 1e-06 
3.0 4.078 0 3.0 1e-06 
0.05 4.079 0 3.0 1e-06 
3.0 4.079 0 3.0 1e-06 
0.05 4.08 0 3.0 1e-06 
3.0 4.08 0 3.0 1e-06 
0.05 4.081 0 3.0 1e-06 
3.0 4.081 0 3.0 1e-06 
0.05 4.082 0 3.0 1e-06 
3.0 4.082 0 3.0 1e-06 
0.05 4.083 0 3.0 1e-06 
3.0 4.083 0 3.0 1e-06 
0.05 4.084 0 3.0 1e-06 
3.0 4.084 0 3.0 1e-06 
0.05 4.085 0 3.0 1e-06 
3.0 4.085 0 3.0 1e-06 
0.05 4.086 0 3.0 1e-06 
3.0 4.086 0 3.0 1e-06 
0.05 4.087 0 3.0 1e-06 
3.0 4.087 0 3.0 1e-06 
0.05 4.088 0 3.0 1e-06 
3.0 4.088 0 3.0 1e-06 
0.05 4.089 0 3.0 1e-06 
3.0 4.089 0 3.0 1e-06 
0.05 4.09 0 3.0 1e-06 
3.0 4.09 0 3.0 1e-06 
0.05 4.091 0 3.0 1e-06 
3.0 4.091 0 3.0 1e-06 
0.05 4.092 0 3.0 1e-06 
3.0 4.092 0 3.0 1e-06 
0.05 4.093 0 3.0 1e-06 
3.0 4.093 0 3.0 1e-06 
0.05 4.094 0 3.0 1e-06 
3.0 4.094 0 3.0 1e-06 
0.05 4.095 0 3.0 1e-06 
3.0 4.095 0 3.0 1e-06 
0.05 4.096 0 3.0 1e-06 
3.0 4.096 0 3.0 1e-06 
0.05 4.097 0 3.0 1e-06 
3.0 4.097 0 3.0 1e-06 
0.05 4.098 0 3.0 1e-06 
3.0 4.098 0 3.0 1e-06 
0.05 4.099 0 3.0 1e-06 
3.0 4.099 0 3.0 1e-06 
0.05 4.1 0 3.0 1e-06 
3.0 4.1 0 3.0 1e-06 
0.05 4.101 0 3.0 1e-06 
3.0 4.101 0 3.0 1e-06 
0.05 4.102 0 3.0 1e-06 
3.0 4.102 0 3.0 1e-06 
0.05 4.103 0 3.0 1e-06 
3.0 4.103 0 3.0 1e-06 
0.05 4.104 0 3.0 1e-06 
3.0 4.104 0 3.0 1e-06 
0.05 4.105 0 3.0 1e-06 
3.0 4.105 0 3.0 1e-06 
0.05 4.106 0 3.0 1e-06 
3.0 4.106 0 3.0 1e-06 
0.05 4.107 0 3.0 1e-06 
3.0 4.107 0 3.0 1e-06 
0.05 4.108 0 3.0 1e-06 
3.0 4.108 0 3.0 1e-06 
0.05 4.109 0 3.0 1e-06 
3.0 4.109 0 3.0 1e-06 
0.05 4.11 0 3.0 1e-06 
3.0 4.11 0 3.0 1e-06 
0.05 4.111 0 3.0 1e-06 
3.0 4.111 0 3.0 1e-06 
0.05 4.112 0 3.0 1e-06 
3.0 4.112 0 3.0 1e-06 
0.05 4.113 0 3.0 1e-06 
3.0 4.113 0 3.0 1e-06 
0.05 4.114 0 3.0 1e-06 
3.0 4.114 0 3.0 1e-06 
0.05 4.115 0 3.0 1e-06 
3.0 4.115 0 3.0 1e-06 
0.05 4.116 0 3.0 1e-06 
3.0 4.116 0 3.0 1e-06 
0.05 4.117 0 3.0 1e-06 
3.0 4.117 0 3.0 1e-06 
0.05 4.118 0 3.0 1e-06 
3.0 4.118 0 3.0 1e-06 
0.05 4.119 0 3.0 1e-06 
3.0 4.119 0 3.0 1e-06 
0.05 4.12 0 3.0 1e-06 
3.0 4.12 0 3.0 1e-06 
0.05 4.121 0 3.0 1e-06 
3.0 4.121 0 3.0 1e-06 
0.05 4.122 0 3.0 1e-06 
3.0 4.122 0 3.0 1e-06 
0.05 4.123 0 3.0 1e-06 
3.0 4.123 0 3.0 1e-06 
0.05 4.124 0 3.0 1e-06 
3.0 4.124 0 3.0 1e-06 
0.05 4.125 0 3.0 1e-06 
3.0 4.125 0 3.0 1e-06 
0.05 4.126 0 3.0 1e-06 
3.0 4.126 0 3.0 1e-06 
0.05 4.127 0 3.0 1e-06 
3.0 4.127 0 3.0 1e-06 
0.05 4.128 0 3.0 1e-06 
3.0 4.128 0 3.0 1e-06 
0.05 4.129 0 3.0 1e-06 
3.0 4.129 0 3.0 1e-06 
0.05 4.13 0 3.0 1e-06 
3.0 4.13 0 3.0 1e-06 
0.05 4.131 0 3.0 1e-06 
3.0 4.131 0 3.0 1e-06 
0.05 4.132 0 3.0 1e-06 
3.0 4.132 0 3.0 1e-06 
0.05 4.133 0 3.0 1e-06 
3.0 4.133 0 3.0 1e-06 
0.05 4.134 0 3.0 1e-06 
3.0 4.134 0 3.0 1e-06 
0.05 4.135 0 3.0 1e-06 
3.0 4.135 0 3.0 1e-06 
0.05 4.136 0 3.0 1e-06 
3.0 4.136 0 3.0 1e-06 
0.05 4.137 0 3.0 1e-06 
3.0 4.137 0 3.0 1e-06 
0.05 4.138 0 3.0 1e-06 
3.0 4.138 0 3.0 1e-06 
0.05 4.139 0 3.0 1e-06 
3.0 4.139 0 3.0 1e-06 
0.05 4.14 0 3.0 1e-06 
3.0 4.14 0 3.0 1e-06 
0.05 4.141 0 3.0 1e-06 
3.0 4.141 0 3.0 1e-06 
0.05 4.142 0 3.0 1e-06 
3.0 4.142 0 3.0 1e-06 
0.05 4.143 0 3.0 1e-06 
3.0 4.143 0 3.0 1e-06 
0.05 4.144 0 3.0 1e-06 
3.0 4.144 0 3.0 1e-06 
0.05 4.145 0 3.0 1e-06 
3.0 4.145 0 3.0 1e-06 
0.05 4.146 0 3.0 1e-06 
3.0 4.146 0 3.0 1e-06 
0.05 4.147 0 3.0 1e-06 
3.0 4.147 0 3.0 1e-06 
0.05 4.148 0 3.0 1e-06 
3.0 4.148 0 3.0 1e-06 
0.05 4.149 0 3.0 1e-06 
3.0 4.149 0 3.0 1e-06 
0.05 4.15 0 3.0 1e-06 
3.0 4.15 0 3.0 1e-06 
0.05 4.151 0 3.0 1e-06 
3.0 4.151 0 3.0 1e-06 
0.05 4.152 0 3.0 1e-06 
3.0 4.152 0 3.0 1e-06 
0.05 4.153 0 3.0 1e-06 
3.0 4.153 0 3.0 1e-06 
0.05 4.154 0 3.0 1e-06 
3.0 4.154 0 3.0 1e-06 
0.05 4.155 0 3.0 1e-06 
3.0 4.155 0 3.0 1e-06 
0.05 4.156 0 3.0 1e-06 
3.0 4.156 0 3.0 1e-06 
0.05 4.157 0 3.0 1e-06 
3.0 4.157 0 3.0 1e-06 
0.05 4.158 0 3.0 1e-06 
3.0 4.158 0 3.0 1e-06 
0.05 4.159 0 3.0 1e-06 
3.0 4.159 0 3.0 1e-06 
0.05 4.16 0 3.0 1e-06 
3.0 4.16 0 3.0 1e-06 
0.05 4.161 0 3.0 1e-06 
3.0 4.161 0 3.0 1e-06 
0.05 4.162 0 3.0 1e-06 
3.0 4.162 0 3.0 1e-06 
0.05 4.163 0 3.0 1e-06 
3.0 4.163 0 3.0 1e-06 
0.05 4.164 0 3.0 1e-06 
3.0 4.164 0 3.0 1e-06 
0.05 4.165 0 3.0 1e-06 
3.0 4.165 0 3.0 1e-06 
0.05 4.166 0 3.0 1e-06 
3.0 4.166 0 3.0 1e-06 
0.05 4.167 0 3.0 1e-06 
3.0 4.167 0 3.0 1e-06 
0.05 4.168 0 3.0 1e-06 
3.0 4.168 0 3.0 1e-06 
0.05 4.169 0 3.0 1e-06 
3.0 4.169 0 3.0 1e-06 
0.05 4.17 0 3.0 1e-06 
3.0 4.17 0 3.0 1e-06 
0.05 4.171 0 3.0 1e-06 
3.0 4.171 0 3.0 1e-06 
0.05 4.172 0 3.0 1e-06 
3.0 4.172 0 3.0 1e-06 
0.05 4.173 0 3.0 1e-06 
3.0 4.173 0 3.0 1e-06 
0.05 4.174 0 3.0 1e-06 
3.0 4.174 0 3.0 1e-06 
0.05 4.175 0 3.0 1e-06 
3.0 4.175 0 3.0 1e-06 
0.05 4.176 0 3.0 1e-06 
3.0 4.176 0 3.0 1e-06 
0.05 4.177 0 3.0 1e-06 
3.0 4.177 0 3.0 1e-06 
0.05 4.178 0 3.0 1e-06 
3.0 4.178 0 3.0 1e-06 
0.05 4.179 0 3.0 1e-06 
3.0 4.179 0 3.0 1e-06 
0.05 4.18 0 3.0 1e-06 
3.0 4.18 0 3.0 1e-06 
0.05 4.181 0 3.0 1e-06 
3.0 4.181 0 3.0 1e-06 
0.05 4.182 0 3.0 1e-06 
3.0 4.182 0 3.0 1e-06 
0.05 4.183 0 3.0 1e-06 
3.0 4.183 0 3.0 1e-06 
0.05 4.184 0 3.0 1e-06 
3.0 4.184 0 3.0 1e-06 
0.05 4.185 0 3.0 1e-06 
3.0 4.185 0 3.0 1e-06 
0.05 4.186 0 3.0 1e-06 
3.0 4.186 0 3.0 1e-06 
0.05 4.187 0 3.0 1e-06 
3.0 4.187 0 3.0 1e-06 
0.05 4.188 0 3.0 1e-06 
3.0 4.188 0 3.0 1e-06 
0.05 4.189 0 3.0 1e-06 
3.0 4.189 0 3.0 1e-06 
0.05 4.19 0 3.0 1e-06 
3.0 4.19 0 3.0 1e-06 
0.05 4.191 0 3.0 1e-06 
3.0 4.191 0 3.0 1e-06 
0.05 4.192 0 3.0 1e-06 
3.0 4.192 0 3.0 1e-06 
0.05 4.193 0 3.0 1e-06 
3.0 4.193 0 3.0 1e-06 
0.05 4.194 0 3.0 1e-06 
3.0 4.194 0 3.0 1e-06 
0.05 4.195 0 3.0 1e-06 
3.0 4.195 0 3.0 1e-06 
0.05 4.196 0 3.0 1e-06 
3.0 4.196 0 3.0 1e-06 
0.05 4.197 0 3.0 1e-06 
3.0 4.197 0 3.0 1e-06 
0.05 4.198 0 3.0 1e-06 
3.0 4.198 0 3.0 1e-06 
0.05 4.199 0 3.0 1e-06 
3.0 4.199 0 3.0 1e-06 
0.05 4.2 0 3.0 1e-06 
3.0 4.2 0 3.0 1e-06 
0.05 4.201 0 3.0 1e-06 
3.0 4.201 0 3.0 1e-06 
0.05 4.202 0 3.0 1e-06 
3.0 4.202 0 3.0 1e-06 
0.05 4.203 0 3.0 1e-06 
3.0 4.203 0 3.0 1e-06 
0.05 4.204 0 3.0 1e-06 
3.0 4.204 0 3.0 1e-06 
0.05 4.205 0 3.0 1e-06 
3.0 4.205 0 3.0 1e-06 
0.05 4.206 0 3.0 1e-06 
3.0 4.206 0 3.0 1e-06 
0.05 4.207 0 3.0 1e-06 
3.0 4.207 0 3.0 1e-06 
0.05 4.208 0 3.0 1e-06 
3.0 4.208 0 3.0 1e-06 
0.05 4.209 0 3.0 1e-06 
3.0 4.209 0 3.0 1e-06 
0.05 4.21 0 3.0 1e-06 
3.0 4.21 0 3.0 1e-06 
0.05 4.211 0 3.0 1e-06 
3.0 4.211 0 3.0 1e-06 
0.05 4.212 0 3.0 1e-06 
3.0 4.212 0 3.0 1e-06 
0.05 4.213 0 3.0 1e-06 
3.0 4.213 0 3.0 1e-06 
0.05 4.214 0 3.0 1e-06 
3.0 4.214 0 3.0 1e-06 
0.05 4.215 0 3.0 1e-06 
3.0 4.215 0 3.0 1e-06 
0.05 4.216 0 3.0 1e-06 
3.0 4.216 0 3.0 1e-06 
0.05 4.217 0 3.0 1e-06 
3.0 4.217 0 3.0 1e-06 
0.05 4.218 0 3.0 1e-06 
3.0 4.218 0 3.0 1e-06 
0.05 4.219 0 3.0 1e-06 
3.0 4.219 0 3.0 1e-06 
0.05 4.22 0 3.0 1e-06 
3.0 4.22 0 3.0 1e-06 
0.05 4.221 0 3.0 1e-06 
3.0 4.221 0 3.0 1e-06 
0.05 4.222 0 3.0 1e-06 
3.0 4.222 0 3.0 1e-06 
0.05 4.223 0 3.0 1e-06 
3.0 4.223 0 3.0 1e-06 
0.05 4.224 0 3.0 1e-06 
3.0 4.224 0 3.0 1e-06 
0.05 4.225 0 3.0 1e-06 
3.0 4.225 0 3.0 1e-06 
0.05 4.226 0 3.0 1e-06 
3.0 4.226 0 3.0 1e-06 
0.05 4.227 0 3.0 1e-06 
3.0 4.227 0 3.0 1e-06 
0.05 4.228 0 3.0 1e-06 
3.0 4.228 0 3.0 1e-06 
0.05 4.229 0 3.0 1e-06 
3.0 4.229 0 3.0 1e-06 
0.05 4.23 0 3.0 1e-06 
3.0 4.23 0 3.0 1e-06 
0.05 4.231 0 3.0 1e-06 
3.0 4.231 0 3.0 1e-06 
0.05 4.232 0 3.0 1e-06 
3.0 4.232 0 3.0 1e-06 
0.05 4.233 0 3.0 1e-06 
3.0 4.233 0 3.0 1e-06 
0.05 4.234 0 3.0 1e-06 
3.0 4.234 0 3.0 1e-06 
0.05 4.235 0 3.0 1e-06 
3.0 4.235 0 3.0 1e-06 
0.05 4.236 0 3.0 1e-06 
3.0 4.236 0 3.0 1e-06 
0.05 4.237 0 3.0 1e-06 
3.0 4.237 0 3.0 1e-06 
0.05 4.238 0 3.0 1e-06 
3.0 4.238 0 3.0 1e-06 
0.05 4.239 0 3.0 1e-06 
3.0 4.239 0 3.0 1e-06 
0.05 4.24 0 3.0 1e-06 
3.0 4.24 0 3.0 1e-06 
0.05 4.241 0 3.0 1e-06 
3.0 4.241 0 3.0 1e-06 
0.05 4.242 0 3.0 1e-06 
3.0 4.242 0 3.0 1e-06 
0.05 4.243 0 3.0 1e-06 
3.0 4.243 0 3.0 1e-06 
0.05 4.244 0 3.0 1e-06 
3.0 4.244 0 3.0 1e-06 
0.05 4.245 0 3.0 1e-06 
3.0 4.245 0 3.0 1e-06 
0.05 4.246 0 3.0 1e-06 
3.0 4.246 0 3.0 1e-06 
0.05 4.247 0 3.0 1e-06 
3.0 4.247 0 3.0 1e-06 
0.05 4.248 0 3.0 1e-06 
3.0 4.248 0 3.0 1e-06 
0.05 4.249 0 3.0 1e-06 
3.0 4.249 0 3.0 1e-06 
0.05 4.25 0 3.0 1e-06 
3.0 4.25 0 3.0 1e-06 
0.05 4.251 0 3.0 1e-06 
3.0 4.251 0 3.0 1e-06 
0.05 4.252 0 3.0 1e-06 
3.0 4.252 0 3.0 1e-06 
0.05 4.253 0 3.0 1e-06 
3.0 4.253 0 3.0 1e-06 
0.05 4.254 0 3.0 1e-06 
3.0 4.254 0 3.0 1e-06 
0.05 4.255 0 3.0 1e-06 
3.0 4.255 0 3.0 1e-06 
0.05 4.256 0 3.0 1e-06 
3.0 4.256 0 3.0 1e-06 
0.05 4.257 0 3.0 1e-06 
3.0 4.257 0 3.0 1e-06 
0.05 4.258 0 3.0 1e-06 
3.0 4.258 0 3.0 1e-06 
0.05 4.259 0 3.0 1e-06 
3.0 4.259 0 3.0 1e-06 
0.05 4.26 0 3.0 1e-06 
3.0 4.26 0 3.0 1e-06 
0.05 4.261 0 3.0 1e-06 
3.0 4.261 0 3.0 1e-06 
0.05 4.262 0 3.0 1e-06 
3.0 4.262 0 3.0 1e-06 
0.05 4.263 0 3.0 1e-06 
3.0 4.263 0 3.0 1e-06 
0.05 4.264 0 3.0 1e-06 
3.0 4.264 0 3.0 1e-06 
0.05 4.265 0 3.0 1e-06 
3.0 4.265 0 3.0 1e-06 
0.05 4.266 0 3.0 1e-06 
3.0 4.266 0 3.0 1e-06 
0.05 4.267 0 3.0 1e-06 
3.0 4.267 0 3.0 1e-06 
0.05 4.268 0 3.0 1e-06 
3.0 4.268 0 3.0 1e-06 
0.05 4.269 0 3.0 1e-06 
3.0 4.269 0 3.0 1e-06 
0.05 4.27 0 3.0 1e-06 
3.0 4.27 0 3.0 1e-06 
0.05 4.271 0 3.0 1e-06 
3.0 4.271 0 3.0 1e-06 
0.05 4.272 0 3.0 1e-06 
3.0 4.272 0 3.0 1e-06 
0.05 4.273 0 3.0 1e-06 
3.0 4.273 0 3.0 1e-06 
0.05 4.274 0 3.0 1e-06 
3.0 4.274 0 3.0 1e-06 
0.05 4.275 0 3.0 1e-06 
3.0 4.275 0 3.0 1e-06 
0.05 4.276 0 3.0 1e-06 
3.0 4.276 0 3.0 1e-06 
0.05 4.277 0 3.0 1e-06 
3.0 4.277 0 3.0 1e-06 
0.05 4.278 0 3.0 1e-06 
3.0 4.278 0 3.0 1e-06 
0.05 4.279 0 3.0 1e-06 
3.0 4.279 0 3.0 1e-06 
0.05 4.28 0 3.0 1e-06 
3.0 4.28 0 3.0 1e-06 
0.05 4.281 0 3.0 1e-06 
3.0 4.281 0 3.0 1e-06 
0.05 4.282 0 3.0 1e-06 
3.0 4.282 0 3.0 1e-06 
0.05 4.283 0 3.0 1e-06 
3.0 4.283 0 3.0 1e-06 
0.05 4.284 0 3.0 1e-06 
3.0 4.284 0 3.0 1e-06 
0.05 4.285 0 3.0 1e-06 
3.0 4.285 0 3.0 1e-06 
0.05 4.286 0 3.0 1e-06 
3.0 4.286 0 3.0 1e-06 
0.05 4.287 0 3.0 1e-06 
3.0 4.287 0 3.0 1e-06 
0.05 4.288 0 3.0 1e-06 
3.0 4.288 0 3.0 1e-06 
0.05 4.289 0 3.0 1e-06 
3.0 4.289 0 3.0 1e-06 
0.05 4.29 0 3.0 1e-06 
3.0 4.29 0 3.0 1e-06 
0.05 4.291 0 3.0 1e-06 
3.0 4.291 0 3.0 1e-06 
0.05 4.292 0 3.0 1e-06 
3.0 4.292 0 3.0 1e-06 
0.05 4.293 0 3.0 1e-06 
3.0 4.293 0 3.0 1e-06 
0.05 4.294 0 3.0 1e-06 
3.0 4.294 0 3.0 1e-06 
0.05 4.295 0 3.0 1e-06 
3.0 4.295 0 3.0 1e-06 
0.05 4.296 0 3.0 1e-06 
3.0 4.296 0 3.0 1e-06 
0.05 4.297 0 3.0 1e-06 
3.0 4.297 0 3.0 1e-06 
0.05 4.298 0 3.0 1e-06 
3.0 4.298 0 3.0 1e-06 
0.05 4.299 0 3.0 1e-06 
3.0 4.299 0 3.0 1e-06 
0.05 4.3 0 3.0 1e-06 
3.0 4.3 0 3.0 1e-06 
0.05 4.301 0 3.0 1e-06 
3.0 4.301 0 3.0 1e-06 
0.05 4.302 0 3.0 1e-06 
3.0 4.302 0 3.0 1e-06 
0.05 4.303 0 3.0 1e-06 
3.0 4.303 0 3.0 1e-06 
0.05 4.304 0 3.0 1e-06 
3.0 4.304 0 3.0 1e-06 
0.05 4.305 0 3.0 1e-06 
3.0 4.305 0 3.0 1e-06 
0.05 4.306 0 3.0 1e-06 
3.0 4.306 0 3.0 1e-06 
0.05 4.307 0 3.0 1e-06 
3.0 4.307 0 3.0 1e-06 
0.05 4.308 0 3.0 1e-06 
3.0 4.308 0 3.0 1e-06 
0.05 4.309 0 3.0 1e-06 
3.0 4.309 0 3.0 1e-06 
0.05 4.31 0 3.0 1e-06 
3.0 4.31 0 3.0 1e-06 
0.05 4.311 0 3.0 1e-06 
3.0 4.311 0 3.0 1e-06 
0.05 4.312 0 3.0 1e-06 
3.0 4.312 0 3.0 1e-06 
0.05 4.313 0 3.0 1e-06 
3.0 4.313 0 3.0 1e-06 
0.05 4.314 0 3.0 1e-06 
3.0 4.314 0 3.0 1e-06 
0.05 4.315 0 3.0 1e-06 
3.0 4.315 0 3.0 1e-06 
0.05 4.316 0 3.0 1e-06 
3.0 4.316 0 3.0 1e-06 
0.05 4.317 0 3.0 1e-06 
3.0 4.317 0 3.0 1e-06 
0.05 4.318 0 3.0 1e-06 
3.0 4.318 0 3.0 1e-06 
0.05 4.319 0 3.0 1e-06 
3.0 4.319 0 3.0 1e-06 
0.05 4.32 0 3.0 1e-06 
3.0 4.32 0 3.0 1e-06 
0.05 4.321 0 3.0 1e-06 
3.0 4.321 0 3.0 1e-06 
0.05 4.322 0 3.0 1e-06 
3.0 4.322 0 3.0 1e-06 
0.05 4.323 0 3.0 1e-06 
3.0 4.323 0 3.0 1e-06 
0.05 4.324 0 3.0 1e-06 
3.0 4.324 0 3.0 1e-06 
0.05 4.325 0 3.0 1e-06 
3.0 4.325 0 3.0 1e-06 
0.05 4.326 0 3.0 1e-06 
3.0 4.326 0 3.0 1e-06 
0.05 4.327 0 3.0 1e-06 
3.0 4.327 0 3.0 1e-06 
0.05 4.328 0 3.0 1e-06 
3.0 4.328 0 3.0 1e-06 
0.05 4.329 0 3.0 1e-06 
3.0 4.329 0 3.0 1e-06 
0.05 4.33 0 3.0 1e-06 
3.0 4.33 0 3.0 1e-06 
0.05 4.331 0 3.0 1e-06 
3.0 4.331 0 3.0 1e-06 
0.05 4.332 0 3.0 1e-06 
3.0 4.332 0 3.0 1e-06 
0.05 4.333 0 3.0 1e-06 
3.0 4.333 0 3.0 1e-06 
0.05 4.334 0 3.0 1e-06 
3.0 4.334 0 3.0 1e-06 
0.05 4.335 0 3.0 1e-06 
3.0 4.335 0 3.0 1e-06 
0.05 4.336 0 3.0 1e-06 
3.0 4.336 0 3.0 1e-06 
0.05 4.337 0 3.0 1e-06 
3.0 4.337 0 3.0 1e-06 
0.05 4.338 0 3.0 1e-06 
3.0 4.338 0 3.0 1e-06 
0.05 4.339 0 3.0 1e-06 
3.0 4.339 0 3.0 1e-06 
0.05 4.34 0 3.0 1e-06 
3.0 4.34 0 3.0 1e-06 
0.05 4.341 0 3.0 1e-06 
3.0 4.341 0 3.0 1e-06 
0.05 4.342 0 3.0 1e-06 
3.0 4.342 0 3.0 1e-06 
0.05 4.343 0 3.0 1e-06 
3.0 4.343 0 3.0 1e-06 
0.05 4.344 0 3.0 1e-06 
3.0 4.344 0 3.0 1e-06 
0.05 4.345 0 3.0 1e-06 
3.0 4.345 0 3.0 1e-06 
0.05 4.346 0 3.0 1e-06 
3.0 4.346 0 3.0 1e-06 
0.05 4.347 0 3.0 1e-06 
3.0 4.347 0 3.0 1e-06 
0.05 4.348 0 3.0 1e-06 
3.0 4.348 0 3.0 1e-06 
0.05 4.349 0 3.0 1e-06 
3.0 4.349 0 3.0 1e-06 
0.05 4.35 0 3.0 1e-06 
3.0 4.35 0 3.0 1e-06 
0.05 4.351 0 3.0 1e-06 
3.0 4.351 0 3.0 1e-06 
0.05 4.352 0 3.0 1e-06 
3.0 4.352 0 3.0 1e-06 
0.05 4.353 0 3.0 1e-06 
3.0 4.353 0 3.0 1e-06 
0.05 4.354 0 3.0 1e-06 
3.0 4.354 0 3.0 1e-06 
0.05 4.355 0 3.0 1e-06 
3.0 4.355 0 3.0 1e-06 
0.05 4.356 0 3.0 1e-06 
3.0 4.356 0 3.0 1e-06 
0.05 4.357 0 3.0 1e-06 
3.0 4.357 0 3.0 1e-06 
0.05 4.358 0 3.0 1e-06 
3.0 4.358 0 3.0 1e-06 
0.05 4.359 0 3.0 1e-06 
3.0 4.359 0 3.0 1e-06 
0.05 4.36 0 3.0 1e-06 
3.0 4.36 0 3.0 1e-06 
0.05 4.361 0 3.0 1e-06 
3.0 4.361 0 3.0 1e-06 
0.05 4.362 0 3.0 1e-06 
3.0 4.362 0 3.0 1e-06 
0.05 4.363 0 3.0 1e-06 
3.0 4.363 0 3.0 1e-06 
0.05 4.364 0 3.0 1e-06 
3.0 4.364 0 3.0 1e-06 
0.05 4.365 0 3.0 1e-06 
3.0 4.365 0 3.0 1e-06 
0.05 4.366 0 3.0 1e-06 
3.0 4.366 0 3.0 1e-06 
0.05 4.367 0 3.0 1e-06 
3.0 4.367 0 3.0 1e-06 
0.05 4.368 0 3.0 1e-06 
3.0 4.368 0 3.0 1e-06 
0.05 4.369 0 3.0 1e-06 
3.0 4.369 0 3.0 1e-06 
0.05 4.37 0 3.0 1e-06 
3.0 4.37 0 3.0 1e-06 
0.05 4.371 0 3.0 1e-06 
3.0 4.371 0 3.0 1e-06 
0.05 4.372 0 3.0 1e-06 
3.0 4.372 0 3.0 1e-06 
0.05 4.373 0 3.0 1e-06 
3.0 4.373 0 3.0 1e-06 
0.05 4.374 0 3.0 1e-06 
3.0 4.374 0 3.0 1e-06 
0.05 4.375 0 3.0 1e-06 
3.0 4.375 0 3.0 1e-06 
0.05 4.376 0 3.0 1e-06 
3.0 4.376 0 3.0 1e-06 
0.05 4.377 0 3.0 1e-06 
3.0 4.377 0 3.0 1e-06 
0.05 4.378 0 3.0 1e-06 
3.0 4.378 0 3.0 1e-06 
0.05 4.379 0 3.0 1e-06 
3.0 4.379 0 3.0 1e-06 
0.05 4.38 0 3.0 1e-06 
3.0 4.38 0 3.0 1e-06 
0.05 4.381 0 3.0 1e-06 
3.0 4.381 0 3.0 1e-06 
0.05 4.382 0 3.0 1e-06 
3.0 4.382 0 3.0 1e-06 
0.05 4.383 0 3.0 1e-06 
3.0 4.383 0 3.0 1e-06 
0.05 4.384 0 3.0 1e-06 
3.0 4.384 0 3.0 1e-06 
0.05 4.385 0 3.0 1e-06 
3.0 4.385 0 3.0 1e-06 
0.05 4.386 0 3.0 1e-06 
3.0 4.386 0 3.0 1e-06 
0.05 4.387 0 3.0 1e-06 
3.0 4.387 0 3.0 1e-06 
0.05 4.388 0 3.0 1e-06 
3.0 4.388 0 3.0 1e-06 
0.05 4.389 0 3.0 1e-06 
3.0 4.389 0 3.0 1e-06 
0.05 4.39 0 3.0 1e-06 
3.0 4.39 0 3.0 1e-06 
0.05 4.391 0 3.0 1e-06 
3.0 4.391 0 3.0 1e-06 
0.05 4.392 0 3.0 1e-06 
3.0 4.392 0 3.0 1e-06 
0.05 4.393 0 3.0 1e-06 
3.0 4.393 0 3.0 1e-06 
0.05 4.394 0 3.0 1e-06 
3.0 4.394 0 3.0 1e-06 
0.05 4.395 0 3.0 1e-06 
3.0 4.395 0 3.0 1e-06 
0.05 4.396 0 3.0 1e-06 
3.0 4.396 0 3.0 1e-06 
0.05 4.397 0 3.0 1e-06 
3.0 4.397 0 3.0 1e-06 
0.05 4.398 0 3.0 1e-06 
3.0 4.398 0 3.0 1e-06 
0.05 4.399 0 3.0 1e-06 
3.0 4.399 0 3.0 1e-06 
0.05 4.4 0 3.0 1e-06 
3.0 4.4 0 3.0 1e-06 
0.05 4.401 0 3.0 1e-06 
3.0 4.401 0 3.0 1e-06 
0.05 4.402 0 3.0 1e-06 
3.0 4.402 0 3.0 1e-06 
0.05 4.403 0 3.0 1e-06 
3.0 4.403 0 3.0 1e-06 
0.05 4.404 0 3.0 1e-06 
3.0 4.404 0 3.0 1e-06 
0.05 4.405 0 3.0 1e-06 
3.0 4.405 0 3.0 1e-06 
0.05 4.406 0 3.0 1e-06 
3.0 4.406 0 3.0 1e-06 
0.05 4.407 0 3.0 1e-06 
3.0 4.407 0 3.0 1e-06 
0.05 4.408 0 3.0 1e-06 
3.0 4.408 0 3.0 1e-06 
0.05 4.409 0 3.0 1e-06 
3.0 4.409 0 3.0 1e-06 
0.05 4.41 0 3.0 1e-06 
3.0 4.41 0 3.0 1e-06 
0.05 4.411 0 3.0 1e-06 
3.0 4.411 0 3.0 1e-06 
0.05 4.412 0 3.0 1e-06 
3.0 4.412 0 3.0 1e-06 
0.05 4.413 0 3.0 1e-06 
3.0 4.413 0 3.0 1e-06 
0.05 4.414 0 3.0 1e-06 
3.0 4.414 0 3.0 1e-06 
0.05 4.415 0 3.0 1e-06 
3.0 4.415 0 3.0 1e-06 
0.05 4.416 0 3.0 1e-06 
3.0 4.416 0 3.0 1e-06 
0.05 4.417 0 3.0 1e-06 
3.0 4.417 0 3.0 1e-06 
0.05 4.418 0 3.0 1e-06 
3.0 4.418 0 3.0 1e-06 
0.05 4.419 0 3.0 1e-06 
3.0 4.419 0 3.0 1e-06 
0.05 4.42 0 3.0 1e-06 
3.0 4.42 0 3.0 1e-06 
0.05 4.421 0 3.0 1e-06 
3.0 4.421 0 3.0 1e-06 
0.05 4.422 0 3.0 1e-06 
3.0 4.422 0 3.0 1e-06 
0.05 4.423 0 3.0 1e-06 
3.0 4.423 0 3.0 1e-06 
0.05 4.424 0 3.0 1e-06 
3.0 4.424 0 3.0 1e-06 
0.05 4.425 0 3.0 1e-06 
3.0 4.425 0 3.0 1e-06 
0.05 4.426 0 3.0 1e-06 
3.0 4.426 0 3.0 1e-06 
0.05 4.427 0 3.0 1e-06 
3.0 4.427 0 3.0 1e-06 
0.05 4.428 0 3.0 1e-06 
3.0 4.428 0 3.0 1e-06 
0.05 4.429 0 3.0 1e-06 
3.0 4.429 0 3.0 1e-06 
0.05 4.43 0 3.0 1e-06 
3.0 4.43 0 3.0 1e-06 
0.05 4.431 0 3.0 1e-06 
3.0 4.431 0 3.0 1e-06 
0.05 4.432 0 3.0 1e-06 
3.0 4.432 0 3.0 1e-06 
0.05 4.433 0 3.0 1e-06 
3.0 4.433 0 3.0 1e-06 
0.05 4.434 0 3.0 1e-06 
3.0 4.434 0 3.0 1e-06 
0.05 4.435 0 3.0 1e-06 
3.0 4.435 0 3.0 1e-06 
0.05 4.436 0 3.0 1e-06 
3.0 4.436 0 3.0 1e-06 
0.05 4.437 0 3.0 1e-06 
3.0 4.437 0 3.0 1e-06 
0.05 4.438 0 3.0 1e-06 
3.0 4.438 0 3.0 1e-06 
0.05 4.439 0 3.0 1e-06 
3.0 4.439 0 3.0 1e-06 
0.05 4.44 0 3.0 1e-06 
3.0 4.44 0 3.0 1e-06 
0.05 4.441 0 3.0 1e-06 
3.0 4.441 0 3.0 1e-06 
0.05 4.442 0 3.0 1e-06 
3.0 4.442 0 3.0 1e-06 
0.05 4.443 0 3.0 1e-06 
3.0 4.443 0 3.0 1e-06 
0.05 4.444 0 3.0 1e-06 
3.0 4.444 0 3.0 1e-06 
0.05 4.445 0 3.0 1e-06 
3.0 4.445 0 3.0 1e-06 
0.05 4.446 0 3.0 1e-06 
3.0 4.446 0 3.0 1e-06 
0.05 4.447 0 3.0 1e-06 
3.0 4.447 0 3.0 1e-06 
0.05 4.448 0 3.0 1e-06 
3.0 4.448 0 3.0 1e-06 
0.05 4.449 0 3.0 1e-06 
3.0 4.449 0 3.0 1e-06 
0.05 4.45 0 3.0 1e-06 
3.0 4.45 0 3.0 1e-06 
0.05 4.451 0 3.0 1e-06 
3.0 4.451 0 3.0 1e-06 
0.05 4.452 0 3.0 1e-06 
3.0 4.452 0 3.0 1e-06 
0.05 4.453 0 3.0 1e-06 
3.0 4.453 0 3.0 1e-06 
0.05 4.454 0 3.0 1e-06 
3.0 4.454 0 3.0 1e-06 
0.05 4.455 0 3.0 1e-06 
3.0 4.455 0 3.0 1e-06 
0.05 4.456 0 3.0 1e-06 
3.0 4.456 0 3.0 1e-06 
0.05 4.457 0 3.0 1e-06 
3.0 4.457 0 3.0 1e-06 
0.05 4.458 0 3.0 1e-06 
3.0 4.458 0 3.0 1e-06 
0.05 4.459 0 3.0 1e-06 
3.0 4.459 0 3.0 1e-06 
0.05 4.46 0 3.0 1e-06 
3.0 4.46 0 3.0 1e-06 
0.05 4.461 0 3.0 1e-06 
3.0 4.461 0 3.0 1e-06 
0.05 4.462 0 3.0 1e-06 
3.0 4.462 0 3.0 1e-06 
0.05 4.463 0 3.0 1e-06 
3.0 4.463 0 3.0 1e-06 
0.05 4.464 0 3.0 1e-06 
3.0 4.464 0 3.0 1e-06 
0.05 4.465 0 3.0 1e-06 
3.0 4.465 0 3.0 1e-06 
0.05 4.466 0 3.0 1e-06 
3.0 4.466 0 3.0 1e-06 
0.05 4.467 0 3.0 1e-06 
3.0 4.467 0 3.0 1e-06 
0.05 4.468 0 3.0 1e-06 
3.0 4.468 0 3.0 1e-06 
0.05 4.469 0 3.0 1e-06 
3.0 4.469 0 3.0 1e-06 
0.05 4.47 0 3.0 1e-06 
3.0 4.47 0 3.0 1e-06 
0.05 4.471 0 3.0 1e-06 
3.0 4.471 0 3.0 1e-06 
0.05 4.472 0 3.0 1e-06 
3.0 4.472 0 3.0 1e-06 
0.05 4.473 0 3.0 1e-06 
3.0 4.473 0 3.0 1e-06 
0.05 4.474 0 3.0 1e-06 
3.0 4.474 0 3.0 1e-06 
0.05 4.475 0 3.0 1e-06 
3.0 4.475 0 3.0 1e-06 
0.05 4.476 0 3.0 1e-06 
3.0 4.476 0 3.0 1e-06 
0.05 4.477 0 3.0 1e-06 
3.0 4.477 0 3.0 1e-06 
0.05 4.478 0 3.0 1e-06 
3.0 4.478 0 3.0 1e-06 
0.05 4.479 0 3.0 1e-06 
3.0 4.479 0 3.0 1e-06 
0.05 4.48 0 3.0 1e-06 
3.0 4.48 0 3.0 1e-06 
0.05 4.481 0 3.0 1e-06 
3.0 4.481 0 3.0 1e-06 
0.05 4.482 0 3.0 1e-06 
3.0 4.482 0 3.0 1e-06 
0.05 4.483 0 3.0 1e-06 
3.0 4.483 0 3.0 1e-06 
0.05 4.484 0 3.0 1e-06 
3.0 4.484 0 3.0 1e-06 
0.05 4.485 0 3.0 1e-06 
3.0 4.485 0 3.0 1e-06 
0.05 4.486 0 3.0 1e-06 
3.0 4.486 0 3.0 1e-06 
0.05 4.487 0 3.0 1e-06 
3.0 4.487 0 3.0 1e-06 
0.05 4.488 0 3.0 1e-06 
3.0 4.488 0 3.0 1e-06 
0.05 4.489 0 3.0 1e-06 
3.0 4.489 0 3.0 1e-06 
0.05 4.49 0 3.0 1e-06 
3.0 4.49 0 3.0 1e-06 
0.05 4.491 0 3.0 1e-06 
3.0 4.491 0 3.0 1e-06 
0.05 4.492 0 3.0 1e-06 
3.0 4.492 0 3.0 1e-06 
0.05 4.493 0 3.0 1e-06 
3.0 4.493 0 3.0 1e-06 
0.05 4.494 0 3.0 1e-06 
3.0 4.494 0 3.0 1e-06 
0.05 4.495 0 3.0 1e-06 
3.0 4.495 0 3.0 1e-06 
0.05 4.496 0 3.0 1e-06 
3.0 4.496 0 3.0 1e-06 
0.05 4.497 0 3.0 1e-06 
3.0 4.497 0 3.0 1e-06 
0.05 4.498 0 3.0 1e-06 
3.0 4.498 0 3.0 1e-06 
0.05 4.499 0 3.0 1e-06 
3.0 4.499 0 3.0 1e-06 
0.05 4.5 0 3.0 1e-06 
3.0 4.5 0 3.0 1e-06 
0.05 4.501 0 3.0 1e-06 
3.0 4.501 0 3.0 1e-06 
0.05 4.502 0 3.0 1e-06 
3.0 4.502 0 3.0 1e-06 
0.05 4.503 0 3.0 1e-06 
3.0 4.503 0 3.0 1e-06 
0.05 4.504 0 3.0 1e-06 
3.0 4.504 0 3.0 1e-06 
0.05 4.505 0 3.0 1e-06 
3.0 4.505 0 3.0 1e-06 
0.05 4.506 0 3.0 1e-06 
3.0 4.506 0 3.0 1e-06 
0.05 4.507 0 3.0 1e-06 
3.0 4.507 0 3.0 1e-06 
0.05 4.508 0 3.0 1e-06 
3.0 4.508 0 3.0 1e-06 
0.05 4.509 0 3.0 1e-06 
3.0 4.509 0 3.0 1e-06 
0.05 4.51 0 3.0 1e-06 
3.0 4.51 0 3.0 1e-06 
0.05 4.511 0 3.0 1e-06 
3.0 4.511 0 3.0 1e-06 
0.05 4.512 0 3.0 1e-06 
3.0 4.512 0 3.0 1e-06 
0.05 4.513 0 3.0 1e-06 
3.0 4.513 0 3.0 1e-06 
0.05 4.514 0 3.0 1e-06 
3.0 4.514 0 3.0 1e-06 
0.05 4.515 0 3.0 1e-06 
3.0 4.515 0 3.0 1e-06 
0.05 4.516 0 3.0 1e-06 
3.0 4.516 0 3.0 1e-06 
0.05 4.517 0 3.0 1e-06 
3.0 4.517 0 3.0 1e-06 
0.05 4.518 0 3.0 1e-06 
3.0 4.518 0 3.0 1e-06 
0.05 4.519 0 3.0 1e-06 
3.0 4.519 0 3.0 1e-06 
0.05 4.52 0 3.0 1e-06 
3.0 4.52 0 3.0 1e-06 
0.05 4.521 0 3.0 1e-06 
3.0 4.521 0 3.0 1e-06 
0.05 4.522 0 3.0 1e-06 
3.0 4.522 0 3.0 1e-06 
0.05 4.523 0 3.0 1e-06 
3.0 4.523 0 3.0 1e-06 
0.05 4.524 0 3.0 1e-06 
3.0 4.524 0 3.0 1e-06 
0.05 4.525 0 3.0 1e-06 
3.0 4.525 0 3.0 1e-06 
0.05 4.526 0 3.0 1e-06 
3.0 4.526 0 3.0 1e-06 
0.05 4.527 0 3.0 1e-06 
3.0 4.527 0 3.0 1e-06 
0.05 4.528 0 3.0 1e-06 
3.0 4.528 0 3.0 1e-06 
0.05 4.529 0 3.0 1e-06 
3.0 4.529 0 3.0 1e-06 
0.05 4.53 0 3.0 1e-06 
3.0 4.53 0 3.0 1e-06 
0.05 4.531 0 3.0 1e-06 
3.0 4.531 0 3.0 1e-06 
0.05 4.532 0 3.0 1e-06 
3.0 4.532 0 3.0 1e-06 
0.05 4.533 0 3.0 1e-06 
3.0 4.533 0 3.0 1e-06 
0.05 4.534 0 3.0 1e-06 
3.0 4.534 0 3.0 1e-06 
0.05 4.535 0 3.0 1e-06 
3.0 4.535 0 3.0 1e-06 
0.05 4.536 0 3.0 1e-06 
3.0 4.536 0 3.0 1e-06 
0.05 4.537 0 3.0 1e-06 
3.0 4.537 0 3.0 1e-06 
0.05 4.538 0 3.0 1e-06 
3.0 4.538 0 3.0 1e-06 
0.05 4.539 0 3.0 1e-06 
3.0 4.539 0 3.0 1e-06 
0.05 4.54 0 3.0 1e-06 
3.0 4.54 0 3.0 1e-06 
0.05 4.541 0 3.0 1e-06 
3.0 4.541 0 3.0 1e-06 
0.05 4.542 0 3.0 1e-06 
3.0 4.542 0 3.0 1e-06 
0.05 4.543 0 3.0 1e-06 
3.0 4.543 0 3.0 1e-06 
0.05 4.544 0 3.0 1e-06 
3.0 4.544 0 3.0 1e-06 
0.05 4.545 0 3.0 1e-06 
3.0 4.545 0 3.0 1e-06 
0.05 4.546 0 3.0 1e-06 
3.0 4.546 0 3.0 1e-06 
0.05 4.547 0 3.0 1e-06 
3.0 4.547 0 3.0 1e-06 
0.05 4.548 0 3.0 1e-06 
3.0 4.548 0 3.0 1e-06 
0.05 4.549 0 3.0 1e-06 
3.0 4.549 0 3.0 1e-06 
0.05 4.55 0 3.0 1e-06 
3.0 4.55 0 3.0 1e-06 
0.05 4.551 0 3.0 1e-06 
3.0 4.551 0 3.0 1e-06 
0.05 4.552 0 3.0 1e-06 
3.0 4.552 0 3.0 1e-06 
0.05 4.553 0 3.0 1e-06 
3.0 4.553 0 3.0 1e-06 
0.05 4.554 0 3.0 1e-06 
3.0 4.554 0 3.0 1e-06 
0.05 4.555 0 3.0 1e-06 
3.0 4.555 0 3.0 1e-06 
0.05 4.556 0 3.0 1e-06 
3.0 4.556 0 3.0 1e-06 
0.05 4.557 0 3.0 1e-06 
3.0 4.557 0 3.0 1e-06 
0.05 4.558 0 3.0 1e-06 
3.0 4.558 0 3.0 1e-06 
0.05 4.559 0 3.0 1e-06 
3.0 4.559 0 3.0 1e-06 
0.05 4.56 0 3.0 1e-06 
3.0 4.56 0 3.0 1e-06 
0.05 4.561 0 3.0 1e-06 
3.0 4.561 0 3.0 1e-06 
0.05 4.562 0 3.0 1e-06 
3.0 4.562 0 3.0 1e-06 
0.05 4.563 0 3.0 1e-06 
3.0 4.563 0 3.0 1e-06 
0.05 4.564 0 3.0 1e-06 
3.0 4.564 0 3.0 1e-06 
0.05 4.565 0 3.0 1e-06 
3.0 4.565 0 3.0 1e-06 
0.05 4.566 0 3.0 1e-06 
3.0 4.566 0 3.0 1e-06 
0.05 4.567 0 3.0 1e-06 
3.0 4.567 0 3.0 1e-06 
0.05 4.568 0 3.0 1e-06 
3.0 4.568 0 3.0 1e-06 
0.05 4.569 0 3.0 1e-06 
3.0 4.569 0 3.0 1e-06 
0.05 4.57 0 3.0 1e-06 
3.0 4.57 0 3.0 1e-06 
0.05 4.571 0 3.0 1e-06 
3.0 4.571 0 3.0 1e-06 
0.05 4.572 0 3.0 1e-06 
3.0 4.572 0 3.0 1e-06 
0.05 4.573 0 3.0 1e-06 
3.0 4.573 0 3.0 1e-06 
0.05 4.574 0 3.0 1e-06 
3.0 4.574 0 3.0 1e-06 
0.05 4.575 0 3.0 1e-06 
3.0 4.575 0 3.0 1e-06 
0.05 4.576 0 3.0 1e-06 
3.0 4.576 0 3.0 1e-06 
0.05 4.577 0 3.0 1e-06 
3.0 4.577 0 3.0 1e-06 
0.05 4.578 0 3.0 1e-06 
3.0 4.578 0 3.0 1e-06 
0.05 4.579 0 3.0 1e-06 
3.0 4.579 0 3.0 1e-06 
0.05 4.58 0 3.0 1e-06 
3.0 4.58 0 3.0 1e-06 
0.05 4.581 0 3.0 1e-06 
3.0 4.581 0 3.0 1e-06 
0.05 4.582 0 3.0 1e-06 
3.0 4.582 0 3.0 1e-06 
0.05 4.583 0 3.0 1e-06 
3.0 4.583 0 3.0 1e-06 
0.05 4.584 0 3.0 1e-06 
3.0 4.584 0 3.0 1e-06 
0.05 4.585 0 3.0 1e-06 
3.0 4.585 0 3.0 1e-06 
0.05 4.586 0 3.0 1e-06 
3.0 4.586 0 3.0 1e-06 
0.05 4.587 0 3.0 1e-06 
3.0 4.587 0 3.0 1e-06 
0.05 4.588 0 3.0 1e-06 
3.0 4.588 0 3.0 1e-06 
0.05 4.589 0 3.0 1e-06 
3.0 4.589 0 3.0 1e-06 
0.05 4.59 0 3.0 1e-06 
3.0 4.59 0 3.0 1e-06 
0.05 4.591 0 3.0 1e-06 
3.0 4.591 0 3.0 1e-06 
0.05 4.592 0 3.0 1e-06 
3.0 4.592 0 3.0 1e-06 
0.05 4.593 0 3.0 1e-06 
3.0 4.593 0 3.0 1e-06 
0.05 4.594 0 3.0 1e-06 
3.0 4.594 0 3.0 1e-06 
0.05 4.595 0 3.0 1e-06 
3.0 4.595 0 3.0 1e-06 
0.05 4.596 0 3.0 1e-06 
3.0 4.596 0 3.0 1e-06 
0.05 4.597 0 3.0 1e-06 
3.0 4.597 0 3.0 1e-06 
0.05 4.598 0 3.0 1e-06 
3.0 4.598 0 3.0 1e-06 
0.05 4.599 0 3.0 1e-06 
3.0 4.599 0 3.0 1e-06 
0.05 4.6 0 3.0 1e-06 
3.0 4.6 0 3.0 1e-06 
0.05 4.601 0 3.0 1e-06 
3.0 4.601 0 3.0 1e-06 
0.05 4.602 0 3.0 1e-06 
3.0 4.602 0 3.0 1e-06 
0.05 4.603 0 3.0 1e-06 
3.0 4.603 0 3.0 1e-06 
0.05 4.604 0 3.0 1e-06 
3.0 4.604 0 3.0 1e-06 
0.05 4.605 0 3.0 1e-06 
3.0 4.605 0 3.0 1e-06 
0.05 4.606 0 3.0 1e-06 
3.0 4.606 0 3.0 1e-06 
0.05 4.607 0 3.0 1e-06 
3.0 4.607 0 3.0 1e-06 
0.05 4.608 0 3.0 1e-06 
3.0 4.608 0 3.0 1e-06 
0.05 4.609 0 3.0 1e-06 
3.0 4.609 0 3.0 1e-06 
0.05 4.61 0 3.0 1e-06 
3.0 4.61 0 3.0 1e-06 
0.05 4.611 0 3.0 1e-06 
3.0 4.611 0 3.0 1e-06 
0.05 4.612 0 3.0 1e-06 
3.0 4.612 0 3.0 1e-06 
0.05 4.613 0 3.0 1e-06 
3.0 4.613 0 3.0 1e-06 
0.05 4.614 0 3.0 1e-06 
3.0 4.614 0 3.0 1e-06 
0.05 4.615 0 3.0 1e-06 
3.0 4.615 0 3.0 1e-06 
0.05 4.616 0 3.0 1e-06 
3.0 4.616 0 3.0 1e-06 
0.05 4.617 0 3.0 1e-06 
3.0 4.617 0 3.0 1e-06 
0.05 4.618 0 3.0 1e-06 
3.0 4.618 0 3.0 1e-06 
0.05 4.619 0 3.0 1e-06 
3.0 4.619 0 3.0 1e-06 
0.05 4.62 0 3.0 1e-06 
3.0 4.62 0 3.0 1e-06 
0.05 4.621 0 3.0 1e-06 
3.0 4.621 0 3.0 1e-06 
0.05 4.622 0 3.0 1e-06 
3.0 4.622 0 3.0 1e-06 
0.05 4.623 0 3.0 1e-06 
3.0 4.623 0 3.0 1e-06 
0.05 4.624 0 3.0 1e-06 
3.0 4.624 0 3.0 1e-06 
0.05 4.625 0 3.0 1e-06 
3.0 4.625 0 3.0 1e-06 
0.05 4.626 0 3.0 1e-06 
3.0 4.626 0 3.0 1e-06 
0.05 4.627 0 3.0 1e-06 
3.0 4.627 0 3.0 1e-06 
0.05 4.628 0 3.0 1e-06 
3.0 4.628 0 3.0 1e-06 
0.05 4.629 0 3.0 1e-06 
3.0 4.629 0 3.0 1e-06 
0.05 4.63 0 3.0 1e-06 
3.0 4.63 0 3.0 1e-06 
0.05 4.631 0 3.0 1e-06 
3.0 4.631 0 3.0 1e-06 
0.05 4.632 0 3.0 1e-06 
3.0 4.632 0 3.0 1e-06 
0.05 4.633 0 3.0 1e-06 
3.0 4.633 0 3.0 1e-06 
0.05 4.634 0 3.0 1e-06 
3.0 4.634 0 3.0 1e-06 
0.05 4.635 0 3.0 1e-06 
3.0 4.635 0 3.0 1e-06 
0.05 4.636 0 3.0 1e-06 
3.0 4.636 0 3.0 1e-06 
0.05 4.637 0 3.0 1e-06 
3.0 4.637 0 3.0 1e-06 
0.05 4.638 0 3.0 1e-06 
3.0 4.638 0 3.0 1e-06 
0.05 4.639 0 3.0 1e-06 
3.0 4.639 0 3.0 1e-06 
0.05 4.64 0 3.0 1e-06 
3.0 4.64 0 3.0 1e-06 
0.05 4.641 0 3.0 1e-06 
3.0 4.641 0 3.0 1e-06 
0.05 4.642 0 3.0 1e-06 
3.0 4.642 0 3.0 1e-06 
0.05 4.643 0 3.0 1e-06 
3.0 4.643 0 3.0 1e-06 
0.05 4.644 0 3.0 1e-06 
3.0 4.644 0 3.0 1e-06 
0.05 4.645 0 3.0 1e-06 
3.0 4.645 0 3.0 1e-06 
0.05 4.646 0 3.0 1e-06 
3.0 4.646 0 3.0 1e-06 
0.05 4.647 0 3.0 1e-06 
3.0 4.647 0 3.0 1e-06 
0.05 4.648 0 3.0 1e-06 
3.0 4.648 0 3.0 1e-06 
0.05 4.649 0 3.0 1e-06 
3.0 4.649 0 3.0 1e-06 
0.05 4.65 0 3.0 1e-06 
3.0 4.65 0 3.0 1e-06 
0.05 4.651 0 3.0 1e-06 
3.0 4.651 0 3.0 1e-06 
0.05 4.652 0 3.0 1e-06 
3.0 4.652 0 3.0 1e-06 
0.05 4.653 0 3.0 1e-06 
3.0 4.653 0 3.0 1e-06 
0.05 4.654 0 3.0 1e-06 
3.0 4.654 0 3.0 1e-06 
0.05 4.655 0 3.0 1e-06 
3.0 4.655 0 3.0 1e-06 
0.05 4.656 0 3.0 1e-06 
3.0 4.656 0 3.0 1e-06 
0.05 4.657 0 3.0 1e-06 
3.0 4.657 0 3.0 1e-06 
0.05 4.658 0 3.0 1e-06 
3.0 4.658 0 3.0 1e-06 
0.05 4.659 0 3.0 1e-06 
3.0 4.659 0 3.0 1e-06 
0.05 4.66 0 3.0 1e-06 
3.0 4.66 0 3.0 1e-06 
0.05 4.661 0 3.0 1e-06 
3.0 4.661 0 3.0 1e-06 
0.05 4.662 0 3.0 1e-06 
3.0 4.662 0 3.0 1e-06 
0.05 4.663 0 3.0 1e-06 
3.0 4.663 0 3.0 1e-06 
0.05 4.664 0 3.0 1e-06 
3.0 4.664 0 3.0 1e-06 
0.05 4.665 0 3.0 1e-06 
3.0 4.665 0 3.0 1e-06 
0.05 4.666 0 3.0 1e-06 
3.0 4.666 0 3.0 1e-06 
0.05 4.667 0 3.0 1e-06 
3.0 4.667 0 3.0 1e-06 
0.05 4.668 0 3.0 1e-06 
3.0 4.668 0 3.0 1e-06 
0.05 4.669 0 3.0 1e-06 
3.0 4.669 0 3.0 1e-06 
0.05 4.67 0 3.0 1e-06 
3.0 4.67 0 3.0 1e-06 
0.05 4.671 0 3.0 1e-06 
3.0 4.671 0 3.0 1e-06 
0.05 4.672 0 3.0 1e-06 
3.0 4.672 0 3.0 1e-06 
0.05 4.673 0 3.0 1e-06 
3.0 4.673 0 3.0 1e-06 
0.05 4.674 0 3.0 1e-06 
3.0 4.674 0 3.0 1e-06 
0.05 4.675 0 3.0 1e-06 
3.0 4.675 0 3.0 1e-06 
0.05 4.676 0 3.0 1e-06 
3.0 4.676 0 3.0 1e-06 
0.05 4.677 0 3.0 1e-06 
3.0 4.677 0 3.0 1e-06 
0.05 4.678 0 3.0 1e-06 
3.0 4.678 0 3.0 1e-06 
0.05 4.679 0 3.0 1e-06 
3.0 4.679 0 3.0 1e-06 
0.05 4.68 0 3.0 1e-06 
3.0 4.68 0 3.0 1e-06 
0.05 4.681 0 3.0 1e-06 
3.0 4.681 0 3.0 1e-06 
0.05 4.682 0 3.0 1e-06 
3.0 4.682 0 3.0 1e-06 
0.05 4.683 0 3.0 1e-06 
3.0 4.683 0 3.0 1e-06 
0.05 4.684 0 3.0 1e-06 
3.0 4.684 0 3.0 1e-06 
0.05 4.685 0 3.0 1e-06 
3.0 4.685 0 3.0 1e-06 
0.05 4.686 0 3.0 1e-06 
3.0 4.686 0 3.0 1e-06 
0.05 4.687 0 3.0 1e-06 
3.0 4.687 0 3.0 1e-06 
0.05 4.688 0 3.0 1e-06 
3.0 4.688 0 3.0 1e-06 
0.05 4.689 0 3.0 1e-06 
3.0 4.689 0 3.0 1e-06 
0.05 4.69 0 3.0 1e-06 
3.0 4.69 0 3.0 1e-06 
0.05 4.691 0 3.0 1e-06 
3.0 4.691 0 3.0 1e-06 
0.05 4.692 0 3.0 1e-06 
3.0 4.692 0 3.0 1e-06 
0.05 4.693 0 3.0 1e-06 
3.0 4.693 0 3.0 1e-06 
0.05 4.694 0 3.0 1e-06 
3.0 4.694 0 3.0 1e-06 
0.05 4.695 0 3.0 1e-06 
3.0 4.695 0 3.0 1e-06 
0.05 4.696 0 3.0 1e-06 
3.0 4.696 0 3.0 1e-06 
0.05 4.697 0 3.0 1e-06 
3.0 4.697 0 3.0 1e-06 
0.05 4.698 0 3.0 1e-06 
3.0 4.698 0 3.0 1e-06 
0.05 4.699 0 3.0 1e-06 
3.0 4.699 0 3.0 1e-06 
0.05 4.7 0 3.0 1e-06 
3.0 4.7 0 3.0 1e-06 
0.05 4.701 0 3.0 1e-06 
3.0 4.701 0 3.0 1e-06 
0.05 4.702 0 3.0 1e-06 
3.0 4.702 0 3.0 1e-06 
0.05 4.703 0 3.0 1e-06 
3.0 4.703 0 3.0 1e-06 
0.05 4.704 0 3.0 1e-06 
3.0 4.704 0 3.0 1e-06 
0.05 4.705 0 3.0 1e-06 
3.0 4.705 0 3.0 1e-06 
0.05 4.706 0 3.0 1e-06 
3.0 4.706 0 3.0 1e-06 
0.05 4.707 0 3.0 1e-06 
3.0 4.707 0 3.0 1e-06 
0.05 4.708 0 3.0 1e-06 
3.0 4.708 0 3.0 1e-06 
0.05 4.709 0 3.0 1e-06 
3.0 4.709 0 3.0 1e-06 
0.05 4.71 0 3.0 1e-06 
3.0 4.71 0 3.0 1e-06 
0.05 4.711 0 3.0 1e-06 
3.0 4.711 0 3.0 1e-06 
0.05 4.712 0 3.0 1e-06 
3.0 4.712 0 3.0 1e-06 
0.05 4.713 0 3.0 1e-06 
3.0 4.713 0 3.0 1e-06 
0.05 4.714 0 3.0 1e-06 
3.0 4.714 0 3.0 1e-06 
0.05 4.715 0 3.0 1e-06 
3.0 4.715 0 3.0 1e-06 
0.05 4.716 0 3.0 1e-06 
3.0 4.716 0 3.0 1e-06 
0.05 4.717 0 3.0 1e-06 
3.0 4.717 0 3.0 1e-06 
0.05 4.718 0 3.0 1e-06 
3.0 4.718 0 3.0 1e-06 
0.05 4.719 0 3.0 1e-06 
3.0 4.719 0 3.0 1e-06 
0.05 4.72 0 3.0 1e-06 
3.0 4.72 0 3.0 1e-06 
0.05 4.721 0 3.0 1e-06 
3.0 4.721 0 3.0 1e-06 
0.05 4.722 0 3.0 1e-06 
3.0 4.722 0 3.0 1e-06 
0.05 4.723 0 3.0 1e-06 
3.0 4.723 0 3.0 1e-06 
0.05 4.724 0 3.0 1e-06 
3.0 4.724 0 3.0 1e-06 
0.05 4.725 0 3.0 1e-06 
3.0 4.725 0 3.0 1e-06 
0.05 4.726 0 3.0 1e-06 
3.0 4.726 0 3.0 1e-06 
0.05 4.727 0 3.0 1e-06 
3.0 4.727 0 3.0 1e-06 
0.05 4.728 0 3.0 1e-06 
3.0 4.728 0 3.0 1e-06 
0.05 4.729 0 3.0 1e-06 
3.0 4.729 0 3.0 1e-06 
0.05 4.73 0 3.0 1e-06 
3.0 4.73 0 3.0 1e-06 
0.05 4.731 0 3.0 1e-06 
3.0 4.731 0 3.0 1e-06 
0.05 4.732 0 3.0 1e-06 
3.0 4.732 0 3.0 1e-06 
0.05 4.733 0 3.0 1e-06 
3.0 4.733 0 3.0 1e-06 
0.05 4.734 0 3.0 1e-06 
3.0 4.734 0 3.0 1e-06 
0.05 4.735 0 3.0 1e-06 
3.0 4.735 0 3.0 1e-06 
0.05 4.736 0 3.0 1e-06 
3.0 4.736 0 3.0 1e-06 
0.05 4.737 0 3.0 1e-06 
3.0 4.737 0 3.0 1e-06 
0.05 4.738 0 3.0 1e-06 
3.0 4.738 0 3.0 1e-06 
0.05 4.739 0 3.0 1e-06 
3.0 4.739 0 3.0 1e-06 
0.05 4.74 0 3.0 1e-06 
3.0 4.74 0 3.0 1e-06 
0.05 4.741 0 3.0 1e-06 
3.0 4.741 0 3.0 1e-06 
0.05 4.742 0 3.0 1e-06 
3.0 4.742 0 3.0 1e-06 
0.05 4.743 0 3.0 1e-06 
3.0 4.743 0 3.0 1e-06 
0.05 4.744 0 3.0 1e-06 
3.0 4.744 0 3.0 1e-06 
0.05 4.745 0 3.0 1e-06 
3.0 4.745 0 3.0 1e-06 
0.05 4.746 0 3.0 1e-06 
3.0 4.746 0 3.0 1e-06 
0.05 4.747 0 3.0 1e-06 
3.0 4.747 0 3.0 1e-06 
0.05 4.748 0 3.0 1e-06 
3.0 4.748 0 3.0 1e-06 
0.05 4.749 0 3.0 1e-06 
3.0 4.749 0 3.0 1e-06 
0.05 4.75 0 3.0 1e-06 
3.0 4.75 0 3.0 1e-06 
0.05 4.751 0 3.0 1e-06 
3.0 4.751 0 3.0 1e-06 
0.05 4.752 0 3.0 1e-06 
3.0 4.752 0 3.0 1e-06 
0.05 4.753 0 3.0 1e-06 
3.0 4.753 0 3.0 1e-06 
0.05 4.754 0 3.0 1e-06 
3.0 4.754 0 3.0 1e-06 
0.05 4.755 0 3.0 1e-06 
3.0 4.755 0 3.0 1e-06 
0.05 4.756 0 3.0 1e-06 
3.0 4.756 0 3.0 1e-06 
0.05 4.757 0 3.0 1e-06 
3.0 4.757 0 3.0 1e-06 
0.05 4.758 0 3.0 1e-06 
3.0 4.758 0 3.0 1e-06 
0.05 4.759 0 3.0 1e-06 
3.0 4.759 0 3.0 1e-06 
0.05 4.76 0 3.0 1e-06 
3.0 4.76 0 3.0 1e-06 
0.05 4.761 0 3.0 1e-06 
3.0 4.761 0 3.0 1e-06 
0.05 4.762 0 3.0 1e-06 
3.0 4.762 0 3.0 1e-06 
0.05 4.763 0 3.0 1e-06 
3.0 4.763 0 3.0 1e-06 
0.05 4.764 0 3.0 1e-06 
3.0 4.764 0 3.0 1e-06 
0.05 4.765 0 3.0 1e-06 
3.0 4.765 0 3.0 1e-06 
0.05 4.766 0 3.0 1e-06 
3.0 4.766 0 3.0 1e-06 
0.05 4.767 0 3.0 1e-06 
3.0 4.767 0 3.0 1e-06 
0.05 4.768 0 3.0 1e-06 
3.0 4.768 0 3.0 1e-06 
0.05 4.769 0 3.0 1e-06 
3.0 4.769 0 3.0 1e-06 
0.05 4.77 0 3.0 1e-06 
3.0 4.77 0 3.0 1e-06 
0.05 4.771 0 3.0 1e-06 
3.0 4.771 0 3.0 1e-06 
0.05 4.772 0 3.0 1e-06 
3.0 4.772 0 3.0 1e-06 
0.05 4.773 0 3.0 1e-06 
3.0 4.773 0 3.0 1e-06 
0.05 4.774 0 3.0 1e-06 
3.0 4.774 0 3.0 1e-06 
0.05 4.775 0 3.0 1e-06 
3.0 4.775 0 3.0 1e-06 
0.05 4.776 0 3.0 1e-06 
3.0 4.776 0 3.0 1e-06 
0.05 4.777 0 3.0 1e-06 
3.0 4.777 0 3.0 1e-06 
0.05 4.778 0 3.0 1e-06 
3.0 4.778 0 3.0 1e-06 
0.05 4.779 0 3.0 1e-06 
3.0 4.779 0 3.0 1e-06 
0.05 4.78 0 3.0 1e-06 
3.0 4.78 0 3.0 1e-06 
0.05 4.781 0 3.0 1e-06 
3.0 4.781 0 3.0 1e-06 
0.05 4.782 0 3.0 1e-06 
3.0 4.782 0 3.0 1e-06 
0.05 4.783 0 3.0 1e-06 
3.0 4.783 0 3.0 1e-06 
0.05 4.784 0 3.0 1e-06 
3.0 4.784 0 3.0 1e-06 
0.05 4.785 0 3.0 1e-06 
3.0 4.785 0 3.0 1e-06 
0.05 4.786 0 3.0 1e-06 
3.0 4.786 0 3.0 1e-06 
0.05 4.787 0 3.0 1e-06 
3.0 4.787 0 3.0 1e-06 
0.05 4.788 0 3.0 1e-06 
3.0 4.788 0 3.0 1e-06 
0.05 4.789 0 3.0 1e-06 
3.0 4.789 0 3.0 1e-06 
0.05 4.79 0 3.0 1e-06 
3.0 4.79 0 3.0 1e-06 
0.05 4.791 0 3.0 1e-06 
3.0 4.791 0 3.0 1e-06 
0.05 4.792 0 3.0 1e-06 
3.0 4.792 0 3.0 1e-06 
0.05 4.793 0 3.0 1e-06 
3.0 4.793 0 3.0 1e-06 
0.05 4.794 0 3.0 1e-06 
3.0 4.794 0 3.0 1e-06 
0.05 4.795 0 3.0 1e-06 
3.0 4.795 0 3.0 1e-06 
0.05 4.796 0 3.0 1e-06 
3.0 4.796 0 3.0 1e-06 
0.05 4.797 0 3.0 1e-06 
3.0 4.797 0 3.0 1e-06 
0.05 4.798 0 3.0 1e-06 
3.0 4.798 0 3.0 1e-06 
0.05 4.799 0 3.0 1e-06 
3.0 4.799 0 3.0 1e-06 
0.05 4.8 0 3.0 1e-06 
3.0 4.8 0 3.0 1e-06 
0.05 4.801 0 3.0 1e-06 
3.0 4.801 0 3.0 1e-06 
0.05 4.802 0 3.0 1e-06 
3.0 4.802 0 3.0 1e-06 
0.05 4.803 0 3.0 1e-06 
3.0 4.803 0 3.0 1e-06 
0.05 4.804 0 3.0 1e-06 
3.0 4.804 0 3.0 1e-06 
0.05 4.805 0 3.0 1e-06 
3.0 4.805 0 3.0 1e-06 
0.05 4.806 0 3.0 1e-06 
3.0 4.806 0 3.0 1e-06 
0.05 4.807 0 3.0 1e-06 
3.0 4.807 0 3.0 1e-06 
0.05 4.808 0 3.0 1e-06 
3.0 4.808 0 3.0 1e-06 
0.05 4.809 0 3.0 1e-06 
3.0 4.809 0 3.0 1e-06 
0.05 4.81 0 3.0 1e-06 
3.0 4.81 0 3.0 1e-06 
0.05 4.811 0 3.0 1e-06 
3.0 4.811 0 3.0 1e-06 
0.05 4.812 0 3.0 1e-06 
3.0 4.812 0 3.0 1e-06 
0.05 4.813 0 3.0 1e-06 
3.0 4.813 0 3.0 1e-06 
0.05 4.814 0 3.0 1e-06 
3.0 4.814 0 3.0 1e-06 
0.05 4.815 0 3.0 1e-06 
3.0 4.815 0 3.0 1e-06 
0.05 4.816 0 3.0 1e-06 
3.0 4.816 0 3.0 1e-06 
0.05 4.817 0 3.0 1e-06 
3.0 4.817 0 3.0 1e-06 
0.05 4.818 0 3.0 1e-06 
3.0 4.818 0 3.0 1e-06 
0.05 4.819 0 3.0 1e-06 
3.0 4.819 0 3.0 1e-06 
0.05 4.82 0 3.0 1e-06 
3.0 4.82 0 3.0 1e-06 
0.05 4.821 0 3.0 1e-06 
3.0 4.821 0 3.0 1e-06 
0.05 4.822 0 3.0 1e-06 
3.0 4.822 0 3.0 1e-06 
0.05 4.823 0 3.0 1e-06 
3.0 4.823 0 3.0 1e-06 
0.05 4.824 0 3.0 1e-06 
3.0 4.824 0 3.0 1e-06 
0.05 4.825 0 3.0 1e-06 
3.0 4.825 0 3.0 1e-06 
0.05 4.826 0 3.0 1e-06 
3.0 4.826 0 3.0 1e-06 
0.05 4.827 0 3.0 1e-06 
3.0 4.827 0 3.0 1e-06 
0.05 4.828 0 3.0 1e-06 
3.0 4.828 0 3.0 1e-06 
0.05 4.829 0 3.0 1e-06 
3.0 4.829 0 3.0 1e-06 
0.05 4.83 0 3.0 1e-06 
3.0 4.83 0 3.0 1e-06 
0.05 4.831 0 3.0 1e-06 
3.0 4.831 0 3.0 1e-06 
0.05 4.832 0 3.0 1e-06 
3.0 4.832 0 3.0 1e-06 
0.05 4.833 0 3.0 1e-06 
3.0 4.833 0 3.0 1e-06 
0.05 4.834 0 3.0 1e-06 
3.0 4.834 0 3.0 1e-06 
0.05 4.835 0 3.0 1e-06 
3.0 4.835 0 3.0 1e-06 
0.05 4.836 0 3.0 1e-06 
3.0 4.836 0 3.0 1e-06 
0.05 4.837 0 3.0 1e-06 
3.0 4.837 0 3.0 1e-06 
0.05 4.838 0 3.0 1e-06 
3.0 4.838 0 3.0 1e-06 
0.05 4.839 0 3.0 1e-06 
3.0 4.839 0 3.0 1e-06 
0.05 4.84 0 3.0 1e-06 
3.0 4.84 0 3.0 1e-06 
0.05 4.841 0 3.0 1e-06 
3.0 4.841 0 3.0 1e-06 
0.05 4.842 0 3.0 1e-06 
3.0 4.842 0 3.0 1e-06 
0.05 4.843 0 3.0 1e-06 
3.0 4.843 0 3.0 1e-06 
0.05 4.844 0 3.0 1e-06 
3.0 4.844 0 3.0 1e-06 
0.05 4.845 0 3.0 1e-06 
3.0 4.845 0 3.0 1e-06 
0.05 4.846 0 3.0 1e-06 
3.0 4.846 0 3.0 1e-06 
0.05 4.847 0 3.0 1e-06 
3.0 4.847 0 3.0 1e-06 
0.05 4.848 0 3.0 1e-06 
3.0 4.848 0 3.0 1e-06 
0.05 4.849 0 3.0 1e-06 
3.0 4.849 0 3.0 1e-06 
0.05 4.85 0 3.0 1e-06 
3.0 4.85 0 3.0 1e-06 
0.05 4.851 0 3.0 1e-06 
3.0 4.851 0 3.0 1e-06 
0.05 4.852 0 3.0 1e-06 
3.0 4.852 0 3.0 1e-06 
0.05 4.853 0 3.0 1e-06 
3.0 4.853 0 3.0 1e-06 
0.05 4.854 0 3.0 1e-06 
3.0 4.854 0 3.0 1e-06 
0.05 4.855 0 3.0 1e-06 
3.0 4.855 0 3.0 1e-06 
0.05 4.856 0 3.0 1e-06 
3.0 4.856 0 3.0 1e-06 
0.05 4.857 0 3.0 1e-06 
3.0 4.857 0 3.0 1e-06 
0.05 4.858 0 3.0 1e-06 
3.0 4.858 0 3.0 1e-06 
0.05 4.859 0 3.0 1e-06 
3.0 4.859 0 3.0 1e-06 
0.05 4.86 0 3.0 1e-06 
3.0 4.86 0 3.0 1e-06 
0.05 4.861 0 3.0 1e-06 
3.0 4.861 0 3.0 1e-06 
0.05 4.862 0 3.0 1e-06 
3.0 4.862 0 3.0 1e-06 
0.05 4.863 0 3.0 1e-06 
3.0 4.863 0 3.0 1e-06 
0.05 4.864 0 3.0 1e-06 
3.0 4.864 0 3.0 1e-06 
0.05 4.865 0 3.0 1e-06 
3.0 4.865 0 3.0 1e-06 
0.05 4.866 0 3.0 1e-06 
3.0 4.866 0 3.0 1e-06 
0.05 4.867 0 3.0 1e-06 
3.0 4.867 0 3.0 1e-06 
0.05 4.868 0 3.0 1e-06 
3.0 4.868 0 3.0 1e-06 
0.05 4.869 0 3.0 1e-06 
3.0 4.869 0 3.0 1e-06 
0.05 4.87 0 3.0 1e-06 
3.0 4.87 0 3.0 1e-06 
0.05 4.871 0 3.0 1e-06 
3.0 4.871 0 3.0 1e-06 
0.05 4.872 0 3.0 1e-06 
3.0 4.872 0 3.0 1e-06 
0.05 4.873 0 3.0 1e-06 
3.0 4.873 0 3.0 1e-06 
0.05 4.874 0 3.0 1e-06 
3.0 4.874 0 3.0 1e-06 
0.05 4.875 0 3.0 1e-06 
3.0 4.875 0 3.0 1e-06 
0.05 4.876 0 3.0 1e-06 
3.0 4.876 0 3.0 1e-06 
0.05 4.877 0 3.0 1e-06 
3.0 4.877 0 3.0 1e-06 
0.05 4.878 0 3.0 1e-06 
3.0 4.878 0 3.0 1e-06 
0.05 4.879 0 3.0 1e-06 
3.0 4.879 0 3.0 1e-06 
0.05 4.88 0 3.0 1e-06 
3.0 4.88 0 3.0 1e-06 
0.05 4.881 0 3.0 1e-06 
3.0 4.881 0 3.0 1e-06 
0.05 4.882 0 3.0 1e-06 
3.0 4.882 0 3.0 1e-06 
0.05 4.883 0 3.0 1e-06 
3.0 4.883 0 3.0 1e-06 
0.05 4.884 0 3.0 1e-06 
3.0 4.884 0 3.0 1e-06 
0.05 4.885 0 3.0 1e-06 
3.0 4.885 0 3.0 1e-06 
0.05 4.886 0 3.0 1e-06 
3.0 4.886 0 3.0 1e-06 
0.05 4.887 0 3.0 1e-06 
3.0 4.887 0 3.0 1e-06 
0.05 4.888 0 3.0 1e-06 
3.0 4.888 0 3.0 1e-06 
0.05 4.889 0 3.0 1e-06 
3.0 4.889 0 3.0 1e-06 
0.05 4.89 0 3.0 1e-06 
3.0 4.89 0 3.0 1e-06 
0.05 4.891 0 3.0 1e-06 
3.0 4.891 0 3.0 1e-06 
0.05 4.892 0 3.0 1e-06 
3.0 4.892 0 3.0 1e-06 
0.05 4.893 0 3.0 1e-06 
3.0 4.893 0 3.0 1e-06 
0.05 4.894 0 3.0 1e-06 
3.0 4.894 0 3.0 1e-06 
0.05 4.895 0 3.0 1e-06 
3.0 4.895 0 3.0 1e-06 
0.05 4.896 0 3.0 1e-06 
3.0 4.896 0 3.0 1e-06 
0.05 4.897 0 3.0 1e-06 
3.0 4.897 0 3.0 1e-06 
0.05 4.898 0 3.0 1e-06 
3.0 4.898 0 3.0 1e-06 
0.05 4.899 0 3.0 1e-06 
3.0 4.899 0 3.0 1e-06 
0.05 4.9 0 3.0 1e-06 
3.0 4.9 0 3.0 1e-06 
0.05 4.901 0 3.0 1e-06 
3.0 4.901 0 3.0 1e-06 
0.05 4.902 0 3.0 1e-06 
3.0 4.902 0 3.0 1e-06 
0.05 4.903 0 3.0 1e-06 
3.0 4.903 0 3.0 1e-06 
0.05 4.904 0 3.0 1e-06 
3.0 4.904 0 3.0 1e-06 
0.05 4.905 0 3.0 1e-06 
3.0 4.905 0 3.0 1e-06 
0.05 4.906 0 3.0 1e-06 
3.0 4.906 0 3.0 1e-06 
0.05 4.907 0 3.0 1e-06 
3.0 4.907 0 3.0 1e-06 
0.05 4.908 0 3.0 1e-06 
3.0 4.908 0 3.0 1e-06 
0.05 4.909 0 3.0 1e-06 
3.0 4.909 0 3.0 1e-06 
0.05 4.91 0 3.0 1e-06 
3.0 4.91 0 3.0 1e-06 
0.05 4.911 0 3.0 1e-06 
3.0 4.911 0 3.0 1e-06 
0.05 4.912 0 3.0 1e-06 
3.0 4.912 0 3.0 1e-06 
0.05 4.913 0 3.0 1e-06 
3.0 4.913 0 3.0 1e-06 
0.05 4.914 0 3.0 1e-06 
3.0 4.914 0 3.0 1e-06 
0.05 4.915 0 3.0 1e-06 
3.0 4.915 0 3.0 1e-06 
0.05 4.916 0 3.0 1e-06 
3.0 4.916 0 3.0 1e-06 
0.05 4.917 0 3.0 1e-06 
3.0 4.917 0 3.0 1e-06 
0.05 4.918 0 3.0 1e-06 
3.0 4.918 0 3.0 1e-06 
0.05 4.919 0 3.0 1e-06 
3.0 4.919 0 3.0 1e-06 
0.05 4.92 0 3.0 1e-06 
3.0 4.92 0 3.0 1e-06 
0.05 4.921 0 3.0 1e-06 
3.0 4.921 0 3.0 1e-06 
0.05 4.922 0 3.0 1e-06 
3.0 4.922 0 3.0 1e-06 
0.05 4.923 0 3.0 1e-06 
3.0 4.923 0 3.0 1e-06 
0.05 4.924 0 3.0 1e-06 
3.0 4.924 0 3.0 1e-06 
0.05 4.925 0 3.0 1e-06 
3.0 4.925 0 3.0 1e-06 
0.05 4.926 0 3.0 1e-06 
3.0 4.926 0 3.0 1e-06 
0.05 4.927 0 3.0 1e-06 
3.0 4.927 0 3.0 1e-06 
0.05 4.928 0 3.0 1e-06 
3.0 4.928 0 3.0 1e-06 
0.05 4.929 0 3.0 1e-06 
3.0 4.929 0 3.0 1e-06 
0.05 4.93 0 3.0 1e-06 
3.0 4.93 0 3.0 1e-06 
0.05 4.931 0 3.0 1e-06 
3.0 4.931 0 3.0 1e-06 
0.05 4.932 0 3.0 1e-06 
3.0 4.932 0 3.0 1e-06 
0.05 4.933 0 3.0 1e-06 
3.0 4.933 0 3.0 1e-06 
0.05 4.934 0 3.0 1e-06 
3.0 4.934 0 3.0 1e-06 
0.05 4.935 0 3.0 1e-06 
3.0 4.935 0 3.0 1e-06 
0.05 4.936 0 3.0 1e-06 
3.0 4.936 0 3.0 1e-06 
0.05 4.937 0 3.0 1e-06 
3.0 4.937 0 3.0 1e-06 
0.05 4.938 0 3.0 1e-06 
3.0 4.938 0 3.0 1e-06 
0.05 4.939 0 3.0 1e-06 
3.0 4.939 0 3.0 1e-06 
0.05 4.94 0 3.0 1e-06 
3.0 4.94 0 3.0 1e-06 
0.05 4.941 0 3.0 1e-06 
3.0 4.941 0 3.0 1e-06 
0.05 4.942 0 3.0 1e-06 
3.0 4.942 0 3.0 1e-06 
0.05 4.943 0 3.0 1e-06 
3.0 4.943 0 3.0 1e-06 
0.05 4.944 0 3.0 1e-06 
3.0 4.944 0 3.0 1e-06 
0.05 4.945 0 3.0 1e-06 
3.0 4.945 0 3.0 1e-06 
0.05 4.946 0 3.0 1e-06 
3.0 4.946 0 3.0 1e-06 
0.05 4.947 0 3.0 1e-06 
3.0 4.947 0 3.0 1e-06 
0.05 4.948 0 3.0 1e-06 
3.0 4.948 0 3.0 1e-06 
0.05 4.949 0 3.0 1e-06 
3.0 4.949 0 3.0 1e-06 
0.05 4.95 0 3.0 1e-06 
3.0 4.95 0 3.0 1e-06 
0.05 4.951 0 3.0 1e-06 
3.0 4.951 0 3.0 1e-06 
0.05 4.952 0 3.0 1e-06 
3.0 4.952 0 3.0 1e-06 
0.05 4.953 0 3.0 1e-06 
3.0 4.953 0 3.0 1e-06 
0.05 4.954 0 3.0 1e-06 
3.0 4.954 0 3.0 1e-06 
0.05 4.955 0 3.0 1e-06 
3.0 4.955 0 3.0 1e-06 
0.05 4.956 0 3.0 1e-06 
3.0 4.956 0 3.0 1e-06 
0.05 4.957 0 3.0 1e-06 
3.0 4.957 0 3.0 1e-06 
0.05 4.958 0 3.0 1e-06 
3.0 4.958 0 3.0 1e-06 
0.05 4.959 0 3.0 1e-06 
3.0 4.959 0 3.0 1e-06 
0.05 4.96 0 3.0 1e-06 
3.0 4.96 0 3.0 1e-06 
0.05 4.961 0 3.0 1e-06 
3.0 4.961 0 3.0 1e-06 
0.05 4.962 0 3.0 1e-06 
3.0 4.962 0 3.0 1e-06 
0.05 4.963 0 3.0 1e-06 
3.0 4.963 0 3.0 1e-06 
0.05 4.964 0 3.0 1e-06 
3.0 4.964 0 3.0 1e-06 
0.05 4.965 0 3.0 1e-06 
3.0 4.965 0 3.0 1e-06 
0.05 4.966 0 3.0 1e-06 
3.0 4.966 0 3.0 1e-06 
0.05 4.967 0 3.0 1e-06 
3.0 4.967 0 3.0 1e-06 
0.05 4.968 0 3.0 1e-06 
3.0 4.968 0 3.0 1e-06 
0.05 4.969 0 3.0 1e-06 
3.0 4.969 0 3.0 1e-06 
0.05 4.97 0 3.0 1e-06 
3.0 4.97 0 3.0 1e-06 
0.05 4.971 0 3.0 1e-06 
3.0 4.971 0 3.0 1e-06 
0.05 4.972 0 3.0 1e-06 
3.0 4.972 0 3.0 1e-06 
0.05 4.973 0 3.0 1e-06 
3.0 4.973 0 3.0 1e-06 
0.05 4.974 0 3.0 1e-06 
3.0 4.974 0 3.0 1e-06 
0.05 4.975 0 3.0 1e-06 
3.0 4.975 0 3.0 1e-06 
0.05 4.976 0 3.0 1e-06 
3.0 4.976 0 3.0 1e-06 
0.05 4.977 0 3.0 1e-06 
3.0 4.977 0 3.0 1e-06 
0.05 4.978 0 3.0 1e-06 
3.0 4.978 0 3.0 1e-06 
0.05 4.979 0 3.0 1e-06 
3.0 4.979 0 3.0 1e-06 
0.05 4.98 0 3.0 1e-06 
3.0 4.98 0 3.0 1e-06 
0.05 4.981 0 3.0 1e-06 
3.0 4.981 0 3.0 1e-06 
0.05 4.982 0 3.0 1e-06 
3.0 4.982 0 3.0 1e-06 
0.05 4.983 0 3.0 1e-06 
3.0 4.983 0 3.0 1e-06 
0.05 4.984 0 3.0 1e-06 
3.0 4.984 0 3.0 1e-06 
0.05 4.985 0 3.0 1e-06 
3.0 4.985 0 3.0 1e-06 
0.05 4.986 0 3.0 1e-06 
3.0 4.986 0 3.0 1e-06 
0.05 4.987 0 3.0 1e-06 
3.0 4.987 0 3.0 1e-06 
0.05 4.988 0 3.0 1e-06 
3.0 4.988 0 3.0 1e-06 
0.05 4.989 0 3.0 1e-06 
3.0 4.989 0 3.0 1e-06 
0.05 4.99 0 3.0 1e-06 
3.0 4.99 0 3.0 1e-06 
0.05 4.991 0 3.0 1e-06 
3.0 4.991 0 3.0 1e-06 
0.05 4.992 0 3.0 1e-06 
3.0 4.992 0 3.0 1e-06 
0.05 4.993 0 3.0 1e-06 
3.0 4.993 0 3.0 1e-06 
0.05 4.994 0 3.0 1e-06 
3.0 4.994 0 3.0 1e-06 
0.05 4.995 0 3.0 1e-06 
3.0 4.995 0 3.0 1e-06 
0.05 4.996 0 3.0 1e-06 
3.0 4.996 0 3.0 1e-06 
0.05 4.997 0 3.0 1e-06 
3.0 4.997 0 3.0 1e-06 
0.05 4.998 0 3.0 1e-06 
3.0 4.998 0 3.0 1e-06 
0.05 4.999 0 3.0 1e-06 
3.0 4.999 0 3.0 1e-06 
.ENDDATA 
.dc sweep DATA = datadc 
.print dc X1:IDS 
.end