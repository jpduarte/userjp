*script to generate hspice simulation using cmdp, Juan Duarte 
*Date: 11/25/2015, time: 11:58:19

.option abstol=1e-6 reltol=1e-6 post ingold 
.option measform=1 
.temp 27 

.hdl "/users/jpduarte/research/BSIMIMG/code/bsimimg.va" 
.include "/users/jpduarte/research/userjp/project4/modelcards/modelcardsimple.nmos" 

.PARAM Vd_value = 0 
.PARAM Vgf_value = 0 
.PARAM Vs_value = 0 
.PARAM Vgb_value = 0 
.PARAM L_value = 1e-06 

Vd Vd 0.0 dc = Vd_value 
Vgf Vgf 0.0 dc = Vgf_value 
Vs Vs 0.0 dc = Vs_value 
Vgb Vgb 0.0 dc = Vgb_value 

X1 Vd Vgf Vs Vgb nmos1 L = 'L_value'

.DATA datadc Vd_value Vgf_value Vs_value Vgb_value L_value 
0.0 -1.5 0 -2.0 1e-06 
0.0 -1.4999 0 -2.0 1e-06 
0.0 -1.4998 0 -2.0 1e-06 
0.0 -1.4997 0 -2.0 1e-06 
0.0 -1.4996 0 -2.0 1e-06 
0.0 -1.4995 0 -2.0 1e-06 
0.0 -1.4994 0 -2.0 1e-06 
0.0 -1.4993 0 -2.0 1e-06 
0.0 -1.4992 0 -2.0 1e-06 
0.0 -1.4991 0 -2.0 1e-06 
0.0 -1.499 0 -2.0 1e-06 
0.0 -1.4989 0 -2.0 1e-06 
0.0 -1.4988 0 -2.0 1e-06 
0.0 -1.4987 0 -2.0 1e-06 
0.0 -1.4986 0 -2.0 1e-06 
0.0 -1.4985 0 -2.0 1e-06 
0.0 -1.4984 0 -2.0 1e-06 
0.0 -1.4983 0 -2.0 1e-06 
0.0 -1.4982 0 -2.0 1e-06 
0.0 -1.4981 0 -2.0 1e-06 
0.0 -1.498 0 -2.0 1e-06 
0.0 -1.4979 0 -2.0 1e-06 
0.0 -1.4978 0 -2.0 1e-06 
0.0 -1.4977 0 -2.0 1e-06 
0.0 -1.4976 0 -2.0 1e-06 
0.0 -1.4975 0 -2.0 1e-06 
0.0 -1.4974 0 -2.0 1e-06 
0.0 -1.4973 0 -2.0 1e-06 
0.0 -1.4972 0 -2.0 1e-06 
0.0 -1.4971 0 -2.0 1e-06 
0.0 -1.497 0 -2.0 1e-06 
0.0 -1.4969 0 -2.0 1e-06 
0.0 -1.4968 0 -2.0 1e-06 
0.0 -1.4967 0 -2.0 1e-06 
0.0 -1.4966 0 -2.0 1e-06 
0.0 -1.4965 0 -2.0 1e-06 
0.0 -1.4964 0 -2.0 1e-06 
0.0 -1.4963 0 -2.0 1e-06 
0.0 -1.4962 0 -2.0 1e-06 
0.0 -1.4961 0 -2.0 1e-06 
0.0 -1.496 0 -2.0 1e-06 
0.0 -1.4959 0 -2.0 1e-06 
0.0 -1.4958 0 -2.0 1e-06 
0.0 -1.4957 0 -2.0 1e-06 
0.0 -1.4956 0 -2.0 1e-06 
0.0 -1.4955 0 -2.0 1e-06 
0.0 -1.4954 0 -2.0 1e-06 
0.0 -1.4953 0 -2.0 1e-06 
0.0 -1.4952 0 -2.0 1e-06 
0.0 -1.4951 0 -2.0 1e-06 
0.0 -1.495 0 -2.0 1e-06 
0.0 -1.4949 0 -2.0 1e-06 
0.0 -1.4948 0 -2.0 1e-06 
0.0 -1.4947 0 -2.0 1e-06 
0.0 -1.4946 0 -2.0 1e-06 
0.0 -1.4945 0 -2.0 1e-06 
0.0 -1.4944 0 -2.0 1e-06 
0.0 -1.4943 0 -2.0 1e-06 
0.0 -1.4942 0 -2.0 1e-06 
0.0 -1.4941 0 -2.0 1e-06 
0.0 -1.494 0 -2.0 1e-06 
0.0 -1.4939 0 -2.0 1e-06 
0.0 -1.4938 0 -2.0 1e-06 
0.0 -1.4937 0 -2.0 1e-06 
0.0 -1.4936 0 -2.0 1e-06 
0.0 -1.4935 0 -2.0 1e-06 
0.0 -1.4934 0 -2.0 1e-06 
0.0 -1.4933 0 -2.0 1e-06 
0.0 -1.4932 0 -2.0 1e-06 
0.0 -1.4931 0 -2.0 1e-06 
0.0 -1.493 0 -2.0 1e-06 
0.0 -1.4929 0 -2.0 1e-06 
0.0 -1.4928 0 -2.0 1e-06 
0.0 -1.4927 0 -2.0 1e-06 
0.0 -1.4926 0 -2.0 1e-06 
0.0 -1.4925 0 -2.0 1e-06 
0.0 -1.4924 0 -2.0 1e-06 
0.0 -1.4923 0 -2.0 1e-06 
0.0 -1.4922 0 -2.0 1e-06 
0.0 -1.4921 0 -2.0 1e-06 
0.0 -1.492 0 -2.0 1e-06 
0.0 -1.4919 0 -2.0 1e-06 
0.0 -1.4918 0 -2.0 1e-06 
0.0 -1.4917 0 -2.0 1e-06 
0.0 -1.4916 0 -2.0 1e-06 
0.0 -1.4915 0 -2.0 1e-06 
0.0 -1.4914 0 -2.0 1e-06 
0.0 -1.4913 0 -2.0 1e-06 
0.0 -1.4912 0 -2.0 1e-06 
0.0 -1.4911 0 -2.0 1e-06 
0.0 -1.491 0 -2.0 1e-06 
0.0 -1.4909 0 -2.0 1e-06 
0.0 -1.4908 0 -2.0 1e-06 
0.0 -1.4907 0 -2.0 1e-06 
0.0 -1.4906 0 -2.0 1e-06 
0.0 -1.4905 0 -2.0 1e-06 
0.0 -1.4904 0 -2.0 1e-06 
0.0 -1.4903 0 -2.0 1e-06 
0.0 -1.4902 0 -2.0 1e-06 
0.0 -1.4901 0 -2.0 1e-06 
0.0 -1.49 0 -2.0 1e-06 
0.0 -1.4899 0 -2.0 1e-06 
0.0 -1.4898 0 -2.0 1e-06 
0.0 -1.4897 0 -2.0 1e-06 
0.0 -1.4896 0 -2.0 1e-06 
0.0 -1.4895 0 -2.0 1e-06 
0.0 -1.4894 0 -2.0 1e-06 
0.0 -1.4893 0 -2.0 1e-06 
0.0 -1.4892 0 -2.0 1e-06 
0.0 -1.4891 0 -2.0 1e-06 
0.0 -1.489 0 -2.0 1e-06 
0.0 -1.4889 0 -2.0 1e-06 
0.0 -1.4888 0 -2.0 1e-06 
0.0 -1.4887 0 -2.0 1e-06 
0.0 -1.4886 0 -2.0 1e-06 
0.0 -1.4885 0 -2.0 1e-06 
0.0 -1.4884 0 -2.0 1e-06 
0.0 -1.4883 0 -2.0 1e-06 
0.0 -1.4882 0 -2.0 1e-06 
0.0 -1.4881 0 -2.0 1e-06 
0.0 -1.488 0 -2.0 1e-06 
0.0 -1.4879 0 -2.0 1e-06 
0.0 -1.4878 0 -2.0 1e-06 
0.0 -1.4877 0 -2.0 1e-06 
0.0 -1.4876 0 -2.0 1e-06 
0.0 -1.4875 0 -2.0 1e-06 
0.0 -1.4874 0 -2.0 1e-06 
0.0 -1.4873 0 -2.0 1e-06 
0.0 -1.4872 0 -2.0 1e-06 
0.0 -1.4871 0 -2.0 1e-06 
0.0 -1.487 0 -2.0 1e-06 
0.0 -1.4869 0 -2.0 1e-06 
0.0 -1.4868 0 -2.0 1e-06 
0.0 -1.4867 0 -2.0 1e-06 
0.0 -1.4866 0 -2.0 1e-06 
0.0 -1.4865 0 -2.0 1e-06 
0.0 -1.4864 0 -2.0 1e-06 
0.0 -1.4863 0 -2.0 1e-06 
0.0 -1.4862 0 -2.0 1e-06 
0.0 -1.4861 0 -2.0 1e-06 
0.0 -1.486 0 -2.0 1e-06 
0.0 -1.4859 0 -2.0 1e-06 
0.0 -1.4858 0 -2.0 1e-06 
0.0 -1.4857 0 -2.0 1e-06 
0.0 -1.4856 0 -2.0 1e-06 
0.0 -1.4855 0 -2.0 1e-06 
0.0 -1.4854 0 -2.0 1e-06 
0.0 -1.4853 0 -2.0 1e-06 
0.0 -1.4852 0 -2.0 1e-06 
0.0 -1.4851 0 -2.0 1e-06 
0.0 -1.485 0 -2.0 1e-06 
0.0 -1.4849 0 -2.0 1e-06 
0.0 -1.4848 0 -2.0 1e-06 
0.0 -1.4847 0 -2.0 1e-06 
0.0 -1.4846 0 -2.0 1e-06 
0.0 -1.4845 0 -2.0 1e-06 
0.0 -1.4844 0 -2.0 1e-06 
0.0 -1.4843 0 -2.0 1e-06 
0.0 -1.4842 0 -2.0 1e-06 
0.0 -1.4841 0 -2.0 1e-06 
0.0 -1.484 0 -2.0 1e-06 
0.0 -1.4839 0 -2.0 1e-06 
0.0 -1.4838 0 -2.0 1e-06 
0.0 -1.4837 0 -2.0 1e-06 
0.0 -1.4836 0 -2.0 1e-06 
0.0 -1.4835 0 -2.0 1e-06 
0.0 -1.4834 0 -2.0 1e-06 
0.0 -1.4833 0 -2.0 1e-06 
0.0 -1.4832 0 -2.0 1e-06 
0.0 -1.4831 0 -2.0 1e-06 
0.0 -1.483 0 -2.0 1e-06 
0.0 -1.4829 0 -2.0 1e-06 
0.0 -1.4828 0 -2.0 1e-06 
0.0 -1.4827 0 -2.0 1e-06 
0.0 -1.4826 0 -2.0 1e-06 
0.0 -1.4825 0 -2.0 1e-06 
0.0 -1.4824 0 -2.0 1e-06 
0.0 -1.4823 0 -2.0 1e-06 
0.0 -1.4822 0 -2.0 1e-06 
0.0 -1.4821 0 -2.0 1e-06 
0.0 -1.482 0 -2.0 1e-06 
0.0 -1.4819 0 -2.0 1e-06 
0.0 -1.4818 0 -2.0 1e-06 
0.0 -1.4817 0 -2.0 1e-06 
0.0 -1.4816 0 -2.0 1e-06 
0.0 -1.4815 0 -2.0 1e-06 
0.0 -1.4814 0 -2.0 1e-06 
0.0 -1.4813 0 -2.0 1e-06 
0.0 -1.4812 0 -2.0 1e-06 
0.0 -1.4811 0 -2.0 1e-06 
0.0 -1.481 0 -2.0 1e-06 
0.0 -1.4809 0 -2.0 1e-06 
0.0 -1.4808 0 -2.0 1e-06 
0.0 -1.4807 0 -2.0 1e-06 
0.0 -1.4806 0 -2.0 1e-06 
0.0 -1.4805 0 -2.0 1e-06 
0.0 -1.4804 0 -2.0 1e-06 
0.0 -1.4803 0 -2.0 1e-06 
0.0 -1.4802 0 -2.0 1e-06 
0.0 -1.4801 0 -2.0 1e-06 
0.0 -1.48 0 -2.0 1e-06 
0.0 -1.4799 0 -2.0 1e-06 
0.0 -1.4798 0 -2.0 1e-06 
0.0 -1.4797 0 -2.0 1e-06 
0.0 -1.4796 0 -2.0 1e-06 
0.0 -1.4795 0 -2.0 1e-06 
0.0 -1.4794 0 -2.0 1e-06 
0.0 -1.4793 0 -2.0 1e-06 
0.0 -1.4792 0 -2.0 1e-06 
0.0 -1.4791 0 -2.0 1e-06 
0.0 -1.479 0 -2.0 1e-06 
0.0 -1.4789 0 -2.0 1e-06 
0.0 -1.4788 0 -2.0 1e-06 
0.0 -1.4787 0 -2.0 1e-06 
0.0 -1.4786 0 -2.0 1e-06 
0.0 -1.4785 0 -2.0 1e-06 
0.0 -1.4784 0 -2.0 1e-06 
0.0 -1.4783 0 -2.0 1e-06 
0.0 -1.4782 0 -2.0 1e-06 
0.0 -1.4781 0 -2.0 1e-06 
0.0 -1.478 0 -2.0 1e-06 
0.0 -1.4779 0 -2.0 1e-06 
0.0 -1.4778 0 -2.0 1e-06 
0.0 -1.4777 0 -2.0 1e-06 
0.0 -1.4776 0 -2.0 1e-06 
0.0 -1.4775 0 -2.0 1e-06 
0.0 -1.4774 0 -2.0 1e-06 
0.0 -1.4773 0 -2.0 1e-06 
0.0 -1.4772 0 -2.0 1e-06 
0.0 -1.4771 0 -2.0 1e-06 
0.0 -1.477 0 -2.0 1e-06 
0.0 -1.4769 0 -2.0 1e-06 
0.0 -1.4768 0 -2.0 1e-06 
0.0 -1.4767 0 -2.0 1e-06 
0.0 -1.4766 0 -2.0 1e-06 
0.0 -1.4765 0 -2.0 1e-06 
0.0 -1.4764 0 -2.0 1e-06 
0.0 -1.4763 0 -2.0 1e-06 
0.0 -1.4762 0 -2.0 1e-06 
0.0 -1.4761 0 -2.0 1e-06 
0.0 -1.476 0 -2.0 1e-06 
0.0 -1.4759 0 -2.0 1e-06 
0.0 -1.4758 0 -2.0 1e-06 
0.0 -1.4757 0 -2.0 1e-06 
0.0 -1.4756 0 -2.0 1e-06 
0.0 -1.4755 0 -2.0 1e-06 
0.0 -1.4754 0 -2.0 1e-06 
0.0 -1.4753 0 -2.0 1e-06 
0.0 -1.4752 0 -2.0 1e-06 
0.0 -1.4751 0 -2.0 1e-06 
0.0 -1.475 0 -2.0 1e-06 
0.0 -1.4749 0 -2.0 1e-06 
0.0 -1.4748 0 -2.0 1e-06 
0.0 -1.4747 0 -2.0 1e-06 
0.0 -1.4746 0 -2.0 1e-06 
0.0 -1.4745 0 -2.0 1e-06 
0.0 -1.4744 0 -2.0 1e-06 
0.0 -1.4743 0 -2.0 1e-06 
0.0 -1.4742 0 -2.0 1e-06 
0.0 -1.4741 0 -2.0 1e-06 
0.0 -1.474 0 -2.0 1e-06 
0.0 -1.4739 0 -2.0 1e-06 
0.0 -1.4738 0 -2.0 1e-06 
0.0 -1.4737 0 -2.0 1e-06 
0.0 -1.4736 0 -2.0 1e-06 
0.0 -1.4735 0 -2.0 1e-06 
0.0 -1.4734 0 -2.0 1e-06 
0.0 -1.4733 0 -2.0 1e-06 
0.0 -1.4732 0 -2.0 1e-06 
0.0 -1.4731 0 -2.0 1e-06 
0.0 -1.473 0 -2.0 1e-06 
0.0 -1.4729 0 -2.0 1e-06 
0.0 -1.4728 0 -2.0 1e-06 
0.0 -1.4727 0 -2.0 1e-06 
0.0 -1.4726 0 -2.0 1e-06 
0.0 -1.4725 0 -2.0 1e-06 
0.0 -1.4724 0 -2.0 1e-06 
0.0 -1.4723 0 -2.0 1e-06 
0.0 -1.4722 0 -2.0 1e-06 
0.0 -1.4721 0 -2.0 1e-06 
0.0 -1.472 0 -2.0 1e-06 
0.0 -1.4719 0 -2.0 1e-06 
0.0 -1.4718 0 -2.0 1e-06 
0.0 -1.4717 0 -2.0 1e-06 
0.0 -1.4716 0 -2.0 1e-06 
0.0 -1.4715 0 -2.0 1e-06 
0.0 -1.4714 0 -2.0 1e-06 
0.0 -1.4713 0 -2.0 1e-06 
0.0 -1.4712 0 -2.0 1e-06 
0.0 -1.4711 0 -2.0 1e-06 
0.0 -1.471 0 -2.0 1e-06 
0.0 -1.4709 0 -2.0 1e-06 
0.0 -1.4708 0 -2.0 1e-06 
0.0 -1.4707 0 -2.0 1e-06 
0.0 -1.4706 0 -2.0 1e-06 
0.0 -1.4705 0 -2.0 1e-06 
0.0 -1.4704 0 -2.0 1e-06 
0.0 -1.4703 0 -2.0 1e-06 
0.0 -1.4702 0 -2.0 1e-06 
0.0 -1.4701 0 -2.0 1e-06 
0.0 -1.47 0 -2.0 1e-06 
0.0 -1.4699 0 -2.0 1e-06 
0.0 -1.4698 0 -2.0 1e-06 
0.0 -1.4697 0 -2.0 1e-06 
0.0 -1.4696 0 -2.0 1e-06 
0.0 -1.4695 0 -2.0 1e-06 
0.0 -1.4694 0 -2.0 1e-06 
0.0 -1.4693 0 -2.0 1e-06 
0.0 -1.4692 0 -2.0 1e-06 
0.0 -1.4691 0 -2.0 1e-06 
0.0 -1.469 0 -2.0 1e-06 
0.0 -1.4689 0 -2.0 1e-06 
0.0 -1.4688 0 -2.0 1e-06 
0.0 -1.4687 0 -2.0 1e-06 
0.0 -1.4686 0 -2.0 1e-06 
0.0 -1.4685 0 -2.0 1e-06 
0.0 -1.4684 0 -2.0 1e-06 
0.0 -1.4683 0 -2.0 1e-06 
0.0 -1.4682 0 -2.0 1e-06 
0.0 -1.4681 0 -2.0 1e-06 
0.0 -1.468 0 -2.0 1e-06 
0.0 -1.4679 0 -2.0 1e-06 
0.0 -1.4678 0 -2.0 1e-06 
0.0 -1.4677 0 -2.0 1e-06 
0.0 -1.4676 0 -2.0 1e-06 
0.0 -1.4675 0 -2.0 1e-06 
0.0 -1.4674 0 -2.0 1e-06 
0.0 -1.4673 0 -2.0 1e-06 
0.0 -1.4672 0 -2.0 1e-06 
0.0 -1.4671 0 -2.0 1e-06 
0.0 -1.467 0 -2.0 1e-06 
0.0 -1.4669 0 -2.0 1e-06 
0.0 -1.4668 0 -2.0 1e-06 
0.0 -1.4667 0 -2.0 1e-06 
0.0 -1.4666 0 -2.0 1e-06 
0.0 -1.4665 0 -2.0 1e-06 
0.0 -1.4664 0 -2.0 1e-06 
0.0 -1.4663 0 -2.0 1e-06 
0.0 -1.4662 0 -2.0 1e-06 
0.0 -1.4661 0 -2.0 1e-06 
0.0 -1.466 0 -2.0 1e-06 
0.0 -1.4659 0 -2.0 1e-06 
0.0 -1.4658 0 -2.0 1e-06 
0.0 -1.4657 0 -2.0 1e-06 
0.0 -1.4656 0 -2.0 1e-06 
0.0 -1.4655 0 -2.0 1e-06 
0.0 -1.4654 0 -2.0 1e-06 
0.0 -1.4653 0 -2.0 1e-06 
0.0 -1.4652 0 -2.0 1e-06 
0.0 -1.4651 0 -2.0 1e-06 
0.0 -1.465 0 -2.0 1e-06 
0.0 -1.4649 0 -2.0 1e-06 
0.0 -1.4648 0 -2.0 1e-06 
0.0 -1.4647 0 -2.0 1e-06 
0.0 -1.4646 0 -2.0 1e-06 
0.0 -1.4645 0 -2.0 1e-06 
0.0 -1.4644 0 -2.0 1e-06 
0.0 -1.4643 0 -2.0 1e-06 
0.0 -1.4642 0 -2.0 1e-06 
0.0 -1.4641 0 -2.0 1e-06 
0.0 -1.464 0 -2.0 1e-06 
0.0 -1.4639 0 -2.0 1e-06 
0.0 -1.4638 0 -2.0 1e-06 
0.0 -1.4637 0 -2.0 1e-06 
0.0 -1.4636 0 -2.0 1e-06 
0.0 -1.4635 0 -2.0 1e-06 
0.0 -1.4634 0 -2.0 1e-06 
0.0 -1.4633 0 -2.0 1e-06 
0.0 -1.4632 0 -2.0 1e-06 
0.0 -1.4631 0 -2.0 1e-06 
0.0 -1.463 0 -2.0 1e-06 
0.0 -1.4629 0 -2.0 1e-06 
0.0 -1.4628 0 -2.0 1e-06 
0.0 -1.4627 0 -2.0 1e-06 
0.0 -1.4626 0 -2.0 1e-06 
0.0 -1.4625 0 -2.0 1e-06 
0.0 -1.4624 0 -2.0 1e-06 
0.0 -1.4623 0 -2.0 1e-06 
0.0 -1.4622 0 -2.0 1e-06 
0.0 -1.4621 0 -2.0 1e-06 
0.0 -1.462 0 -2.0 1e-06 
0.0 -1.4619 0 -2.0 1e-06 
0.0 -1.4618 0 -2.0 1e-06 
0.0 -1.4617 0 -2.0 1e-06 
0.0 -1.4616 0 -2.0 1e-06 
0.0 -1.4615 0 -2.0 1e-06 
0.0 -1.4614 0 -2.0 1e-06 
0.0 -1.4613 0 -2.0 1e-06 
0.0 -1.4612 0 -2.0 1e-06 
0.0 -1.4611 0 -2.0 1e-06 
0.0 -1.461 0 -2.0 1e-06 
0.0 -1.4609 0 -2.0 1e-06 
0.0 -1.4608 0 -2.0 1e-06 
0.0 -1.4607 0 -2.0 1e-06 
0.0 -1.4606 0 -2.0 1e-06 
0.0 -1.4605 0 -2.0 1e-06 
0.0 -1.4604 0 -2.0 1e-06 
0.0 -1.4603 0 -2.0 1e-06 
0.0 -1.4602 0 -2.0 1e-06 
0.0 -1.4601 0 -2.0 1e-06 
0.0 -1.46 0 -2.0 1e-06 
0.0 -1.4599 0 -2.0 1e-06 
0.0 -1.4598 0 -2.0 1e-06 
0.0 -1.4597 0 -2.0 1e-06 
0.0 -1.4596 0 -2.0 1e-06 
0.0 -1.4595 0 -2.0 1e-06 
0.0 -1.4594 0 -2.0 1e-06 
0.0 -1.4593 0 -2.0 1e-06 
0.0 -1.4592 0 -2.0 1e-06 
0.0 -1.4591 0 -2.0 1e-06 
0.0 -1.459 0 -2.0 1e-06 
0.0 -1.4589 0 -2.0 1e-06 
0.0 -1.4588 0 -2.0 1e-06 
0.0 -1.4587 0 -2.0 1e-06 
0.0 -1.4586 0 -2.0 1e-06 
0.0 -1.4585 0 -2.0 1e-06 
0.0 -1.4584 0 -2.0 1e-06 
0.0 -1.4583 0 -2.0 1e-06 
0.0 -1.4582 0 -2.0 1e-06 
0.0 -1.4581 0 -2.0 1e-06 
0.0 -1.458 0 -2.0 1e-06 
0.0 -1.4579 0 -2.0 1e-06 
0.0 -1.4578 0 -2.0 1e-06 
0.0 -1.4577 0 -2.0 1e-06 
0.0 -1.4576 0 -2.0 1e-06 
0.0 -1.4575 0 -2.0 1e-06 
0.0 -1.4574 0 -2.0 1e-06 
0.0 -1.4573 0 -2.0 1e-06 
0.0 -1.4572 0 -2.0 1e-06 
0.0 -1.4571 0 -2.0 1e-06 
0.0 -1.457 0 -2.0 1e-06 
0.0 -1.4569 0 -2.0 1e-06 
0.0 -1.4568 0 -2.0 1e-06 
0.0 -1.4567 0 -2.0 1e-06 
0.0 -1.4566 0 -2.0 1e-06 
0.0 -1.4565 0 -2.0 1e-06 
0.0 -1.4564 0 -2.0 1e-06 
0.0 -1.4563 0 -2.0 1e-06 
0.0 -1.4562 0 -2.0 1e-06 
0.0 -1.4561 0 -2.0 1e-06 
0.0 -1.456 0 -2.0 1e-06 
0.0 -1.4559 0 -2.0 1e-06 
0.0 -1.4558 0 -2.0 1e-06 
0.0 -1.4557 0 -2.0 1e-06 
0.0 -1.4556 0 -2.0 1e-06 
0.0 -1.4555 0 -2.0 1e-06 
0.0 -1.4554 0 -2.0 1e-06 
0.0 -1.4553 0 -2.0 1e-06 
0.0 -1.4552 0 -2.0 1e-06 
0.0 -1.4551 0 -2.0 1e-06 
0.0 -1.455 0 -2.0 1e-06 
0.0 -1.4549 0 -2.0 1e-06 
0.0 -1.4548 0 -2.0 1e-06 
0.0 -1.4547 0 -2.0 1e-06 
0.0 -1.4546 0 -2.0 1e-06 
0.0 -1.4545 0 -2.0 1e-06 
0.0 -1.4544 0 -2.0 1e-06 
0.0 -1.4543 0 -2.0 1e-06 
0.0 -1.4542 0 -2.0 1e-06 
0.0 -1.4541 0 -2.0 1e-06 
0.0 -1.454 0 -2.0 1e-06 
0.0 -1.4539 0 -2.0 1e-06 
0.0 -1.4538 0 -2.0 1e-06 
0.0 -1.4537 0 -2.0 1e-06 
0.0 -1.4536 0 -2.0 1e-06 
0.0 -1.4535 0 -2.0 1e-06 
0.0 -1.4534 0 -2.0 1e-06 
0.0 -1.4533 0 -2.0 1e-06 
0.0 -1.4532 0 -2.0 1e-06 
0.0 -1.4531 0 -2.0 1e-06 
0.0 -1.453 0 -2.0 1e-06 
0.0 -1.4529 0 -2.0 1e-06 
0.0 -1.4528 0 -2.0 1e-06 
0.0 -1.4527 0 -2.0 1e-06 
0.0 -1.4526 0 -2.0 1e-06 
0.0 -1.4525 0 -2.0 1e-06 
0.0 -1.4524 0 -2.0 1e-06 
0.0 -1.4523 0 -2.0 1e-06 
0.0 -1.4522 0 -2.0 1e-06 
0.0 -1.4521 0 -2.0 1e-06 
0.0 -1.452 0 -2.0 1e-06 
0.0 -1.4519 0 -2.0 1e-06 
0.0 -1.4518 0 -2.0 1e-06 
0.0 -1.4517 0 -2.0 1e-06 
0.0 -1.4516 0 -2.0 1e-06 
0.0 -1.4515 0 -2.0 1e-06 
0.0 -1.4514 0 -2.0 1e-06 
0.0 -1.4513 0 -2.0 1e-06 
0.0 -1.4512 0 -2.0 1e-06 
0.0 -1.4511 0 -2.0 1e-06 
0.0 -1.451 0 -2.0 1e-06 
0.0 -1.4509 0 -2.0 1e-06 
0.0 -1.4508 0 -2.0 1e-06 
0.0 -1.4507 0 -2.0 1e-06 
0.0 -1.4506 0 -2.0 1e-06 
0.0 -1.4505 0 -2.0 1e-06 
0.0 -1.4504 0 -2.0 1e-06 
0.0 -1.4503 0 -2.0 1e-06 
0.0 -1.4502 0 -2.0 1e-06 
0.0 -1.4501 0 -2.0 1e-06 
0.0 -1.45 0 -2.0 1e-06 
0.0 -1.4499 0 -2.0 1e-06 
0.0 -1.4498 0 -2.0 1e-06 
0.0 -1.4497 0 -2.0 1e-06 
0.0 -1.4496 0 -2.0 1e-06 
0.0 -1.4495 0 -2.0 1e-06 
0.0 -1.4494 0 -2.0 1e-06 
0.0 -1.4493 0 -2.0 1e-06 
0.0 -1.4492 0 -2.0 1e-06 
0.0 -1.4491 0 -2.0 1e-06 
0.0 -1.449 0 -2.0 1e-06 
0.0 -1.4489 0 -2.0 1e-06 
0.0 -1.4488 0 -2.0 1e-06 
0.0 -1.4487 0 -2.0 1e-06 
0.0 -1.4486 0 -2.0 1e-06 
0.0 -1.4485 0 -2.0 1e-06 
0.0 -1.4484 0 -2.0 1e-06 
0.0 -1.4483 0 -2.0 1e-06 
0.0 -1.4482 0 -2.0 1e-06 
0.0 -1.4481 0 -2.0 1e-06 
0.0 -1.448 0 -2.0 1e-06 
0.0 -1.4479 0 -2.0 1e-06 
0.0 -1.4478 0 -2.0 1e-06 
0.0 -1.4477 0 -2.0 1e-06 
0.0 -1.4476 0 -2.0 1e-06 
0.0 -1.4475 0 -2.0 1e-06 
0.0 -1.4474 0 -2.0 1e-06 
0.0 -1.4473 0 -2.0 1e-06 
0.0 -1.4472 0 -2.0 1e-06 
0.0 -1.4471 0 -2.0 1e-06 
0.0 -1.447 0 -2.0 1e-06 
0.0 -1.4469 0 -2.0 1e-06 
0.0 -1.4468 0 -2.0 1e-06 
0.0 -1.4467 0 -2.0 1e-06 
0.0 -1.4466 0 -2.0 1e-06 
0.0 -1.4465 0 -2.0 1e-06 
0.0 -1.4464 0 -2.0 1e-06 
0.0 -1.4463 0 -2.0 1e-06 
0.0 -1.4462 0 -2.0 1e-06 
0.0 -1.4461 0 -2.0 1e-06 
0.0 -1.446 0 -2.0 1e-06 
0.0 -1.4459 0 -2.0 1e-06 
0.0 -1.4458 0 -2.0 1e-06 
0.0 -1.4457 0 -2.0 1e-06 
0.0 -1.4456 0 -2.0 1e-06 
0.0 -1.4455 0 -2.0 1e-06 
0.0 -1.4454 0 -2.0 1e-06 
0.0 -1.4453 0 -2.0 1e-06 
0.0 -1.4452 0 -2.0 1e-06 
0.0 -1.4451 0 -2.0 1e-06 
0.0 -1.445 0 -2.0 1e-06 
0.0 -1.4449 0 -2.0 1e-06 
0.0 -1.4448 0 -2.0 1e-06 
0.0 -1.4447 0 -2.0 1e-06 
0.0 -1.4446 0 -2.0 1e-06 
0.0 -1.4445 0 -2.0 1e-06 
0.0 -1.4444 0 -2.0 1e-06 
0.0 -1.4443 0 -2.0 1e-06 
0.0 -1.4442 0 -2.0 1e-06 
0.0 -1.4441 0 -2.0 1e-06 
0.0 -1.444 0 -2.0 1e-06 
0.0 -1.4439 0 -2.0 1e-06 
0.0 -1.4438 0 -2.0 1e-06 
0.0 -1.4437 0 -2.0 1e-06 
0.0 -1.4436 0 -2.0 1e-06 
0.0 -1.4435 0 -2.0 1e-06 
0.0 -1.4434 0 -2.0 1e-06 
0.0 -1.4433 0 -2.0 1e-06 
0.0 -1.4432 0 -2.0 1e-06 
0.0 -1.4431 0 -2.0 1e-06 
0.0 -1.443 0 -2.0 1e-06 
0.0 -1.4429 0 -2.0 1e-06 
0.0 -1.4428 0 -2.0 1e-06 
0.0 -1.4427 0 -2.0 1e-06 
0.0 -1.4426 0 -2.0 1e-06 
0.0 -1.4425 0 -2.0 1e-06 
0.0 -1.4424 0 -2.0 1e-06 
0.0 -1.4423 0 -2.0 1e-06 
0.0 -1.4422 0 -2.0 1e-06 
0.0 -1.4421 0 -2.0 1e-06 
0.0 -1.442 0 -2.0 1e-06 
0.0 -1.4419 0 -2.0 1e-06 
0.0 -1.4418 0 -2.0 1e-06 
0.0 -1.4417 0 -2.0 1e-06 
0.0 -1.4416 0 -2.0 1e-06 
0.0 -1.4415 0 -2.0 1e-06 
0.0 -1.4414 0 -2.0 1e-06 
0.0 -1.4413 0 -2.0 1e-06 
0.0 -1.4412 0 -2.0 1e-06 
0.0 -1.4411 0 -2.0 1e-06 
0.0 -1.441 0 -2.0 1e-06 
0.0 -1.4409 0 -2.0 1e-06 
0.0 -1.4408 0 -2.0 1e-06 
0.0 -1.4407 0 -2.0 1e-06 
0.0 -1.4406 0 -2.0 1e-06 
0.0 -1.4405 0 -2.0 1e-06 
0.0 -1.4404 0 -2.0 1e-06 
0.0 -1.4403 0 -2.0 1e-06 
0.0 -1.4402 0 -2.0 1e-06 
0.0 -1.4401 0 -2.0 1e-06 
0.0 -1.44 0 -2.0 1e-06 
0.0 -1.4399 0 -2.0 1e-06 
0.0 -1.4398 0 -2.0 1e-06 
0.0 -1.4397 0 -2.0 1e-06 
0.0 -1.4396 0 -2.0 1e-06 
0.0 -1.4395 0 -2.0 1e-06 
0.0 -1.4394 0 -2.0 1e-06 
0.0 -1.4393 0 -2.0 1e-06 
0.0 -1.4392 0 -2.0 1e-06 
0.0 -1.4391 0 -2.0 1e-06 
0.0 -1.439 0 -2.0 1e-06 
0.0 -1.4389 0 -2.0 1e-06 
0.0 -1.4388 0 -2.0 1e-06 
0.0 -1.4387 0 -2.0 1e-06 
0.0 -1.4386 0 -2.0 1e-06 
0.0 -1.4385 0 -2.0 1e-06 
0.0 -1.4384 0 -2.0 1e-06 
0.0 -1.4383 0 -2.0 1e-06 
0.0 -1.4382 0 -2.0 1e-06 
0.0 -1.4381 0 -2.0 1e-06 
0.0 -1.438 0 -2.0 1e-06 
0.0 -1.4379 0 -2.0 1e-06 
0.0 -1.4378 0 -2.0 1e-06 
0.0 -1.4377 0 -2.0 1e-06 
0.0 -1.4376 0 -2.0 1e-06 
0.0 -1.4375 0 -2.0 1e-06 
0.0 -1.4374 0 -2.0 1e-06 
0.0 -1.4373 0 -2.0 1e-06 
0.0 -1.4372 0 -2.0 1e-06 
0.0 -1.4371 0 -2.0 1e-06 
0.0 -1.437 0 -2.0 1e-06 
0.0 -1.4369 0 -2.0 1e-06 
0.0 -1.4368 0 -2.0 1e-06 
0.0 -1.4367 0 -2.0 1e-06 
0.0 -1.4366 0 -2.0 1e-06 
0.0 -1.4365 0 -2.0 1e-06 
0.0 -1.4364 0 -2.0 1e-06 
0.0 -1.4363 0 -2.0 1e-06 
0.0 -1.4362 0 -2.0 1e-06 
0.0 -1.4361 0 -2.0 1e-06 
0.0 -1.436 0 -2.0 1e-06 
0.0 -1.4359 0 -2.0 1e-06 
0.0 -1.4358 0 -2.0 1e-06 
0.0 -1.4357 0 -2.0 1e-06 
0.0 -1.4356 0 -2.0 1e-06 
0.0 -1.4355 0 -2.0 1e-06 
0.0 -1.4354 0 -2.0 1e-06 
0.0 -1.4353 0 -2.0 1e-06 
0.0 -1.4352 0 -2.0 1e-06 
0.0 -1.4351 0 -2.0 1e-06 
0.0 -1.435 0 -2.0 1e-06 
0.0 -1.4349 0 -2.0 1e-06 
0.0 -1.4348 0 -2.0 1e-06 
0.0 -1.4347 0 -2.0 1e-06 
0.0 -1.4346 0 -2.0 1e-06 
0.0 -1.4345 0 -2.0 1e-06 
0.0 -1.4344 0 -2.0 1e-06 
0.0 -1.4343 0 -2.0 1e-06 
0.0 -1.4342 0 -2.0 1e-06 
0.0 -1.4341 0 -2.0 1e-06 
0.0 -1.434 0 -2.0 1e-06 
0.0 -1.4339 0 -2.0 1e-06 
0.0 -1.4338 0 -2.0 1e-06 
0.0 -1.4337 0 -2.0 1e-06 
0.0 -1.4336 0 -2.0 1e-06 
0.0 -1.4335 0 -2.0 1e-06 
0.0 -1.4334 0 -2.0 1e-06 
0.0 -1.4333 0 -2.0 1e-06 
0.0 -1.4332 0 -2.0 1e-06 
0.0 -1.4331 0 -2.0 1e-06 
0.0 -1.433 0 -2.0 1e-06 
0.0 -1.4329 0 -2.0 1e-06 
0.0 -1.4328 0 -2.0 1e-06 
0.0 -1.4327 0 -2.0 1e-06 
0.0 -1.4326 0 -2.0 1e-06 
0.0 -1.4325 0 -2.0 1e-06 
0.0 -1.4324 0 -2.0 1e-06 
0.0 -1.4323 0 -2.0 1e-06 
0.0 -1.4322 0 -2.0 1e-06 
0.0 -1.4321 0 -2.0 1e-06 
0.0 -1.432 0 -2.0 1e-06 
0.0 -1.4319 0 -2.0 1e-06 
0.0 -1.4318 0 -2.0 1e-06 
0.0 -1.4317 0 -2.0 1e-06 
0.0 -1.4316 0 -2.0 1e-06 
0.0 -1.4315 0 -2.0 1e-06 
0.0 -1.4314 0 -2.0 1e-06 
0.0 -1.4313 0 -2.0 1e-06 
0.0 -1.4312 0 -2.0 1e-06 
0.0 -1.4311 0 -2.0 1e-06 
0.0 -1.431 0 -2.0 1e-06 
0.0 -1.4309 0 -2.0 1e-06 
0.0 -1.4308 0 -2.0 1e-06 
0.0 -1.4307 0 -2.0 1e-06 
0.0 -1.4306 0 -2.0 1e-06 
0.0 -1.4305 0 -2.0 1e-06 
0.0 -1.4304 0 -2.0 1e-06 
0.0 -1.4303 0 -2.0 1e-06 
0.0 -1.4302 0 -2.0 1e-06 
0.0 -1.4301 0 -2.0 1e-06 
0.0 -1.43 0 -2.0 1e-06 
0.0 -1.4299 0 -2.0 1e-06 
0.0 -1.4298 0 -2.0 1e-06 
0.0 -1.4297 0 -2.0 1e-06 
0.0 -1.4296 0 -2.0 1e-06 
0.0 -1.4295 0 -2.0 1e-06 
0.0 -1.4294 0 -2.0 1e-06 
0.0 -1.4293 0 -2.0 1e-06 
0.0 -1.4292 0 -2.0 1e-06 
0.0 -1.4291 0 -2.0 1e-06 
0.0 -1.429 0 -2.0 1e-06 
0.0 -1.4289 0 -2.0 1e-06 
0.0 -1.4288 0 -2.0 1e-06 
0.0 -1.4287 0 -2.0 1e-06 
0.0 -1.4286 0 -2.0 1e-06 
0.0 -1.4285 0 -2.0 1e-06 
0.0 -1.4284 0 -2.0 1e-06 
0.0 -1.4283 0 -2.0 1e-06 
0.0 -1.4282 0 -2.0 1e-06 
0.0 -1.4281 0 -2.0 1e-06 
0.0 -1.428 0 -2.0 1e-06 
0.0 -1.4279 0 -2.0 1e-06 
0.0 -1.4278 0 -2.0 1e-06 
0.0 -1.4277 0 -2.0 1e-06 
0.0 -1.4276 0 -2.0 1e-06 
0.0 -1.4275 0 -2.0 1e-06 
0.0 -1.4274 0 -2.0 1e-06 
0.0 -1.4273 0 -2.0 1e-06 
0.0 -1.4272 0 -2.0 1e-06 
0.0 -1.4271 0 -2.0 1e-06 
0.0 -1.427 0 -2.0 1e-06 
0.0 -1.4269 0 -2.0 1e-06 
0.0 -1.4268 0 -2.0 1e-06 
0.0 -1.4267 0 -2.0 1e-06 
0.0 -1.4266 0 -2.0 1e-06 
0.0 -1.4265 0 -2.0 1e-06 
0.0 -1.4264 0 -2.0 1e-06 
0.0 -1.4263 0 -2.0 1e-06 
0.0 -1.4262 0 -2.0 1e-06 
0.0 -1.4261 0 -2.0 1e-06 
0.0 -1.426 0 -2.0 1e-06 
0.0 -1.4259 0 -2.0 1e-06 
0.0 -1.4258 0 -2.0 1e-06 
0.0 -1.4257 0 -2.0 1e-06 
0.0 -1.4256 0 -2.0 1e-06 
0.0 -1.4255 0 -2.0 1e-06 
0.0 -1.4254 0 -2.0 1e-06 
0.0 -1.4253 0 -2.0 1e-06 
0.0 -1.4252 0 -2.0 1e-06 
0.0 -1.4251 0 -2.0 1e-06 
0.0 -1.425 0 -2.0 1e-06 
0.0 -1.4249 0 -2.0 1e-06 
0.0 -1.4248 0 -2.0 1e-06 
0.0 -1.4247 0 -2.0 1e-06 
0.0 -1.4246 0 -2.0 1e-06 
0.0 -1.4245 0 -2.0 1e-06 
0.0 -1.4244 0 -2.0 1e-06 
0.0 -1.4243 0 -2.0 1e-06 
0.0 -1.4242 0 -2.0 1e-06 
0.0 -1.4241 0 -2.0 1e-06 
0.0 -1.424 0 -2.0 1e-06 
0.0 -1.4239 0 -2.0 1e-06 
0.0 -1.4238 0 -2.0 1e-06 
0.0 -1.4237 0 -2.0 1e-06 
0.0 -1.4236 0 -2.0 1e-06 
0.0 -1.4235 0 -2.0 1e-06 
0.0 -1.4234 0 -2.0 1e-06 
0.0 -1.4233 0 -2.0 1e-06 
0.0 -1.4232 0 -2.0 1e-06 
0.0 -1.4231 0 -2.0 1e-06 
0.0 -1.423 0 -2.0 1e-06 
0.0 -1.4229 0 -2.0 1e-06 
0.0 -1.4228 0 -2.0 1e-06 
0.0 -1.4227 0 -2.0 1e-06 
0.0 -1.4226 0 -2.0 1e-06 
0.0 -1.4225 0 -2.0 1e-06 
0.0 -1.4224 0 -2.0 1e-06 
0.0 -1.4223 0 -2.0 1e-06 
0.0 -1.4222 0 -2.0 1e-06 
0.0 -1.4221 0 -2.0 1e-06 
0.0 -1.422 0 -2.0 1e-06 
0.0 -1.4219 0 -2.0 1e-06 
0.0 -1.4218 0 -2.0 1e-06 
0.0 -1.4217 0 -2.0 1e-06 
0.0 -1.4216 0 -2.0 1e-06 
0.0 -1.4215 0 -2.0 1e-06 
0.0 -1.4214 0 -2.0 1e-06 
0.0 -1.4213 0 -2.0 1e-06 
0.0 -1.4212 0 -2.0 1e-06 
0.0 -1.4211 0 -2.0 1e-06 
0.0 -1.421 0 -2.0 1e-06 
0.0 -1.4209 0 -2.0 1e-06 
0.0 -1.4208 0 -2.0 1e-06 
0.0 -1.4207 0 -2.0 1e-06 
0.0 -1.4206 0 -2.0 1e-06 
0.0 -1.4205 0 -2.0 1e-06 
0.0 -1.4204 0 -2.0 1e-06 
0.0 -1.4203 0 -2.0 1e-06 
0.0 -1.4202 0 -2.0 1e-06 
0.0 -1.4201 0 -2.0 1e-06 
0.0 -1.42 0 -2.0 1e-06 
0.0 -1.4199 0 -2.0 1e-06 
0.0 -1.4198 0 -2.0 1e-06 
0.0 -1.4197 0 -2.0 1e-06 
0.0 -1.4196 0 -2.0 1e-06 
0.0 -1.4195 0 -2.0 1e-06 
0.0 -1.4194 0 -2.0 1e-06 
0.0 -1.4193 0 -2.0 1e-06 
0.0 -1.4192 0 -2.0 1e-06 
0.0 -1.4191 0 -2.0 1e-06 
0.0 -1.419 0 -2.0 1e-06 
0.0 -1.4189 0 -2.0 1e-06 
0.0 -1.4188 0 -2.0 1e-06 
0.0 -1.4187 0 -2.0 1e-06 
0.0 -1.4186 0 -2.0 1e-06 
0.0 -1.4185 0 -2.0 1e-06 
0.0 -1.4184 0 -2.0 1e-06 
0.0 -1.4183 0 -2.0 1e-06 
0.0 -1.4182 0 -2.0 1e-06 
0.0 -1.4181 0 -2.0 1e-06 
0.0 -1.418 0 -2.0 1e-06 
0.0 -1.4179 0 -2.0 1e-06 
0.0 -1.4178 0 -2.0 1e-06 
0.0 -1.4177 0 -2.0 1e-06 
0.0 -1.4176 0 -2.0 1e-06 
0.0 -1.4175 0 -2.0 1e-06 
0.0 -1.4174 0 -2.0 1e-06 
0.0 -1.4173 0 -2.0 1e-06 
0.0 -1.4172 0 -2.0 1e-06 
0.0 -1.4171 0 -2.0 1e-06 
0.0 -1.417 0 -2.0 1e-06 
0.0 -1.4169 0 -2.0 1e-06 
0.0 -1.4168 0 -2.0 1e-06 
0.0 -1.4167 0 -2.0 1e-06 
0.0 -1.4166 0 -2.0 1e-06 
0.0 -1.4165 0 -2.0 1e-06 
0.0 -1.4164 0 -2.0 1e-06 
0.0 -1.4163 0 -2.0 1e-06 
0.0 -1.4162 0 -2.0 1e-06 
0.0 -1.4161 0 -2.0 1e-06 
0.0 -1.416 0 -2.0 1e-06 
0.0 -1.4159 0 -2.0 1e-06 
0.0 -1.4158 0 -2.0 1e-06 
0.0 -1.4157 0 -2.0 1e-06 
0.0 -1.4156 0 -2.0 1e-06 
0.0 -1.4155 0 -2.0 1e-06 
0.0 -1.4154 0 -2.0 1e-06 
0.0 -1.4153 0 -2.0 1e-06 
0.0 -1.4152 0 -2.0 1e-06 
0.0 -1.4151 0 -2.0 1e-06 
0.0 -1.415 0 -2.0 1e-06 
0.0 -1.4149 0 -2.0 1e-06 
0.0 -1.4148 0 -2.0 1e-06 
0.0 -1.4147 0 -2.0 1e-06 
0.0 -1.4146 0 -2.0 1e-06 
0.0 -1.4145 0 -2.0 1e-06 
0.0 -1.4144 0 -2.0 1e-06 
0.0 -1.4143 0 -2.0 1e-06 
0.0 -1.4142 0 -2.0 1e-06 
0.0 -1.4141 0 -2.0 1e-06 
0.0 -1.414 0 -2.0 1e-06 
0.0 -1.4139 0 -2.0 1e-06 
0.0 -1.4138 0 -2.0 1e-06 
0.0 -1.4137 0 -2.0 1e-06 
0.0 -1.4136 0 -2.0 1e-06 
0.0 -1.4135 0 -2.0 1e-06 
0.0 -1.4134 0 -2.0 1e-06 
0.0 -1.4133 0 -2.0 1e-06 
0.0 -1.4132 0 -2.0 1e-06 
0.0 -1.4131 0 -2.0 1e-06 
0.0 -1.413 0 -2.0 1e-06 
0.0 -1.4129 0 -2.0 1e-06 
0.0 -1.4128 0 -2.0 1e-06 
0.0 -1.4127 0 -2.0 1e-06 
0.0 -1.4126 0 -2.0 1e-06 
0.0 -1.4125 0 -2.0 1e-06 
0.0 -1.4124 0 -2.0 1e-06 
0.0 -1.4123 0 -2.0 1e-06 
0.0 -1.4122 0 -2.0 1e-06 
0.0 -1.4121 0 -2.0 1e-06 
0.0 -1.412 0 -2.0 1e-06 
0.0 -1.4119 0 -2.0 1e-06 
0.0 -1.4118 0 -2.0 1e-06 
0.0 -1.4117 0 -2.0 1e-06 
0.0 -1.4116 0 -2.0 1e-06 
0.0 -1.4115 0 -2.0 1e-06 
0.0 -1.4114 0 -2.0 1e-06 
0.0 -1.4113 0 -2.0 1e-06 
0.0 -1.4112 0 -2.0 1e-06 
0.0 -1.4111 0 -2.0 1e-06 
0.0 -1.411 0 -2.0 1e-06 
0.0 -1.4109 0 -2.0 1e-06 
0.0 -1.4108 0 -2.0 1e-06 
0.0 -1.4107 0 -2.0 1e-06 
0.0 -1.4106 0 -2.0 1e-06 
0.0 -1.4105 0 -2.0 1e-06 
0.0 -1.4104 0 -2.0 1e-06 
0.0 -1.4103 0 -2.0 1e-06 
0.0 -1.4102 0 -2.0 1e-06 
0.0 -1.4101 0 -2.0 1e-06 
0.0 -1.41 0 -2.0 1e-06 
0.0 -1.4099 0 -2.0 1e-06 
0.0 -1.4098 0 -2.0 1e-06 
0.0 -1.4097 0 -2.0 1e-06 
0.0 -1.4096 0 -2.0 1e-06 
0.0 -1.4095 0 -2.0 1e-06 
0.0 -1.4094 0 -2.0 1e-06 
0.0 -1.4093 0 -2.0 1e-06 
0.0 -1.4092 0 -2.0 1e-06 
0.0 -1.4091 0 -2.0 1e-06 
0.0 -1.409 0 -2.0 1e-06 
0.0 -1.4089 0 -2.0 1e-06 
0.0 -1.4088 0 -2.0 1e-06 
0.0 -1.4087 0 -2.0 1e-06 
0.0 -1.4086 0 -2.0 1e-06 
0.0 -1.4085 0 -2.0 1e-06 
0.0 -1.4084 0 -2.0 1e-06 
0.0 -1.4083 0 -2.0 1e-06 
0.0 -1.4082 0 -2.0 1e-06 
0.0 -1.4081 0 -2.0 1e-06 
0.0 -1.408 0 -2.0 1e-06 
0.0 -1.4079 0 -2.0 1e-06 
0.0 -1.4078 0 -2.0 1e-06 
0.0 -1.4077 0 -2.0 1e-06 
0.0 -1.4076 0 -2.0 1e-06 
0.0 -1.4075 0 -2.0 1e-06 
0.0 -1.4074 0 -2.0 1e-06 
0.0 -1.4073 0 -2.0 1e-06 
0.0 -1.4072 0 -2.0 1e-06 
0.0 -1.4071 0 -2.0 1e-06 
0.0 -1.407 0 -2.0 1e-06 
0.0 -1.4069 0 -2.0 1e-06 
0.0 -1.4068 0 -2.0 1e-06 
0.0 -1.4067 0 -2.0 1e-06 
0.0 -1.4066 0 -2.0 1e-06 
0.0 -1.4065 0 -2.0 1e-06 
0.0 -1.4064 0 -2.0 1e-06 
0.0 -1.4063 0 -2.0 1e-06 
0.0 -1.4062 0 -2.0 1e-06 
0.0 -1.4061 0 -2.0 1e-06 
0.0 -1.406 0 -2.0 1e-06 
0.0 -1.4059 0 -2.0 1e-06 
0.0 -1.4058 0 -2.0 1e-06 
0.0 -1.4057 0 -2.0 1e-06 
0.0 -1.4056 0 -2.0 1e-06 
0.0 -1.4055 0 -2.0 1e-06 
0.0 -1.4054 0 -2.0 1e-06 
0.0 -1.4053 0 -2.0 1e-06 
0.0 -1.4052 0 -2.0 1e-06 
0.0 -1.4051 0 -2.0 1e-06 
0.0 -1.405 0 -2.0 1e-06 
0.0 -1.4049 0 -2.0 1e-06 
0.0 -1.4048 0 -2.0 1e-06 
0.0 -1.4047 0 -2.0 1e-06 
0.0 -1.4046 0 -2.0 1e-06 
0.0 -1.4045 0 -2.0 1e-06 
0.0 -1.4044 0 -2.0 1e-06 
0.0 -1.4043 0 -2.0 1e-06 
0.0 -1.4042 0 -2.0 1e-06 
0.0 -1.4041 0 -2.0 1e-06 
0.0 -1.404 0 -2.0 1e-06 
0.0 -1.4039 0 -2.0 1e-06 
0.0 -1.4038 0 -2.0 1e-06 
0.0 -1.4037 0 -2.0 1e-06 
0.0 -1.4036 0 -2.0 1e-06 
0.0 -1.4035 0 -2.0 1e-06 
0.0 -1.4034 0 -2.0 1e-06 
0.0 -1.4033 0 -2.0 1e-06 
0.0 -1.4032 0 -2.0 1e-06 
0.0 -1.4031 0 -2.0 1e-06 
0.0 -1.403 0 -2.0 1e-06 
0.0 -1.4029 0 -2.0 1e-06 
0.0 -1.4028 0 -2.0 1e-06 
0.0 -1.4027 0 -2.0 1e-06 
0.0 -1.4026 0 -2.0 1e-06 
0.0 -1.4025 0 -2.0 1e-06 
0.0 -1.4024 0 -2.0 1e-06 
0.0 -1.4023 0 -2.0 1e-06 
0.0 -1.4022 0 -2.0 1e-06 
0.0 -1.4021 0 -2.0 1e-06 
0.0 -1.402 0 -2.0 1e-06 
0.0 -1.4019 0 -2.0 1e-06 
0.0 -1.4018 0 -2.0 1e-06 
0.0 -1.4017 0 -2.0 1e-06 
0.0 -1.4016 0 -2.0 1e-06 
0.0 -1.4015 0 -2.0 1e-06 
0.0 -1.4014 0 -2.0 1e-06 
0.0 -1.4013 0 -2.0 1e-06 
0.0 -1.4012 0 -2.0 1e-06 
0.0 -1.4011 0 -2.0 1e-06 
0.0 -1.401 0 -2.0 1e-06 
0.0 -1.4009 0 -2.0 1e-06 
0.0 -1.4008 0 -2.0 1e-06 
0.0 -1.4007 0 -2.0 1e-06 
0.0 -1.4006 0 -2.0 1e-06 
0.0 -1.4005 0 -2.0 1e-06 
0.0 -1.4004 0 -2.0 1e-06 
0.0 -1.4003 0 -2.0 1e-06 
0.0 -1.4002 0 -2.0 1e-06 
0.0 -1.4001 0 -2.0 1e-06 
0.0 -1.4 0 -2.0 1e-06 
0.0 -1.3999 0 -2.0 1e-06 
0.0 -1.3998 0 -2.0 1e-06 
0.0 -1.3997 0 -2.0 1e-06 
0.0 -1.3996 0 -2.0 1e-06 
0.0 -1.3995 0 -2.0 1e-06 
0.0 -1.3994 0 -2.0 1e-06 
0.0 -1.3993 0 -2.0 1e-06 
0.0 -1.3992 0 -2.0 1e-06 
0.0 -1.3991 0 -2.0 1e-06 
0.0 -1.399 0 -2.0 1e-06 
0.0 -1.3989 0 -2.0 1e-06 
0.0 -1.3988 0 -2.0 1e-06 
0.0 -1.3987 0 -2.0 1e-06 
0.0 -1.3986 0 -2.0 1e-06 
0.0 -1.3985 0 -2.0 1e-06 
0.0 -1.3984 0 -2.0 1e-06 
0.0 -1.3983 0 -2.0 1e-06 
0.0 -1.3982 0 -2.0 1e-06 
0.0 -1.3981 0 -2.0 1e-06 
0.0 -1.398 0 -2.0 1e-06 
0.0 -1.3979 0 -2.0 1e-06 
0.0 -1.3978 0 -2.0 1e-06 
0.0 -1.3977 0 -2.0 1e-06 
0.0 -1.3976 0 -2.0 1e-06 
0.0 -1.3975 0 -2.0 1e-06 
0.0 -1.3974 0 -2.0 1e-06 
0.0 -1.3973 0 -2.0 1e-06 
0.0 -1.3972 0 -2.0 1e-06 
0.0 -1.3971 0 -2.0 1e-06 
0.0 -1.397 0 -2.0 1e-06 
0.0 -1.3969 0 -2.0 1e-06 
0.0 -1.3968 0 -2.0 1e-06 
0.0 -1.3967 0 -2.0 1e-06 
0.0 -1.3966 0 -2.0 1e-06 
0.0 -1.3965 0 -2.0 1e-06 
0.0 -1.3964 0 -2.0 1e-06 
0.0 -1.3963 0 -2.0 1e-06 
0.0 -1.3962 0 -2.0 1e-06 
0.0 -1.3961 0 -2.0 1e-06 
0.0 -1.396 0 -2.0 1e-06 
0.0 -1.3959 0 -2.0 1e-06 
0.0 -1.3958 0 -2.0 1e-06 
0.0 -1.3957 0 -2.0 1e-06 
0.0 -1.3956 0 -2.0 1e-06 
0.0 -1.3955 0 -2.0 1e-06 
0.0 -1.3954 0 -2.0 1e-06 
0.0 -1.3953 0 -2.0 1e-06 
0.0 -1.3952 0 -2.0 1e-06 
0.0 -1.3951 0 -2.0 1e-06 
0.0 -1.395 0 -2.0 1e-06 
0.0 -1.3949 0 -2.0 1e-06 
0.0 -1.3948 0 -2.0 1e-06 
0.0 -1.3947 0 -2.0 1e-06 
0.0 -1.3946 0 -2.0 1e-06 
0.0 -1.3945 0 -2.0 1e-06 
0.0 -1.3944 0 -2.0 1e-06 
0.0 -1.3943 0 -2.0 1e-06 
0.0 -1.3942 0 -2.0 1e-06 
0.0 -1.3941 0 -2.0 1e-06 
0.0 -1.394 0 -2.0 1e-06 
0.0 -1.3939 0 -2.0 1e-06 
0.0 -1.3938 0 -2.0 1e-06 
0.0 -1.3937 0 -2.0 1e-06 
0.0 -1.3936 0 -2.0 1e-06 
0.0 -1.3935 0 -2.0 1e-06 
0.0 -1.3934 0 -2.0 1e-06 
0.0 -1.3933 0 -2.0 1e-06 
0.0 -1.3932 0 -2.0 1e-06 
0.0 -1.3931 0 -2.0 1e-06 
0.0 -1.393 0 -2.0 1e-06 
0.0 -1.3929 0 -2.0 1e-06 
0.0 -1.3928 0 -2.0 1e-06 
0.0 -1.3927 0 -2.0 1e-06 
0.0 -1.3926 0 -2.0 1e-06 
0.0 -1.3925 0 -2.0 1e-06 
0.0 -1.3924 0 -2.0 1e-06 
0.0 -1.3923 0 -2.0 1e-06 
0.0 -1.3922 0 -2.0 1e-06 
0.0 -1.3921 0 -2.0 1e-06 
0.0 -1.392 0 -2.0 1e-06 
0.0 -1.3919 0 -2.0 1e-06 
0.0 -1.3918 0 -2.0 1e-06 
0.0 -1.3917 0 -2.0 1e-06 
0.0 -1.3916 0 -2.0 1e-06 
0.0 -1.3915 0 -2.0 1e-06 
0.0 -1.3914 0 -2.0 1e-06 
0.0 -1.3913 0 -2.0 1e-06 
0.0 -1.3912 0 -2.0 1e-06 
0.0 -1.3911 0 -2.0 1e-06 
0.0 -1.391 0 -2.0 1e-06 
0.0 -1.3909 0 -2.0 1e-06 
0.0 -1.3908 0 -2.0 1e-06 
0.0 -1.3907 0 -2.0 1e-06 
0.0 -1.3906 0 -2.0 1e-06 
0.0 -1.3905 0 -2.0 1e-06 
0.0 -1.3904 0 -2.0 1e-06 
0.0 -1.3903 0 -2.0 1e-06 
0.0 -1.3902 0 -2.0 1e-06 
0.0 -1.3901 0 -2.0 1e-06 
0.0 -1.39 0 -2.0 1e-06 
0.0 -1.3899 0 -2.0 1e-06 
0.0 -1.3898 0 -2.0 1e-06 
0.0 -1.3897 0 -2.0 1e-06 
0.0 -1.3896 0 -2.0 1e-06 
0.0 -1.3895 0 -2.0 1e-06 
0.0 -1.3894 0 -2.0 1e-06 
0.0 -1.3893 0 -2.0 1e-06 
0.0 -1.3892 0 -2.0 1e-06 
0.0 -1.3891 0 -2.0 1e-06 
0.0 -1.389 0 -2.0 1e-06 
0.0 -1.3889 0 -2.0 1e-06 
0.0 -1.3888 0 -2.0 1e-06 
0.0 -1.3887 0 -2.0 1e-06 
0.0 -1.3886 0 -2.0 1e-06 
0.0 -1.3885 0 -2.0 1e-06 
0.0 -1.3884 0 -2.0 1e-06 
0.0 -1.3883 0 -2.0 1e-06 
0.0 -1.3882 0 -2.0 1e-06 
0.0 -1.3881 0 -2.0 1e-06 
0.0 -1.388 0 -2.0 1e-06 
0.0 -1.3879 0 -2.0 1e-06 
0.0 -1.3878 0 -2.0 1e-06 
0.0 -1.3877 0 -2.0 1e-06 
0.0 -1.3876 0 -2.0 1e-06 
0.0 -1.3875 0 -2.0 1e-06 
0.0 -1.3874 0 -2.0 1e-06 
0.0 -1.3873 0 -2.0 1e-06 
0.0 -1.3872 0 -2.0 1e-06 
0.0 -1.3871 0 -2.0 1e-06 
0.0 -1.387 0 -2.0 1e-06 
0.0 -1.3869 0 -2.0 1e-06 
0.0 -1.3868 0 -2.0 1e-06 
0.0 -1.3867 0 -2.0 1e-06 
0.0 -1.3866 0 -2.0 1e-06 
0.0 -1.3865 0 -2.0 1e-06 
0.0 -1.3864 0 -2.0 1e-06 
0.0 -1.3863 0 -2.0 1e-06 
0.0 -1.3862 0 -2.0 1e-06 
0.0 -1.3861 0 -2.0 1e-06 
0.0 -1.386 0 -2.0 1e-06 
0.0 -1.3859 0 -2.0 1e-06 
0.0 -1.3858 0 -2.0 1e-06 
0.0 -1.3857 0 -2.0 1e-06 
0.0 -1.3856 0 -2.0 1e-06 
0.0 -1.3855 0 -2.0 1e-06 
0.0 -1.3854 0 -2.0 1e-06 
0.0 -1.3853 0 -2.0 1e-06 
0.0 -1.3852 0 -2.0 1e-06 
0.0 -1.3851 0 -2.0 1e-06 
0.0 -1.385 0 -2.0 1e-06 
0.0 -1.3849 0 -2.0 1e-06 
0.0 -1.3848 0 -2.0 1e-06 
0.0 -1.3847 0 -2.0 1e-06 
0.0 -1.3846 0 -2.0 1e-06 
0.0 -1.3845 0 -2.0 1e-06 
0.0 -1.3844 0 -2.0 1e-06 
0.0 -1.3843 0 -2.0 1e-06 
0.0 -1.3842 0 -2.0 1e-06 
0.0 -1.3841 0 -2.0 1e-06 
0.0 -1.384 0 -2.0 1e-06 
0.0 -1.3839 0 -2.0 1e-06 
0.0 -1.3838 0 -2.0 1e-06 
0.0 -1.3837 0 -2.0 1e-06 
0.0 -1.3836 0 -2.0 1e-06 
0.0 -1.3835 0 -2.0 1e-06 
0.0 -1.3834 0 -2.0 1e-06 
0.0 -1.3833 0 -2.0 1e-06 
0.0 -1.3832 0 -2.0 1e-06 
0.0 -1.3831 0 -2.0 1e-06 
0.0 -1.383 0 -2.0 1e-06 
0.0 -1.3829 0 -2.0 1e-06 
0.0 -1.3828 0 -2.0 1e-06 
0.0 -1.3827 0 -2.0 1e-06 
0.0 -1.3826 0 -2.0 1e-06 
0.0 -1.3825 0 -2.0 1e-06 
0.0 -1.3824 0 -2.0 1e-06 
0.0 -1.3823 0 -2.0 1e-06 
0.0 -1.3822 0 -2.0 1e-06 
0.0 -1.3821 0 -2.0 1e-06 
0.0 -1.382 0 -2.0 1e-06 
0.0 -1.3819 0 -2.0 1e-06 
0.0 -1.3818 0 -2.0 1e-06 
0.0 -1.3817 0 -2.0 1e-06 
0.0 -1.3816 0 -2.0 1e-06 
0.0 -1.3815 0 -2.0 1e-06 
0.0 -1.3814 0 -2.0 1e-06 
0.0 -1.3813 0 -2.0 1e-06 
0.0 -1.3812 0 -2.0 1e-06 
0.0 -1.3811 0 -2.0 1e-06 
0.0 -1.381 0 -2.0 1e-06 
0.0 -1.3809 0 -2.0 1e-06 
0.0 -1.3808 0 -2.0 1e-06 
0.0 -1.3807 0 -2.0 1e-06 
0.0 -1.3806 0 -2.0 1e-06 
0.0 -1.3805 0 -2.0 1e-06 
0.0 -1.3804 0 -2.0 1e-06 
0.0 -1.3803 0 -2.0 1e-06 
0.0 -1.3802 0 -2.0 1e-06 
0.0 -1.3801 0 -2.0 1e-06 
0.0 -1.38 0 -2.0 1e-06 
0.0 -1.3799 0 -2.0 1e-06 
0.0 -1.3798 0 -2.0 1e-06 
0.0 -1.3797 0 -2.0 1e-06 
0.0 -1.3796 0 -2.0 1e-06 
0.0 -1.3795 0 -2.0 1e-06 
0.0 -1.3794 0 -2.0 1e-06 
0.0 -1.3793 0 -2.0 1e-06 
0.0 -1.3792 0 -2.0 1e-06 
0.0 -1.3791 0 -2.0 1e-06 
0.0 -1.379 0 -2.0 1e-06 
0.0 -1.3789 0 -2.0 1e-06 
0.0 -1.3788 0 -2.0 1e-06 
0.0 -1.3787 0 -2.0 1e-06 
0.0 -1.3786 0 -2.0 1e-06 
0.0 -1.3785 0 -2.0 1e-06 
0.0 -1.3784 0 -2.0 1e-06 
0.0 -1.3783 0 -2.0 1e-06 
0.0 -1.3782 0 -2.0 1e-06 
0.0 -1.3781 0 -2.0 1e-06 
0.0 -1.378 0 -2.0 1e-06 
0.0 -1.3779 0 -2.0 1e-06 
0.0 -1.3778 0 -2.0 1e-06 
0.0 -1.3777 0 -2.0 1e-06 
0.0 -1.3776 0 -2.0 1e-06 
0.0 -1.3775 0 -2.0 1e-06 
0.0 -1.3774 0 -2.0 1e-06 
0.0 -1.3773 0 -2.0 1e-06 
0.0 -1.3772 0 -2.0 1e-06 
0.0 -1.3771 0 -2.0 1e-06 
0.0 -1.377 0 -2.0 1e-06 
0.0 -1.3769 0 -2.0 1e-06 
0.0 -1.3768 0 -2.0 1e-06 
0.0 -1.3767 0 -2.0 1e-06 
0.0 -1.3766 0 -2.0 1e-06 
0.0 -1.3765 0 -2.0 1e-06 
0.0 -1.3764 0 -2.0 1e-06 
0.0 -1.3763 0 -2.0 1e-06 
0.0 -1.3762 0 -2.0 1e-06 
0.0 -1.3761 0 -2.0 1e-06 
0.0 -1.376 0 -2.0 1e-06 
0.0 -1.3759 0 -2.0 1e-06 
0.0 -1.3758 0 -2.0 1e-06 
0.0 -1.3757 0 -2.0 1e-06 
0.0 -1.3756 0 -2.0 1e-06 
0.0 -1.3755 0 -2.0 1e-06 
0.0 -1.3754 0 -2.0 1e-06 
0.0 -1.3753 0 -2.0 1e-06 
0.0 -1.3752 0 -2.0 1e-06 
0.0 -1.3751 0 -2.0 1e-06 
0.0 -1.375 0 -2.0 1e-06 
0.0 -1.3749 0 -2.0 1e-06 
0.0 -1.3748 0 -2.0 1e-06 
0.0 -1.3747 0 -2.0 1e-06 
0.0 -1.3746 0 -2.0 1e-06 
0.0 -1.3745 0 -2.0 1e-06 
0.0 -1.3744 0 -2.0 1e-06 
0.0 -1.3743 0 -2.0 1e-06 
0.0 -1.3742 0 -2.0 1e-06 
0.0 -1.3741 0 -2.0 1e-06 
0.0 -1.374 0 -2.0 1e-06 
0.0 -1.3739 0 -2.0 1e-06 
0.0 -1.3738 0 -2.0 1e-06 
0.0 -1.3737 0 -2.0 1e-06 
0.0 -1.3736 0 -2.0 1e-06 
0.0 -1.3735 0 -2.0 1e-06 
0.0 -1.3734 0 -2.0 1e-06 
0.0 -1.3733 0 -2.0 1e-06 
0.0 -1.3732 0 -2.0 1e-06 
0.0 -1.3731 0 -2.0 1e-06 
0.0 -1.373 0 -2.0 1e-06 
0.0 -1.3729 0 -2.0 1e-06 
0.0 -1.3728 0 -2.0 1e-06 
0.0 -1.3727 0 -2.0 1e-06 
0.0 -1.3726 0 -2.0 1e-06 
0.0 -1.3725 0 -2.0 1e-06 
0.0 -1.3724 0 -2.0 1e-06 
0.0 -1.3723 0 -2.0 1e-06 
0.0 -1.3722 0 -2.0 1e-06 
0.0 -1.3721 0 -2.0 1e-06 
0.0 -1.372 0 -2.0 1e-06 
0.0 -1.3719 0 -2.0 1e-06 
0.0 -1.3718 0 -2.0 1e-06 
0.0 -1.3717 0 -2.0 1e-06 
0.0 -1.3716 0 -2.0 1e-06 
0.0 -1.3715 0 -2.0 1e-06 
0.0 -1.3714 0 -2.0 1e-06 
0.0 -1.3713 0 -2.0 1e-06 
0.0 -1.3712 0 -2.0 1e-06 
0.0 -1.3711 0 -2.0 1e-06 
0.0 -1.371 0 -2.0 1e-06 
0.0 -1.3709 0 -2.0 1e-06 
0.0 -1.3708 0 -2.0 1e-06 
0.0 -1.3707 0 -2.0 1e-06 
0.0 -1.3706 0 -2.0 1e-06 
0.0 -1.3705 0 -2.0 1e-06 
0.0 -1.3704 0 -2.0 1e-06 
0.0 -1.3703 0 -2.0 1e-06 
0.0 -1.3702 0 -2.0 1e-06 
0.0 -1.3701 0 -2.0 1e-06 
0.0 -1.37 0 -2.0 1e-06 
0.0 -1.3699 0 -2.0 1e-06 
0.0 -1.3698 0 -2.0 1e-06 
0.0 -1.3697 0 -2.0 1e-06 
0.0 -1.3696 0 -2.0 1e-06 
0.0 -1.3695 0 -2.0 1e-06 
0.0 -1.3694 0 -2.0 1e-06 
0.0 -1.3693 0 -2.0 1e-06 
0.0 -1.3692 0 -2.0 1e-06 
0.0 -1.3691 0 -2.0 1e-06 
0.0 -1.369 0 -2.0 1e-06 
0.0 -1.3689 0 -2.0 1e-06 
0.0 -1.3688 0 -2.0 1e-06 
0.0 -1.3687 0 -2.0 1e-06 
0.0 -1.3686 0 -2.0 1e-06 
0.0 -1.3685 0 -2.0 1e-06 
0.0 -1.3684 0 -2.0 1e-06 
0.0 -1.3683 0 -2.0 1e-06 
0.0 -1.3682 0 -2.0 1e-06 
0.0 -1.3681 0 -2.0 1e-06 
0.0 -1.368 0 -2.0 1e-06 
0.0 -1.3679 0 -2.0 1e-06 
0.0 -1.3678 0 -2.0 1e-06 
0.0 -1.3677 0 -2.0 1e-06 
0.0 -1.3676 0 -2.0 1e-06 
0.0 -1.3675 0 -2.0 1e-06 
0.0 -1.3674 0 -2.0 1e-06 
0.0 -1.3673 0 -2.0 1e-06 
0.0 -1.3672 0 -2.0 1e-06 
0.0 -1.3671 0 -2.0 1e-06 
0.0 -1.367 0 -2.0 1e-06 
0.0 -1.3669 0 -2.0 1e-06 
0.0 -1.3668 0 -2.0 1e-06 
0.0 -1.3667 0 -2.0 1e-06 
0.0 -1.3666 0 -2.0 1e-06 
0.0 -1.3665 0 -2.0 1e-06 
0.0 -1.3664 0 -2.0 1e-06 
0.0 -1.3663 0 -2.0 1e-06 
0.0 -1.3662 0 -2.0 1e-06 
0.0 -1.3661 0 -2.0 1e-06 
0.0 -1.366 0 -2.0 1e-06 
0.0 -1.3659 0 -2.0 1e-06 
0.0 -1.3658 0 -2.0 1e-06 
0.0 -1.3657 0 -2.0 1e-06 
0.0 -1.3656 0 -2.0 1e-06 
0.0 -1.3655 0 -2.0 1e-06 
0.0 -1.3654 0 -2.0 1e-06 
0.0 -1.3653 0 -2.0 1e-06 
0.0 -1.3652 0 -2.0 1e-06 
0.0 -1.3651 0 -2.0 1e-06 
0.0 -1.365 0 -2.0 1e-06 
0.0 -1.3649 0 -2.0 1e-06 
0.0 -1.3648 0 -2.0 1e-06 
0.0 -1.3647 0 -2.0 1e-06 
0.0 -1.3646 0 -2.0 1e-06 
0.0 -1.3645 0 -2.0 1e-06 
0.0 -1.3644 0 -2.0 1e-06 
0.0 -1.3643 0 -2.0 1e-06 
0.0 -1.3642 0 -2.0 1e-06 
0.0 -1.3641 0 -2.0 1e-06 
0.0 -1.364 0 -2.0 1e-06 
0.0 -1.3639 0 -2.0 1e-06 
0.0 -1.3638 0 -2.0 1e-06 
0.0 -1.3637 0 -2.0 1e-06 
0.0 -1.3636 0 -2.0 1e-06 
0.0 -1.3635 0 -2.0 1e-06 
0.0 -1.3634 0 -2.0 1e-06 
0.0 -1.3633 0 -2.0 1e-06 
0.0 -1.3632 0 -2.0 1e-06 
0.0 -1.3631 0 -2.0 1e-06 
0.0 -1.363 0 -2.0 1e-06 
0.0 -1.3629 0 -2.0 1e-06 
0.0 -1.3628 0 -2.0 1e-06 
0.0 -1.3627 0 -2.0 1e-06 
0.0 -1.3626 0 -2.0 1e-06 
0.0 -1.3625 0 -2.0 1e-06 
0.0 -1.3624 0 -2.0 1e-06 
0.0 -1.3623 0 -2.0 1e-06 
0.0 -1.3622 0 -2.0 1e-06 
0.0 -1.3621 0 -2.0 1e-06 
0.0 -1.362 0 -2.0 1e-06 
0.0 -1.3619 0 -2.0 1e-06 
0.0 -1.3618 0 -2.0 1e-06 
0.0 -1.3617 0 -2.0 1e-06 
0.0 -1.3616 0 -2.0 1e-06 
0.0 -1.3615 0 -2.0 1e-06 
0.0 -1.3614 0 -2.0 1e-06 
0.0 -1.3613 0 -2.0 1e-06 
0.0 -1.3612 0 -2.0 1e-06 
0.0 -1.3611 0 -2.0 1e-06 
0.0 -1.361 0 -2.0 1e-06 
0.0 -1.3609 0 -2.0 1e-06 
0.0 -1.3608 0 -2.0 1e-06 
0.0 -1.3607 0 -2.0 1e-06 
0.0 -1.3606 0 -2.0 1e-06 
0.0 -1.3605 0 -2.0 1e-06 
0.0 -1.3604 0 -2.0 1e-06 
0.0 -1.3603 0 -2.0 1e-06 
0.0 -1.3602 0 -2.0 1e-06 
0.0 -1.3601 0 -2.0 1e-06 
0.0 -1.36 0 -2.0 1e-06 
0.0 -1.3599 0 -2.0 1e-06 
0.0 -1.3598 0 -2.0 1e-06 
0.0 -1.3597 0 -2.0 1e-06 
0.0 -1.3596 0 -2.0 1e-06 
0.0 -1.3595 0 -2.0 1e-06 
0.0 -1.3594 0 -2.0 1e-06 
0.0 -1.3593 0 -2.0 1e-06 
0.0 -1.3592 0 -2.0 1e-06 
0.0 -1.3591 0 -2.0 1e-06 
0.0 -1.359 0 -2.0 1e-06 
0.0 -1.3589 0 -2.0 1e-06 
0.0 -1.3588 0 -2.0 1e-06 
0.0 -1.3587 0 -2.0 1e-06 
0.0 -1.3586 0 -2.0 1e-06 
0.0 -1.3585 0 -2.0 1e-06 
0.0 -1.3584 0 -2.0 1e-06 
0.0 -1.3583 0 -2.0 1e-06 
0.0 -1.3582 0 -2.0 1e-06 
0.0 -1.3581 0 -2.0 1e-06 
0.0 -1.358 0 -2.0 1e-06 
0.0 -1.3579 0 -2.0 1e-06 
0.0 -1.3578 0 -2.0 1e-06 
0.0 -1.3577 0 -2.0 1e-06 
0.0 -1.3576 0 -2.0 1e-06 
0.0 -1.3575 0 -2.0 1e-06 
0.0 -1.3574 0 -2.0 1e-06 
0.0 -1.3573 0 -2.0 1e-06 
0.0 -1.3572 0 -2.0 1e-06 
0.0 -1.3571 0 -2.0 1e-06 
0.0 -1.357 0 -2.0 1e-06 
0.0 -1.3569 0 -2.0 1e-06 
0.0 -1.3568 0 -2.0 1e-06 
0.0 -1.3567 0 -2.0 1e-06 
0.0 -1.3566 0 -2.0 1e-06 
0.0 -1.3565 0 -2.0 1e-06 
0.0 -1.3564 0 -2.0 1e-06 
0.0 -1.3563 0 -2.0 1e-06 
0.0 -1.3562 0 -2.0 1e-06 
0.0 -1.3561 0 -2.0 1e-06 
0.0 -1.356 0 -2.0 1e-06 
0.0 -1.3559 0 -2.0 1e-06 
0.0 -1.3558 0 -2.0 1e-06 
0.0 -1.3557 0 -2.0 1e-06 
0.0 -1.3556 0 -2.0 1e-06 
0.0 -1.3555 0 -2.0 1e-06 
0.0 -1.3554 0 -2.0 1e-06 
0.0 -1.3553 0 -2.0 1e-06 
0.0 -1.3552 0 -2.0 1e-06 
0.0 -1.3551 0 -2.0 1e-06 
0.0 -1.355 0 -2.0 1e-06 
0.0 -1.3549 0 -2.0 1e-06 
0.0 -1.3548 0 -2.0 1e-06 
0.0 -1.3547 0 -2.0 1e-06 
0.0 -1.3546 0 -2.0 1e-06 
0.0 -1.3545 0 -2.0 1e-06 
0.0 -1.3544 0 -2.0 1e-06 
0.0 -1.3543 0 -2.0 1e-06 
0.0 -1.3542 0 -2.0 1e-06 
0.0 -1.3541 0 -2.0 1e-06 
0.0 -1.354 0 -2.0 1e-06 
0.0 -1.3539 0 -2.0 1e-06 
0.0 -1.3538 0 -2.0 1e-06 
0.0 -1.3537 0 -2.0 1e-06 
0.0 -1.3536 0 -2.0 1e-06 
0.0 -1.3535 0 -2.0 1e-06 
0.0 -1.3534 0 -2.0 1e-06 
0.0 -1.3533 0 -2.0 1e-06 
0.0 -1.3532 0 -2.0 1e-06 
0.0 -1.3531 0 -2.0 1e-06 
0.0 -1.353 0 -2.0 1e-06 
0.0 -1.3529 0 -2.0 1e-06 
0.0 -1.3528 0 -2.0 1e-06 
0.0 -1.3527 0 -2.0 1e-06 
0.0 -1.3526 0 -2.0 1e-06 
0.0 -1.3525 0 -2.0 1e-06 
0.0 -1.3524 0 -2.0 1e-06 
0.0 -1.3523 0 -2.0 1e-06 
0.0 -1.3522 0 -2.0 1e-06 
0.0 -1.3521 0 -2.0 1e-06 
0.0 -1.352 0 -2.0 1e-06 
0.0 -1.3519 0 -2.0 1e-06 
0.0 -1.3518 0 -2.0 1e-06 
0.0 -1.3517 0 -2.0 1e-06 
0.0 -1.3516 0 -2.0 1e-06 
0.0 -1.3515 0 -2.0 1e-06 
0.0 -1.3514 0 -2.0 1e-06 
0.0 -1.3513 0 -2.0 1e-06 
0.0 -1.3512 0 -2.0 1e-06 
0.0 -1.3511 0 -2.0 1e-06 
0.0 -1.351 0 -2.0 1e-06 
0.0 -1.3509 0 -2.0 1e-06 
0.0 -1.3508 0 -2.0 1e-06 
0.0 -1.3507 0 -2.0 1e-06 
0.0 -1.3506 0 -2.0 1e-06 
0.0 -1.3505 0 -2.0 1e-06 
0.0 -1.3504 0 -2.0 1e-06 
0.0 -1.3503 0 -2.0 1e-06 
0.0 -1.3502 0 -2.0 1e-06 
0.0 -1.3501 0 -2.0 1e-06 
0.0 -1.35 0 -2.0 1e-06 
0.0 -1.3499 0 -2.0 1e-06 
0.0 -1.3498 0 -2.0 1e-06 
0.0 -1.3497 0 -2.0 1e-06 
0.0 -1.3496 0 -2.0 1e-06 
0.0 -1.3495 0 -2.0 1e-06 
0.0 -1.3494 0 -2.0 1e-06 
0.0 -1.3493 0 -2.0 1e-06 
0.0 -1.3492 0 -2.0 1e-06 
0.0 -1.3491 0 -2.0 1e-06 
0.0 -1.349 0 -2.0 1e-06 
0.0 -1.3489 0 -2.0 1e-06 
0.0 -1.3488 0 -2.0 1e-06 
0.0 -1.3487 0 -2.0 1e-06 
0.0 -1.3486 0 -2.0 1e-06 
0.0 -1.3485 0 -2.0 1e-06 
0.0 -1.3484 0 -2.0 1e-06 
0.0 -1.3483 0 -2.0 1e-06 
0.0 -1.3482 0 -2.0 1e-06 
0.0 -1.3481 0 -2.0 1e-06 
0.0 -1.348 0 -2.0 1e-06 
0.0 -1.3479 0 -2.0 1e-06 
0.0 -1.3478 0 -2.0 1e-06 
0.0 -1.3477 0 -2.0 1e-06 
0.0 -1.3476 0 -2.0 1e-06 
0.0 -1.3475 0 -2.0 1e-06 
0.0 -1.3474 0 -2.0 1e-06 
0.0 -1.3473 0 -2.0 1e-06 
0.0 -1.3472 0 -2.0 1e-06 
0.0 -1.3471 0 -2.0 1e-06 
0.0 -1.347 0 -2.0 1e-06 
0.0 -1.3469 0 -2.0 1e-06 
0.0 -1.3468 0 -2.0 1e-06 
0.0 -1.3467 0 -2.0 1e-06 
0.0 -1.3466 0 -2.0 1e-06 
0.0 -1.3465 0 -2.0 1e-06 
0.0 -1.3464 0 -2.0 1e-06 
0.0 -1.3463 0 -2.0 1e-06 
0.0 -1.3462 0 -2.0 1e-06 
0.0 -1.3461 0 -2.0 1e-06 
0.0 -1.346 0 -2.0 1e-06 
0.0 -1.3459 0 -2.0 1e-06 
0.0 -1.3458 0 -2.0 1e-06 
0.0 -1.3457 0 -2.0 1e-06 
0.0 -1.3456 0 -2.0 1e-06 
0.0 -1.3455 0 -2.0 1e-06 
0.0 -1.3454 0 -2.0 1e-06 
0.0 -1.3453 0 -2.0 1e-06 
0.0 -1.3452 0 -2.0 1e-06 
0.0 -1.3451 0 -2.0 1e-06 
0.0 -1.345 0 -2.0 1e-06 
0.0 -1.3449 0 -2.0 1e-06 
0.0 -1.3448 0 -2.0 1e-06 
0.0 -1.3447 0 -2.0 1e-06 
0.0 -1.3446 0 -2.0 1e-06 
0.0 -1.3445 0 -2.0 1e-06 
0.0 -1.3444 0 -2.0 1e-06 
0.0 -1.3443 0 -2.0 1e-06 
0.0 -1.3442 0 -2.0 1e-06 
0.0 -1.3441 0 -2.0 1e-06 
0.0 -1.344 0 -2.0 1e-06 
0.0 -1.3439 0 -2.0 1e-06 
0.0 -1.3438 0 -2.0 1e-06 
0.0 -1.3437 0 -2.0 1e-06 
0.0 -1.3436 0 -2.0 1e-06 
0.0 -1.3435 0 -2.0 1e-06 
0.0 -1.3434 0 -2.0 1e-06 
0.0 -1.3433 0 -2.0 1e-06 
0.0 -1.3432 0 -2.0 1e-06 
0.0 -1.3431 0 -2.0 1e-06 
0.0 -1.343 0 -2.0 1e-06 
0.0 -1.3429 0 -2.0 1e-06 
0.0 -1.3428 0 -2.0 1e-06 
0.0 -1.3427 0 -2.0 1e-06 
0.0 -1.3426 0 -2.0 1e-06 
0.0 -1.3425 0 -2.0 1e-06 
0.0 -1.3424 0 -2.0 1e-06 
0.0 -1.3423 0 -2.0 1e-06 
0.0 -1.3422 0 -2.0 1e-06 
0.0 -1.3421 0 -2.0 1e-06 
0.0 -1.342 0 -2.0 1e-06 
0.0 -1.3419 0 -2.0 1e-06 
0.0 -1.3418 0 -2.0 1e-06 
0.0 -1.3417 0 -2.0 1e-06 
0.0 -1.3416 0 -2.0 1e-06 
0.0 -1.3415 0 -2.0 1e-06 
0.0 -1.3414 0 -2.0 1e-06 
0.0 -1.3413 0 -2.0 1e-06 
0.0 -1.3412 0 -2.0 1e-06 
0.0 -1.3411 0 -2.0 1e-06 
0.0 -1.341 0 -2.0 1e-06 
0.0 -1.3409 0 -2.0 1e-06 
0.0 -1.3408 0 -2.0 1e-06 
0.0 -1.3407 0 -2.0 1e-06 
0.0 -1.3406 0 -2.0 1e-06 
0.0 -1.3405 0 -2.0 1e-06 
0.0 -1.3404 0 -2.0 1e-06 
0.0 -1.3403 0 -2.0 1e-06 
0.0 -1.3402 0 -2.0 1e-06 
0.0 -1.3401 0 -2.0 1e-06 
0.0 -1.34 0 -2.0 1e-06 
0.0 -1.3399 0 -2.0 1e-06 
0.0 -1.3398 0 -2.0 1e-06 
0.0 -1.3397 0 -2.0 1e-06 
0.0 -1.3396 0 -2.0 1e-06 
0.0 -1.3395 0 -2.0 1e-06 
0.0 -1.3394 0 -2.0 1e-06 
0.0 -1.3393 0 -2.0 1e-06 
0.0 -1.3392 0 -2.0 1e-06 
0.0 -1.3391 0 -2.0 1e-06 
0.0 -1.339 0 -2.0 1e-06 
0.0 -1.3389 0 -2.0 1e-06 
0.0 -1.3388 0 -2.0 1e-06 
0.0 -1.3387 0 -2.0 1e-06 
0.0 -1.3386 0 -2.0 1e-06 
0.0 -1.3385 0 -2.0 1e-06 
0.0 -1.3384 0 -2.0 1e-06 
0.0 -1.3383 0 -2.0 1e-06 
0.0 -1.3382 0 -2.0 1e-06 
0.0 -1.3381 0 -2.0 1e-06 
0.0 -1.338 0 -2.0 1e-06 
0.0 -1.3379 0 -2.0 1e-06 
0.0 -1.3378 0 -2.0 1e-06 
0.0 -1.3377 0 -2.0 1e-06 
0.0 -1.3376 0 -2.0 1e-06 
0.0 -1.3375 0 -2.0 1e-06 
0.0 -1.3374 0 -2.0 1e-06 
0.0 -1.3373 0 -2.0 1e-06 
0.0 -1.3372 0 -2.0 1e-06 
0.0 -1.3371 0 -2.0 1e-06 
0.0 -1.337 0 -2.0 1e-06 
0.0 -1.3369 0 -2.0 1e-06 
0.0 -1.3368 0 -2.0 1e-06 
0.0 -1.3367 0 -2.0 1e-06 
0.0 -1.3366 0 -2.0 1e-06 
0.0 -1.3365 0 -2.0 1e-06 
0.0 -1.3364 0 -2.0 1e-06 
0.0 -1.3363 0 -2.0 1e-06 
0.0 -1.3362 0 -2.0 1e-06 
0.0 -1.3361 0 -2.0 1e-06 
0.0 -1.336 0 -2.0 1e-06 
0.0 -1.3359 0 -2.0 1e-06 
0.0 -1.3358 0 -2.0 1e-06 
0.0 -1.3357 0 -2.0 1e-06 
0.0 -1.3356 0 -2.0 1e-06 
0.0 -1.3355 0 -2.0 1e-06 
0.0 -1.3354 0 -2.0 1e-06 
0.0 -1.3353 0 -2.0 1e-06 
0.0 -1.3352 0 -2.0 1e-06 
0.0 -1.3351 0 -2.0 1e-06 
0.0 -1.335 0 -2.0 1e-06 
0.0 -1.3349 0 -2.0 1e-06 
0.0 -1.3348 0 -2.0 1e-06 
0.0 -1.3347 0 -2.0 1e-06 
0.0 -1.3346 0 -2.0 1e-06 
0.0 -1.3345 0 -2.0 1e-06 
0.0 -1.3344 0 -2.0 1e-06 
0.0 -1.3343 0 -2.0 1e-06 
0.0 -1.3342 0 -2.0 1e-06 
0.0 -1.3341 0 -2.0 1e-06 
0.0 -1.334 0 -2.0 1e-06 
0.0 -1.3339 0 -2.0 1e-06 
0.0 -1.3338 0 -2.0 1e-06 
0.0 -1.3337 0 -2.0 1e-06 
0.0 -1.3336 0 -2.0 1e-06 
0.0 -1.3335 0 -2.0 1e-06 
0.0 -1.3334 0 -2.0 1e-06 
0.0 -1.3333 0 -2.0 1e-06 
0.0 -1.3332 0 -2.0 1e-06 
0.0 -1.3331 0 -2.0 1e-06 
0.0 -1.333 0 -2.0 1e-06 
0.0 -1.3329 0 -2.0 1e-06 
0.0 -1.3328 0 -2.0 1e-06 
0.0 -1.3327 0 -2.0 1e-06 
0.0 -1.3326 0 -2.0 1e-06 
0.0 -1.3325 0 -2.0 1e-06 
0.0 -1.3324 0 -2.0 1e-06 
0.0 -1.3323 0 -2.0 1e-06 
0.0 -1.3322 0 -2.0 1e-06 
0.0 -1.3321 0 -2.0 1e-06 
0.0 -1.332 0 -2.0 1e-06 
0.0 -1.3319 0 -2.0 1e-06 
0.0 -1.3318 0 -2.0 1e-06 
0.0 -1.3317 0 -2.0 1e-06 
0.0 -1.3316 0 -2.0 1e-06 
0.0 -1.3315 0 -2.0 1e-06 
0.0 -1.3314 0 -2.0 1e-06 
0.0 -1.3313 0 -2.0 1e-06 
0.0 -1.3312 0 -2.0 1e-06 
0.0 -1.3311 0 -2.0 1e-06 
0.0 -1.331 0 -2.0 1e-06 
0.0 -1.3309 0 -2.0 1e-06 
0.0 -1.3308 0 -2.0 1e-06 
0.0 -1.3307 0 -2.0 1e-06 
0.0 -1.3306 0 -2.0 1e-06 
0.0 -1.3305 0 -2.0 1e-06 
0.0 -1.3304 0 -2.0 1e-06 
0.0 -1.3303 0 -2.0 1e-06 
0.0 -1.3302 0 -2.0 1e-06 
0.0 -1.3301 0 -2.0 1e-06 
0.0 -1.33 0 -2.0 1e-06 
0.0 -1.3299 0 -2.0 1e-06 
0.0 -1.3298 0 -2.0 1e-06 
0.0 -1.3297 0 -2.0 1e-06 
0.0 -1.3296 0 -2.0 1e-06 
0.0 -1.3295 0 -2.0 1e-06 
0.0 -1.3294 0 -2.0 1e-06 
0.0 -1.3293 0 -2.0 1e-06 
0.0 -1.3292 0 -2.0 1e-06 
0.0 -1.3291 0 -2.0 1e-06 
0.0 -1.329 0 -2.0 1e-06 
0.0 -1.3289 0 -2.0 1e-06 
0.0 -1.3288 0 -2.0 1e-06 
0.0 -1.3287 0 -2.0 1e-06 
0.0 -1.3286 0 -2.0 1e-06 
0.0 -1.3285 0 -2.0 1e-06 
0.0 -1.3284 0 -2.0 1e-06 
0.0 -1.3283 0 -2.0 1e-06 
0.0 -1.3282 0 -2.0 1e-06 
0.0 -1.3281 0 -2.0 1e-06 
0.0 -1.328 0 -2.0 1e-06 
0.0 -1.3279 0 -2.0 1e-06 
0.0 -1.3278 0 -2.0 1e-06 
0.0 -1.3277 0 -2.0 1e-06 
0.0 -1.3276 0 -2.0 1e-06 
0.0 -1.3275 0 -2.0 1e-06 
0.0 -1.3274 0 -2.0 1e-06 
0.0 -1.3273 0 -2.0 1e-06 
0.0 -1.3272 0 -2.0 1e-06 
0.0 -1.3271 0 -2.0 1e-06 
0.0 -1.327 0 -2.0 1e-06 
0.0 -1.3269 0 -2.0 1e-06 
0.0 -1.3268 0 -2.0 1e-06 
0.0 -1.3267 0 -2.0 1e-06 
0.0 -1.3266 0 -2.0 1e-06 
0.0 -1.3265 0 -2.0 1e-06 
0.0 -1.3264 0 -2.0 1e-06 
0.0 -1.3263 0 -2.0 1e-06 
0.0 -1.3262 0 -2.0 1e-06 
0.0 -1.3261 0 -2.0 1e-06 
0.0 -1.326 0 -2.0 1e-06 
0.0 -1.3259 0 -2.0 1e-06 
0.0 -1.3258 0 -2.0 1e-06 
0.0 -1.3257 0 -2.0 1e-06 
0.0 -1.3256 0 -2.0 1e-06 
0.0 -1.3255 0 -2.0 1e-06 
0.0 -1.3254 0 -2.0 1e-06 
0.0 -1.3253 0 -2.0 1e-06 
0.0 -1.3252 0 -2.0 1e-06 
0.0 -1.3251 0 -2.0 1e-06 
0.0 -1.325 0 -2.0 1e-06 
0.0 -1.3249 0 -2.0 1e-06 
0.0 -1.3248 0 -2.0 1e-06 
0.0 -1.3247 0 -2.0 1e-06 
0.0 -1.3246 0 -2.0 1e-06 
0.0 -1.3245 0 -2.0 1e-06 
0.0 -1.3244 0 -2.0 1e-06 
0.0 -1.3243 0 -2.0 1e-06 
0.0 -1.3242 0 -2.0 1e-06 
0.0 -1.3241 0 -2.0 1e-06 
0.0 -1.324 0 -2.0 1e-06 
0.0 -1.3239 0 -2.0 1e-06 
0.0 -1.3238 0 -2.0 1e-06 
0.0 -1.3237 0 -2.0 1e-06 
0.0 -1.3236 0 -2.0 1e-06 
0.0 -1.3235 0 -2.0 1e-06 
0.0 -1.3234 0 -2.0 1e-06 
0.0 -1.3233 0 -2.0 1e-06 
0.0 -1.3232 0 -2.0 1e-06 
0.0 -1.3231 0 -2.0 1e-06 
0.0 -1.323 0 -2.0 1e-06 
0.0 -1.3229 0 -2.0 1e-06 
0.0 -1.3228 0 -2.0 1e-06 
0.0 -1.3227 0 -2.0 1e-06 
0.0 -1.3226 0 -2.0 1e-06 
0.0 -1.3225 0 -2.0 1e-06 
0.0 -1.3224 0 -2.0 1e-06 
0.0 -1.3223 0 -2.0 1e-06 
0.0 -1.3222 0 -2.0 1e-06 
0.0 -1.3221 0 -2.0 1e-06 
0.0 -1.322 0 -2.0 1e-06 
0.0 -1.3219 0 -2.0 1e-06 
0.0 -1.3218 0 -2.0 1e-06 
0.0 -1.3217 0 -2.0 1e-06 
0.0 -1.3216 0 -2.0 1e-06 
0.0 -1.3215 0 -2.0 1e-06 
0.0 -1.3214 0 -2.0 1e-06 
0.0 -1.3213 0 -2.0 1e-06 
0.0 -1.3212 0 -2.0 1e-06 
0.0 -1.3211 0 -2.0 1e-06 
0.0 -1.321 0 -2.0 1e-06 
0.0 -1.3209 0 -2.0 1e-06 
0.0 -1.3208 0 -2.0 1e-06 
0.0 -1.3207 0 -2.0 1e-06 
0.0 -1.3206 0 -2.0 1e-06 
0.0 -1.3205 0 -2.0 1e-06 
0.0 -1.3204 0 -2.0 1e-06 
0.0 -1.3203 0 -2.0 1e-06 
0.0 -1.3202 0 -2.0 1e-06 
0.0 -1.3201 0 -2.0 1e-06 
0.0 -1.32 0 -2.0 1e-06 
0.0 -1.3199 0 -2.0 1e-06 
0.0 -1.3198 0 -2.0 1e-06 
0.0 -1.3197 0 -2.0 1e-06 
0.0 -1.3196 0 -2.0 1e-06 
0.0 -1.3195 0 -2.0 1e-06 
0.0 -1.3194 0 -2.0 1e-06 
0.0 -1.3193 0 -2.0 1e-06 
0.0 -1.3192 0 -2.0 1e-06 
0.0 -1.3191 0 -2.0 1e-06 
0.0 -1.319 0 -2.0 1e-06 
0.0 -1.3189 0 -2.0 1e-06 
0.0 -1.3188 0 -2.0 1e-06 
0.0 -1.3187 0 -2.0 1e-06 
0.0 -1.3186 0 -2.0 1e-06 
0.0 -1.3185 0 -2.0 1e-06 
0.0 -1.3184 0 -2.0 1e-06 
0.0 -1.3183 0 -2.0 1e-06 
0.0 -1.3182 0 -2.0 1e-06 
0.0 -1.3181 0 -2.0 1e-06 
0.0 -1.318 0 -2.0 1e-06 
0.0 -1.3179 0 -2.0 1e-06 
0.0 -1.3178 0 -2.0 1e-06 
0.0 -1.3177 0 -2.0 1e-06 
0.0 -1.3176 0 -2.0 1e-06 
0.0 -1.3175 0 -2.0 1e-06 
0.0 -1.3174 0 -2.0 1e-06 
0.0 -1.3173 0 -2.0 1e-06 
0.0 -1.3172 0 -2.0 1e-06 
0.0 -1.3171 0 -2.0 1e-06 
0.0 -1.317 0 -2.0 1e-06 
0.0 -1.3169 0 -2.0 1e-06 
0.0 -1.3168 0 -2.0 1e-06 
0.0 -1.3167 0 -2.0 1e-06 
0.0 -1.3166 0 -2.0 1e-06 
0.0 -1.3165 0 -2.0 1e-06 
0.0 -1.3164 0 -2.0 1e-06 
0.0 -1.3163 0 -2.0 1e-06 
0.0 -1.3162 0 -2.0 1e-06 
0.0 -1.3161 0 -2.0 1e-06 
0.0 -1.316 0 -2.0 1e-06 
0.0 -1.3159 0 -2.0 1e-06 
0.0 -1.3158 0 -2.0 1e-06 
0.0 -1.3157 0 -2.0 1e-06 
0.0 -1.3156 0 -2.0 1e-06 
0.0 -1.3155 0 -2.0 1e-06 
0.0 -1.3154 0 -2.0 1e-06 
0.0 -1.3153 0 -2.0 1e-06 
0.0 -1.3152 0 -2.0 1e-06 
0.0 -1.3151 0 -2.0 1e-06 
0.0 -1.315 0 -2.0 1e-06 
0.0 -1.3149 0 -2.0 1e-06 
0.0 -1.3148 0 -2.0 1e-06 
0.0 -1.3147 0 -2.0 1e-06 
0.0 -1.3146 0 -2.0 1e-06 
0.0 -1.3145 0 -2.0 1e-06 
0.0 -1.3144 0 -2.0 1e-06 
0.0 -1.3143 0 -2.0 1e-06 
0.0 -1.3142 0 -2.0 1e-06 
0.0 -1.3141 0 -2.0 1e-06 
0.0 -1.314 0 -2.0 1e-06 
0.0 -1.3139 0 -2.0 1e-06 
0.0 -1.3138 0 -2.0 1e-06 
0.0 -1.3137 0 -2.0 1e-06 
0.0 -1.3136 0 -2.0 1e-06 
0.0 -1.3135 0 -2.0 1e-06 
0.0 -1.3134 0 -2.0 1e-06 
0.0 -1.3133 0 -2.0 1e-06 
0.0 -1.3132 0 -2.0 1e-06 
0.0 -1.3131 0 -2.0 1e-06 
0.0 -1.313 0 -2.0 1e-06 
0.0 -1.3129 0 -2.0 1e-06 
0.0 -1.3128 0 -2.0 1e-06 
0.0 -1.3127 0 -2.0 1e-06 
0.0 -1.3126 0 -2.0 1e-06 
0.0 -1.3125 0 -2.0 1e-06 
0.0 -1.3124 0 -2.0 1e-06 
0.0 -1.3123 0 -2.0 1e-06 
0.0 -1.3122 0 -2.0 1e-06 
0.0 -1.3121 0 -2.0 1e-06 
0.0 -1.312 0 -2.0 1e-06 
0.0 -1.3119 0 -2.0 1e-06 
0.0 -1.3118 0 -2.0 1e-06 
0.0 -1.3117 0 -2.0 1e-06 
0.0 -1.3116 0 -2.0 1e-06 
0.0 -1.3115 0 -2.0 1e-06 
0.0 -1.3114 0 -2.0 1e-06 
0.0 -1.3113 0 -2.0 1e-06 
0.0 -1.3112 0 -2.0 1e-06 
0.0 -1.3111 0 -2.0 1e-06 
0.0 -1.311 0 -2.0 1e-06 
0.0 -1.3109 0 -2.0 1e-06 
0.0 -1.3108 0 -2.0 1e-06 
0.0 -1.3107 0 -2.0 1e-06 
0.0 -1.3106 0 -2.0 1e-06 
0.0 -1.3105 0 -2.0 1e-06 
0.0 -1.3104 0 -2.0 1e-06 
0.0 -1.3103 0 -2.0 1e-06 
0.0 -1.3102 0 -2.0 1e-06 
0.0 -1.3101 0 -2.0 1e-06 
0.0 -1.31 0 -2.0 1e-06 
0.0 -1.3099 0 -2.0 1e-06 
0.0 -1.3098 0 -2.0 1e-06 
0.0 -1.3097 0 -2.0 1e-06 
0.0 -1.3096 0 -2.0 1e-06 
0.0 -1.3095 0 -2.0 1e-06 
0.0 -1.3094 0 -2.0 1e-06 
0.0 -1.3093 0 -2.0 1e-06 
0.0 -1.3092 0 -2.0 1e-06 
0.0 -1.3091 0 -2.0 1e-06 
0.0 -1.309 0 -2.0 1e-06 
0.0 -1.3089 0 -2.0 1e-06 
0.0 -1.3088 0 -2.0 1e-06 
0.0 -1.3087 0 -2.0 1e-06 
0.0 -1.3086 0 -2.0 1e-06 
0.0 -1.3085 0 -2.0 1e-06 
0.0 -1.3084 0 -2.0 1e-06 
0.0 -1.3083 0 -2.0 1e-06 
0.0 -1.3082 0 -2.0 1e-06 
0.0 -1.3081 0 -2.0 1e-06 
0.0 -1.308 0 -2.0 1e-06 
0.0 -1.3079 0 -2.0 1e-06 
0.0 -1.3078 0 -2.0 1e-06 
0.0 -1.3077 0 -2.0 1e-06 
0.0 -1.3076 0 -2.0 1e-06 
0.0 -1.3075 0 -2.0 1e-06 
0.0 -1.3074 0 -2.0 1e-06 
0.0 -1.3073 0 -2.0 1e-06 
0.0 -1.3072 0 -2.0 1e-06 
0.0 -1.3071 0 -2.0 1e-06 
0.0 -1.307 0 -2.0 1e-06 
0.0 -1.3069 0 -2.0 1e-06 
0.0 -1.3068 0 -2.0 1e-06 
0.0 -1.3067 0 -2.0 1e-06 
0.0 -1.3066 0 -2.0 1e-06 
0.0 -1.3065 0 -2.0 1e-06 
0.0 -1.3064 0 -2.0 1e-06 
0.0 -1.3063 0 -2.0 1e-06 
0.0 -1.3062 0 -2.0 1e-06 
0.0 -1.3061 0 -2.0 1e-06 
0.0 -1.306 0 -2.0 1e-06 
0.0 -1.3059 0 -2.0 1e-06 
0.0 -1.3058 0 -2.0 1e-06 
0.0 -1.3057 0 -2.0 1e-06 
0.0 -1.3056 0 -2.0 1e-06 
0.0 -1.3055 0 -2.0 1e-06 
0.0 -1.3054 0 -2.0 1e-06 
0.0 -1.3053 0 -2.0 1e-06 
0.0 -1.3052 0 -2.0 1e-06 
0.0 -1.3051 0 -2.0 1e-06 
0.0 -1.305 0 -2.0 1e-06 
0.0 -1.3049 0 -2.0 1e-06 
0.0 -1.3048 0 -2.0 1e-06 
0.0 -1.3047 0 -2.0 1e-06 
0.0 -1.3046 0 -2.0 1e-06 
0.0 -1.3045 0 -2.0 1e-06 
0.0 -1.3044 0 -2.0 1e-06 
0.0 -1.3043 0 -2.0 1e-06 
0.0 -1.3042 0 -2.0 1e-06 
0.0 -1.3041 0 -2.0 1e-06 
0.0 -1.304 0 -2.0 1e-06 
0.0 -1.3039 0 -2.0 1e-06 
0.0 -1.3038 0 -2.0 1e-06 
0.0 -1.3037 0 -2.0 1e-06 
0.0 -1.3036 0 -2.0 1e-06 
0.0 -1.3035 0 -2.0 1e-06 
0.0 -1.3034 0 -2.0 1e-06 
0.0 -1.3033 0 -2.0 1e-06 
0.0 -1.3032 0 -2.0 1e-06 
0.0 -1.3031 0 -2.0 1e-06 
0.0 -1.303 0 -2.0 1e-06 
0.0 -1.3029 0 -2.0 1e-06 
0.0 -1.3028 0 -2.0 1e-06 
0.0 -1.3027 0 -2.0 1e-06 
0.0 -1.3026 0 -2.0 1e-06 
0.0 -1.3025 0 -2.0 1e-06 
0.0 -1.3024 0 -2.0 1e-06 
0.0 -1.3023 0 -2.0 1e-06 
0.0 -1.3022 0 -2.0 1e-06 
0.0 -1.3021 0 -2.0 1e-06 
0.0 -1.302 0 -2.0 1e-06 
0.0 -1.3019 0 -2.0 1e-06 
0.0 -1.3018 0 -2.0 1e-06 
0.0 -1.3017 0 -2.0 1e-06 
0.0 -1.3016 0 -2.0 1e-06 
0.0 -1.3015 0 -2.0 1e-06 
0.0 -1.3014 0 -2.0 1e-06 
0.0 -1.3013 0 -2.0 1e-06 
0.0 -1.3012 0 -2.0 1e-06 
0.0 -1.3011 0 -2.0 1e-06 
0.0 -1.301 0 -2.0 1e-06 
0.0 -1.3009 0 -2.0 1e-06 
0.0 -1.3008 0 -2.0 1e-06 
0.0 -1.3007 0 -2.0 1e-06 
0.0 -1.3006 0 -2.0 1e-06 
0.0 -1.3005 0 -2.0 1e-06 
0.0 -1.3004 0 -2.0 1e-06 
0.0 -1.3003 0 -2.0 1e-06 
0.0 -1.3002 0 -2.0 1e-06 
0.0 -1.3001 0 -2.0 1e-06 
0.0 -1.3 0 -2.0 1e-06 
0.0 -1.2999 0 -2.0 1e-06 
0.0 -1.2998 0 -2.0 1e-06 
0.0 -1.2997 0 -2.0 1e-06 
0.0 -1.2996 0 -2.0 1e-06 
0.0 -1.2995 0 -2.0 1e-06 
0.0 -1.2994 0 -2.0 1e-06 
0.0 -1.2993 0 -2.0 1e-06 
0.0 -1.2992 0 -2.0 1e-06 
0.0 -1.2991 0 -2.0 1e-06 
0.0 -1.299 0 -2.0 1e-06 
0.0 -1.2989 0 -2.0 1e-06 
0.0 -1.2988 0 -2.0 1e-06 
0.0 -1.2987 0 -2.0 1e-06 
0.0 -1.2986 0 -2.0 1e-06 
0.0 -1.2985 0 -2.0 1e-06 
0.0 -1.2984 0 -2.0 1e-06 
0.0 -1.2983 0 -2.0 1e-06 
0.0 -1.2982 0 -2.0 1e-06 
0.0 -1.2981 0 -2.0 1e-06 
0.0 -1.298 0 -2.0 1e-06 
0.0 -1.2979 0 -2.0 1e-06 
0.0 -1.2978 0 -2.0 1e-06 
0.0 -1.2977 0 -2.0 1e-06 
0.0 -1.2976 0 -2.0 1e-06 
0.0 -1.2975 0 -2.0 1e-06 
0.0 -1.2974 0 -2.0 1e-06 
0.0 -1.2973 0 -2.0 1e-06 
0.0 -1.2972 0 -2.0 1e-06 
0.0 -1.2971 0 -2.0 1e-06 
0.0 -1.297 0 -2.0 1e-06 
0.0 -1.2969 0 -2.0 1e-06 
0.0 -1.2968 0 -2.0 1e-06 
0.0 -1.2967 0 -2.0 1e-06 
0.0 -1.2966 0 -2.0 1e-06 
0.0 -1.2965 0 -2.0 1e-06 
0.0 -1.2964 0 -2.0 1e-06 
0.0 -1.2963 0 -2.0 1e-06 
0.0 -1.2962 0 -2.0 1e-06 
0.0 -1.2961 0 -2.0 1e-06 
0.0 -1.296 0 -2.0 1e-06 
0.0 -1.2959 0 -2.0 1e-06 
0.0 -1.2958 0 -2.0 1e-06 
0.0 -1.2957 0 -2.0 1e-06 
0.0 -1.2956 0 -2.0 1e-06 
0.0 -1.2955 0 -2.0 1e-06 
0.0 -1.2954 0 -2.0 1e-06 
0.0 -1.2953 0 -2.0 1e-06 
0.0 -1.2952 0 -2.0 1e-06 
0.0 -1.2951 0 -2.0 1e-06 
0.0 -1.295 0 -2.0 1e-06 
0.0 -1.2949 0 -2.0 1e-06 
0.0 -1.2948 0 -2.0 1e-06 
0.0 -1.2947 0 -2.0 1e-06 
0.0 -1.2946 0 -2.0 1e-06 
0.0 -1.2945 0 -2.0 1e-06 
0.0 -1.2944 0 -2.0 1e-06 
0.0 -1.2943 0 -2.0 1e-06 
0.0 -1.2942 0 -2.0 1e-06 
0.0 -1.2941 0 -2.0 1e-06 
0.0 -1.294 0 -2.0 1e-06 
0.0 -1.2939 0 -2.0 1e-06 
0.0 -1.2938 0 -2.0 1e-06 
0.0 -1.2937 0 -2.0 1e-06 
0.0 -1.2936 0 -2.0 1e-06 
0.0 -1.2935 0 -2.0 1e-06 
0.0 -1.2934 0 -2.0 1e-06 
0.0 -1.2933 0 -2.0 1e-06 
0.0 -1.2932 0 -2.0 1e-06 
0.0 -1.2931 0 -2.0 1e-06 
0.0 -1.293 0 -2.0 1e-06 
0.0 -1.2929 0 -2.0 1e-06 
0.0 -1.2928 0 -2.0 1e-06 
0.0 -1.2927 0 -2.0 1e-06 
0.0 -1.2926 0 -2.0 1e-06 
0.0 -1.2925 0 -2.0 1e-06 
0.0 -1.2924 0 -2.0 1e-06 
0.0 -1.2923 0 -2.0 1e-06 
0.0 -1.2922 0 -2.0 1e-06 
0.0 -1.2921 0 -2.0 1e-06 
0.0 -1.292 0 -2.0 1e-06 
0.0 -1.2919 0 -2.0 1e-06 
0.0 -1.2918 0 -2.0 1e-06 
0.0 -1.2917 0 -2.0 1e-06 
0.0 -1.2916 0 -2.0 1e-06 
0.0 -1.2915 0 -2.0 1e-06 
0.0 -1.2914 0 -2.0 1e-06 
0.0 -1.2913 0 -2.0 1e-06 
0.0 -1.2912 0 -2.0 1e-06 
0.0 -1.2911 0 -2.0 1e-06 
0.0 -1.291 0 -2.0 1e-06 
0.0 -1.2909 0 -2.0 1e-06 
0.0 -1.2908 0 -2.0 1e-06 
0.0 -1.2907 0 -2.0 1e-06 
0.0 -1.2906 0 -2.0 1e-06 
0.0 -1.2905 0 -2.0 1e-06 
0.0 -1.2904 0 -2.0 1e-06 
0.0 -1.2903 0 -2.0 1e-06 
0.0 -1.2902 0 -2.0 1e-06 
0.0 -1.2901 0 -2.0 1e-06 
0.0 -1.29 0 -2.0 1e-06 
0.0 -1.2899 0 -2.0 1e-06 
0.0 -1.2898 0 -2.0 1e-06 
0.0 -1.2897 0 -2.0 1e-06 
0.0 -1.2896 0 -2.0 1e-06 
0.0 -1.2895 0 -2.0 1e-06 
0.0 -1.2894 0 -2.0 1e-06 
0.0 -1.2893 0 -2.0 1e-06 
0.0 -1.2892 0 -2.0 1e-06 
0.0 -1.2891 0 -2.0 1e-06 
0.0 -1.289 0 -2.0 1e-06 
0.0 -1.2889 0 -2.0 1e-06 
0.0 -1.2888 0 -2.0 1e-06 
0.0 -1.2887 0 -2.0 1e-06 
0.0 -1.2886 0 -2.0 1e-06 
0.0 -1.2885 0 -2.0 1e-06 
0.0 -1.2884 0 -2.0 1e-06 
0.0 -1.2883 0 -2.0 1e-06 
0.0 -1.2882 0 -2.0 1e-06 
0.0 -1.2881 0 -2.0 1e-06 
0.0 -1.288 0 -2.0 1e-06 
0.0 -1.2879 0 -2.0 1e-06 
0.0 -1.2878 0 -2.0 1e-06 
0.0 -1.2877 0 -2.0 1e-06 
0.0 -1.2876 0 -2.0 1e-06 
0.0 -1.2875 0 -2.0 1e-06 
0.0 -1.2874 0 -2.0 1e-06 
0.0 -1.2873 0 -2.0 1e-06 
0.0 -1.2872 0 -2.0 1e-06 
0.0 -1.2871 0 -2.0 1e-06 
0.0 -1.287 0 -2.0 1e-06 
0.0 -1.2869 0 -2.0 1e-06 
0.0 -1.2868 0 -2.0 1e-06 
0.0 -1.2867 0 -2.0 1e-06 
0.0 -1.2866 0 -2.0 1e-06 
0.0 -1.2865 0 -2.0 1e-06 
0.0 -1.2864 0 -2.0 1e-06 
0.0 -1.2863 0 -2.0 1e-06 
0.0 -1.2862 0 -2.0 1e-06 
0.0 -1.2861 0 -2.0 1e-06 
0.0 -1.286 0 -2.0 1e-06 
0.0 -1.2859 0 -2.0 1e-06 
0.0 -1.2858 0 -2.0 1e-06 
0.0 -1.2857 0 -2.0 1e-06 
0.0 -1.2856 0 -2.0 1e-06 
0.0 -1.2855 0 -2.0 1e-06 
0.0 -1.2854 0 -2.0 1e-06 
0.0 -1.2853 0 -2.0 1e-06 
0.0 -1.2852 0 -2.0 1e-06 
0.0 -1.2851 0 -2.0 1e-06 
0.0 -1.285 0 -2.0 1e-06 
0.0 -1.2849 0 -2.0 1e-06 
0.0 -1.2848 0 -2.0 1e-06 
0.0 -1.2847 0 -2.0 1e-06 
0.0 -1.2846 0 -2.0 1e-06 
0.0 -1.2845 0 -2.0 1e-06 
0.0 -1.2844 0 -2.0 1e-06 
0.0 -1.2843 0 -2.0 1e-06 
0.0 -1.2842 0 -2.0 1e-06 
0.0 -1.2841 0 -2.0 1e-06 
0.0 -1.284 0 -2.0 1e-06 
0.0 -1.2839 0 -2.0 1e-06 
0.0 -1.2838 0 -2.0 1e-06 
0.0 -1.2837 0 -2.0 1e-06 
0.0 -1.2836 0 -2.0 1e-06 
0.0 -1.2835 0 -2.0 1e-06 
0.0 -1.2834 0 -2.0 1e-06 
0.0 -1.2833 0 -2.0 1e-06 
0.0 -1.2832 0 -2.0 1e-06 
0.0 -1.2831 0 -2.0 1e-06 
0.0 -1.283 0 -2.0 1e-06 
0.0 -1.2829 0 -2.0 1e-06 
0.0 -1.2828 0 -2.0 1e-06 
0.0 -1.2827 0 -2.0 1e-06 
0.0 -1.2826 0 -2.0 1e-06 
0.0 -1.2825 0 -2.0 1e-06 
0.0 -1.2824 0 -2.0 1e-06 
0.0 -1.2823 0 -2.0 1e-06 
0.0 -1.2822 0 -2.0 1e-06 
0.0 -1.2821 0 -2.0 1e-06 
0.0 -1.282 0 -2.0 1e-06 
0.0 -1.2819 0 -2.0 1e-06 
0.0 -1.2818 0 -2.0 1e-06 
0.0 -1.2817 0 -2.0 1e-06 
0.0 -1.2816 0 -2.0 1e-06 
0.0 -1.2815 0 -2.0 1e-06 
0.0 -1.2814 0 -2.0 1e-06 
0.0 -1.2813 0 -2.0 1e-06 
0.0 -1.2812 0 -2.0 1e-06 
0.0 -1.2811 0 -2.0 1e-06 
0.0 -1.281 0 -2.0 1e-06 
0.0 -1.2809 0 -2.0 1e-06 
0.0 -1.2808 0 -2.0 1e-06 
0.0 -1.2807 0 -2.0 1e-06 
0.0 -1.2806 0 -2.0 1e-06 
0.0 -1.2805 0 -2.0 1e-06 
0.0 -1.2804 0 -2.0 1e-06 
0.0 -1.2803 0 -2.0 1e-06 
0.0 -1.2802 0 -2.0 1e-06 
0.0 -1.2801 0 -2.0 1e-06 
0.0 -1.28 0 -2.0 1e-06 
0.0 -1.2799 0 -2.0 1e-06 
0.0 -1.2798 0 -2.0 1e-06 
0.0 -1.2797 0 -2.0 1e-06 
0.0 -1.2796 0 -2.0 1e-06 
0.0 -1.2795 0 -2.0 1e-06 
0.0 -1.2794 0 -2.0 1e-06 
0.0 -1.2793 0 -2.0 1e-06 
0.0 -1.2792 0 -2.0 1e-06 
0.0 -1.2791 0 -2.0 1e-06 
0.0 -1.279 0 -2.0 1e-06 
0.0 -1.2789 0 -2.0 1e-06 
0.0 -1.2788 0 -2.0 1e-06 
0.0 -1.2787 0 -2.0 1e-06 
0.0 -1.2786 0 -2.0 1e-06 
0.0 -1.2785 0 -2.0 1e-06 
0.0 -1.2784 0 -2.0 1e-06 
0.0 -1.2783 0 -2.0 1e-06 
0.0 -1.2782 0 -2.0 1e-06 
0.0 -1.2781 0 -2.0 1e-06 
0.0 -1.278 0 -2.0 1e-06 
0.0 -1.2779 0 -2.0 1e-06 
0.0 -1.2778 0 -2.0 1e-06 
0.0 -1.2777 0 -2.0 1e-06 
0.0 -1.2776 0 -2.0 1e-06 
0.0 -1.2775 0 -2.0 1e-06 
0.0 -1.2774 0 -2.0 1e-06 
0.0 -1.2773 0 -2.0 1e-06 
0.0 -1.2772 0 -2.0 1e-06 
0.0 -1.2771 0 -2.0 1e-06 
0.0 -1.277 0 -2.0 1e-06 
0.0 -1.2769 0 -2.0 1e-06 
0.0 -1.2768 0 -2.0 1e-06 
0.0 -1.2767 0 -2.0 1e-06 
0.0 -1.2766 0 -2.0 1e-06 
0.0 -1.2765 0 -2.0 1e-06 
0.0 -1.2764 0 -2.0 1e-06 
0.0 -1.2763 0 -2.0 1e-06 
0.0 -1.2762 0 -2.0 1e-06 
0.0 -1.2761 0 -2.0 1e-06 
0.0 -1.276 0 -2.0 1e-06 
0.0 -1.2759 0 -2.0 1e-06 
0.0 -1.2758 0 -2.0 1e-06 
0.0 -1.2757 0 -2.0 1e-06 
0.0 -1.2756 0 -2.0 1e-06 
0.0 -1.2755 0 -2.0 1e-06 
0.0 -1.2754 0 -2.0 1e-06 
0.0 -1.2753 0 -2.0 1e-06 
0.0 -1.2752 0 -2.0 1e-06 
0.0 -1.2751 0 -2.0 1e-06 
0.0 -1.275 0 -2.0 1e-06 
0.0 -1.2749 0 -2.0 1e-06 
0.0 -1.2748 0 -2.0 1e-06 
0.0 -1.2747 0 -2.0 1e-06 
0.0 -1.2746 0 -2.0 1e-06 
0.0 -1.2745 0 -2.0 1e-06 
0.0 -1.2744 0 -2.0 1e-06 
0.0 -1.2743 0 -2.0 1e-06 
0.0 -1.2742 0 -2.0 1e-06 
0.0 -1.2741 0 -2.0 1e-06 
0.0 -1.274 0 -2.0 1e-06 
0.0 -1.2739 0 -2.0 1e-06 
0.0 -1.2738 0 -2.0 1e-06 
0.0 -1.2737 0 -2.0 1e-06 
0.0 -1.2736 0 -2.0 1e-06 
0.0 -1.2735 0 -2.0 1e-06 
0.0 -1.2734 0 -2.0 1e-06 
0.0 -1.2733 0 -2.0 1e-06 
0.0 -1.2732 0 -2.0 1e-06 
0.0 -1.2731 0 -2.0 1e-06 
0.0 -1.273 0 -2.0 1e-06 
0.0 -1.2729 0 -2.0 1e-06 
0.0 -1.2728 0 -2.0 1e-06 
0.0 -1.2727 0 -2.0 1e-06 
0.0 -1.2726 0 -2.0 1e-06 
0.0 -1.2725 0 -2.0 1e-06 
0.0 -1.2724 0 -2.0 1e-06 
0.0 -1.2723 0 -2.0 1e-06 
0.0 -1.2722 0 -2.0 1e-06 
0.0 -1.2721 0 -2.0 1e-06 
0.0 -1.272 0 -2.0 1e-06 
0.0 -1.2719 0 -2.0 1e-06 
0.0 -1.2718 0 -2.0 1e-06 
0.0 -1.2717 0 -2.0 1e-06 
0.0 -1.2716 0 -2.0 1e-06 
0.0 -1.2715 0 -2.0 1e-06 
0.0 -1.2714 0 -2.0 1e-06 
0.0 -1.2713 0 -2.0 1e-06 
0.0 -1.2712 0 -2.0 1e-06 
0.0 -1.2711 0 -2.0 1e-06 
0.0 -1.271 0 -2.0 1e-06 
0.0 -1.2709 0 -2.0 1e-06 
0.0 -1.2708 0 -2.0 1e-06 
0.0 -1.2707 0 -2.0 1e-06 
0.0 -1.2706 0 -2.0 1e-06 
0.0 -1.2705 0 -2.0 1e-06 
0.0 -1.2704 0 -2.0 1e-06 
0.0 -1.2703 0 -2.0 1e-06 
0.0 -1.2702 0 -2.0 1e-06 
0.0 -1.2701 0 -2.0 1e-06 
0.0 -1.27 0 -2.0 1e-06 
0.0 -1.2699 0 -2.0 1e-06 
0.0 -1.2698 0 -2.0 1e-06 
0.0 -1.2697 0 -2.0 1e-06 
0.0 -1.2696 0 -2.0 1e-06 
0.0 -1.2695 0 -2.0 1e-06 
0.0 -1.2694 0 -2.0 1e-06 
0.0 -1.2693 0 -2.0 1e-06 
0.0 -1.2692 0 -2.0 1e-06 
0.0 -1.2691 0 -2.0 1e-06 
0.0 -1.269 0 -2.0 1e-06 
0.0 -1.2689 0 -2.0 1e-06 
0.0 -1.2688 0 -2.0 1e-06 
0.0 -1.2687 0 -2.0 1e-06 
0.0 -1.2686 0 -2.0 1e-06 
0.0 -1.2685 0 -2.0 1e-06 
0.0 -1.2684 0 -2.0 1e-06 
0.0 -1.2683 0 -2.0 1e-06 
0.0 -1.2682 0 -2.0 1e-06 
0.0 -1.2681 0 -2.0 1e-06 
0.0 -1.268 0 -2.0 1e-06 
0.0 -1.2679 0 -2.0 1e-06 
0.0 -1.2678 0 -2.0 1e-06 
0.0 -1.2677 0 -2.0 1e-06 
0.0 -1.2676 0 -2.0 1e-06 
0.0 -1.2675 0 -2.0 1e-06 
0.0 -1.2674 0 -2.0 1e-06 
0.0 -1.2673 0 -2.0 1e-06 
0.0 -1.2672 0 -2.0 1e-06 
0.0 -1.2671 0 -2.0 1e-06 
0.0 -1.267 0 -2.0 1e-06 
0.0 -1.2669 0 -2.0 1e-06 
0.0 -1.2668 0 -2.0 1e-06 
0.0 -1.2667 0 -2.0 1e-06 
0.0 -1.2666 0 -2.0 1e-06 
0.0 -1.2665 0 -2.0 1e-06 
0.0 -1.2664 0 -2.0 1e-06 
0.0 -1.2663 0 -2.0 1e-06 
0.0 -1.2662 0 -2.0 1e-06 
0.0 -1.2661 0 -2.0 1e-06 
0.0 -1.266 0 -2.0 1e-06 
0.0 -1.2659 0 -2.0 1e-06 
0.0 -1.2658 0 -2.0 1e-06 
0.0 -1.2657 0 -2.0 1e-06 
0.0 -1.2656 0 -2.0 1e-06 
0.0 -1.2655 0 -2.0 1e-06 
0.0 -1.2654 0 -2.0 1e-06 
0.0 -1.2653 0 -2.0 1e-06 
0.0 -1.2652 0 -2.0 1e-06 
0.0 -1.2651 0 -2.0 1e-06 
0.0 -1.265 0 -2.0 1e-06 
0.0 -1.2649 0 -2.0 1e-06 
0.0 -1.2648 0 -2.0 1e-06 
0.0 -1.2647 0 -2.0 1e-06 
0.0 -1.2646 0 -2.0 1e-06 
0.0 -1.2645 0 -2.0 1e-06 
0.0 -1.2644 0 -2.0 1e-06 
0.0 -1.2643 0 -2.0 1e-06 
0.0 -1.2642 0 -2.0 1e-06 
0.0 -1.2641 0 -2.0 1e-06 
0.0 -1.264 0 -2.0 1e-06 
0.0 -1.2639 0 -2.0 1e-06 
0.0 -1.2638 0 -2.0 1e-06 
0.0 -1.2637 0 -2.0 1e-06 
0.0 -1.2636 0 -2.0 1e-06 
0.0 -1.2635 0 -2.0 1e-06 
0.0 -1.2634 0 -2.0 1e-06 
0.0 -1.2633 0 -2.0 1e-06 
0.0 -1.2632 0 -2.0 1e-06 
0.0 -1.2631 0 -2.0 1e-06 
0.0 -1.263 0 -2.0 1e-06 
0.0 -1.2629 0 -2.0 1e-06 
0.0 -1.2628 0 -2.0 1e-06 
0.0 -1.2627 0 -2.0 1e-06 
0.0 -1.2626 0 -2.0 1e-06 
0.0 -1.2625 0 -2.0 1e-06 
0.0 -1.2624 0 -2.0 1e-06 
0.0 -1.2623 0 -2.0 1e-06 
0.0 -1.2622 0 -2.0 1e-06 
0.0 -1.2621 0 -2.0 1e-06 
0.0 -1.262 0 -2.0 1e-06 
0.0 -1.2619 0 -2.0 1e-06 
0.0 -1.2618 0 -2.0 1e-06 
0.0 -1.2617 0 -2.0 1e-06 
0.0 -1.2616 0 -2.0 1e-06 
0.0 -1.2615 0 -2.0 1e-06 
0.0 -1.2614 0 -2.0 1e-06 
0.0 -1.2613 0 -2.0 1e-06 
0.0 -1.2612 0 -2.0 1e-06 
0.0 -1.2611 0 -2.0 1e-06 
0.0 -1.261 0 -2.0 1e-06 
0.0 -1.2609 0 -2.0 1e-06 
0.0 -1.2608 0 -2.0 1e-06 
0.0 -1.2607 0 -2.0 1e-06 
0.0 -1.2606 0 -2.0 1e-06 
0.0 -1.2605 0 -2.0 1e-06 
0.0 -1.2604 0 -2.0 1e-06 
0.0 -1.2603 0 -2.0 1e-06 
0.0 -1.2602 0 -2.0 1e-06 
0.0 -1.2601 0 -2.0 1e-06 
0.0 -1.26 0 -2.0 1e-06 
0.0 -1.2599 0 -2.0 1e-06 
0.0 -1.2598 0 -2.0 1e-06 
0.0 -1.2597 0 -2.0 1e-06 
0.0 -1.2596 0 -2.0 1e-06 
0.0 -1.2595 0 -2.0 1e-06 
0.0 -1.2594 0 -2.0 1e-06 
0.0 -1.2593 0 -2.0 1e-06 
0.0 -1.2592 0 -2.0 1e-06 
0.0 -1.2591 0 -2.0 1e-06 
0.0 -1.259 0 -2.0 1e-06 
0.0 -1.2589 0 -2.0 1e-06 
0.0 -1.2588 0 -2.0 1e-06 
0.0 -1.2587 0 -2.0 1e-06 
0.0 -1.2586 0 -2.0 1e-06 
0.0 -1.2585 0 -2.0 1e-06 
0.0 -1.2584 0 -2.0 1e-06 
0.0 -1.2583 0 -2.0 1e-06 
0.0 -1.2582 0 -2.0 1e-06 
0.0 -1.2581 0 -2.0 1e-06 
0.0 -1.258 0 -2.0 1e-06 
0.0 -1.2579 0 -2.0 1e-06 
0.0 -1.2578 0 -2.0 1e-06 
0.0 -1.2577 0 -2.0 1e-06 
0.0 -1.2576 0 -2.0 1e-06 
0.0 -1.2575 0 -2.0 1e-06 
0.0 -1.2574 0 -2.0 1e-06 
0.0 -1.2573 0 -2.0 1e-06 
0.0 -1.2572 0 -2.0 1e-06 
0.0 -1.2571 0 -2.0 1e-06 
0.0 -1.257 0 -2.0 1e-06 
0.0 -1.2569 0 -2.0 1e-06 
0.0 -1.2568 0 -2.0 1e-06 
0.0 -1.2567 0 -2.0 1e-06 
0.0 -1.2566 0 -2.0 1e-06 
0.0 -1.2565 0 -2.0 1e-06 
0.0 -1.2564 0 -2.0 1e-06 
0.0 -1.2563 0 -2.0 1e-06 
0.0 -1.2562 0 -2.0 1e-06 
0.0 -1.2561 0 -2.0 1e-06 
0.0 -1.256 0 -2.0 1e-06 
0.0 -1.2559 0 -2.0 1e-06 
0.0 -1.2558 0 -2.0 1e-06 
0.0 -1.2557 0 -2.0 1e-06 
0.0 -1.2556 0 -2.0 1e-06 
0.0 -1.2555 0 -2.0 1e-06 
0.0 -1.2554 0 -2.0 1e-06 
0.0 -1.2553 0 -2.0 1e-06 
0.0 -1.2552 0 -2.0 1e-06 
0.0 -1.2551 0 -2.0 1e-06 
0.0 -1.255 0 -2.0 1e-06 
0.0 -1.2549 0 -2.0 1e-06 
0.0 -1.2548 0 -2.0 1e-06 
0.0 -1.2547 0 -2.0 1e-06 
0.0 -1.2546 0 -2.0 1e-06 
0.0 -1.2545 0 -2.0 1e-06 
0.0 -1.2544 0 -2.0 1e-06 
0.0 -1.2543 0 -2.0 1e-06 
0.0 -1.2542 0 -2.0 1e-06 
0.0 -1.2541 0 -2.0 1e-06 
0.0 -1.254 0 -2.0 1e-06 
0.0 -1.2539 0 -2.0 1e-06 
0.0 -1.2538 0 -2.0 1e-06 
0.0 -1.2537 0 -2.0 1e-06 
0.0 -1.2536 0 -2.0 1e-06 
0.0 -1.2535 0 -2.0 1e-06 
0.0 -1.2534 0 -2.0 1e-06 
0.0 -1.2533 0 -2.0 1e-06 
0.0 -1.2532 0 -2.0 1e-06 
0.0 -1.2531 0 -2.0 1e-06 
0.0 -1.253 0 -2.0 1e-06 
0.0 -1.2529 0 -2.0 1e-06 
0.0 -1.2528 0 -2.0 1e-06 
0.0 -1.2527 0 -2.0 1e-06 
0.0 -1.2526 0 -2.0 1e-06 
0.0 -1.2525 0 -2.0 1e-06 
0.0 -1.2524 0 -2.0 1e-06 
0.0 -1.2523 0 -2.0 1e-06 
0.0 -1.2522 0 -2.0 1e-06 
0.0 -1.2521 0 -2.0 1e-06 
0.0 -1.252 0 -2.0 1e-06 
0.0 -1.2519 0 -2.0 1e-06 
0.0 -1.2518 0 -2.0 1e-06 
0.0 -1.2517 0 -2.0 1e-06 
0.0 -1.2516 0 -2.0 1e-06 
0.0 -1.2515 0 -2.0 1e-06 
0.0 -1.2514 0 -2.0 1e-06 
0.0 -1.2513 0 -2.0 1e-06 
0.0 -1.2512 0 -2.0 1e-06 
0.0 -1.2511 0 -2.0 1e-06 
0.0 -1.251 0 -2.0 1e-06 
0.0 -1.2509 0 -2.0 1e-06 
0.0 -1.2508 0 -2.0 1e-06 
0.0 -1.2507 0 -2.0 1e-06 
0.0 -1.2506 0 -2.0 1e-06 
0.0 -1.2505 0 -2.0 1e-06 
0.0 -1.2504 0 -2.0 1e-06 
0.0 -1.2503 0 -2.0 1e-06 
0.0 -1.2502 0 -2.0 1e-06 
0.0 -1.2501 0 -2.0 1e-06 
0.0 -1.25 0 -2.0 1e-06 
0.0 -1.2499 0 -2.0 1e-06 
0.0 -1.2498 0 -2.0 1e-06 
0.0 -1.2497 0 -2.0 1e-06 
0.0 -1.2496 0 -2.0 1e-06 
0.0 -1.2495 0 -2.0 1e-06 
0.0 -1.2494 0 -2.0 1e-06 
0.0 -1.2493 0 -2.0 1e-06 
0.0 -1.2492 0 -2.0 1e-06 
0.0 -1.2491 0 -2.0 1e-06 
0.0 -1.249 0 -2.0 1e-06 
0.0 -1.2489 0 -2.0 1e-06 
0.0 -1.2488 0 -2.0 1e-06 
0.0 -1.2487 0 -2.0 1e-06 
0.0 -1.2486 0 -2.0 1e-06 
0.0 -1.2485 0 -2.0 1e-06 
0.0 -1.2484 0 -2.0 1e-06 
0.0 -1.2483 0 -2.0 1e-06 
0.0 -1.2482 0 -2.0 1e-06 
0.0 -1.2481 0 -2.0 1e-06 
0.0 -1.248 0 -2.0 1e-06 
0.0 -1.2479 0 -2.0 1e-06 
0.0 -1.2478 0 -2.0 1e-06 
0.0 -1.2477 0 -2.0 1e-06 
0.0 -1.2476 0 -2.0 1e-06 
0.0 -1.2475 0 -2.0 1e-06 
0.0 -1.2474 0 -2.0 1e-06 
0.0 -1.2473 0 -2.0 1e-06 
0.0 -1.2472 0 -2.0 1e-06 
0.0 -1.2471 0 -2.0 1e-06 
0.0 -1.247 0 -2.0 1e-06 
0.0 -1.2469 0 -2.0 1e-06 
0.0 -1.2468 0 -2.0 1e-06 
0.0 -1.2467 0 -2.0 1e-06 
0.0 -1.2466 0 -2.0 1e-06 
0.0 -1.2465 0 -2.0 1e-06 
0.0 -1.2464 0 -2.0 1e-06 
0.0 -1.2463 0 -2.0 1e-06 
0.0 -1.2462 0 -2.0 1e-06 
0.0 -1.2461 0 -2.0 1e-06 
0.0 -1.246 0 -2.0 1e-06 
0.0 -1.2459 0 -2.0 1e-06 
0.0 -1.2458 0 -2.0 1e-06 
0.0 -1.2457 0 -2.0 1e-06 
0.0 -1.2456 0 -2.0 1e-06 
0.0 -1.2455 0 -2.0 1e-06 
0.0 -1.2454 0 -2.0 1e-06 
0.0 -1.2453 0 -2.0 1e-06 
0.0 -1.2452 0 -2.0 1e-06 
0.0 -1.2451 0 -2.0 1e-06 
0.0 -1.245 0 -2.0 1e-06 
0.0 -1.2449 0 -2.0 1e-06 
0.0 -1.2448 0 -2.0 1e-06 
0.0 -1.2447 0 -2.0 1e-06 
0.0 -1.2446 0 -2.0 1e-06 
0.0 -1.2445 0 -2.0 1e-06 
0.0 -1.2444 0 -2.0 1e-06 
0.0 -1.2443 0 -2.0 1e-06 
0.0 -1.2442 0 -2.0 1e-06 
0.0 -1.2441 0 -2.0 1e-06 
0.0 -1.244 0 -2.0 1e-06 
0.0 -1.2439 0 -2.0 1e-06 
0.0 -1.2438 0 -2.0 1e-06 
0.0 -1.2437 0 -2.0 1e-06 
0.0 -1.2436 0 -2.0 1e-06 
0.0 -1.2435 0 -2.0 1e-06 
0.0 -1.2434 0 -2.0 1e-06 
0.0 -1.2433 0 -2.0 1e-06 
0.0 -1.2432 0 -2.0 1e-06 
0.0 -1.2431 0 -2.0 1e-06 
0.0 -1.243 0 -2.0 1e-06 
0.0 -1.2429 0 -2.0 1e-06 
0.0 -1.2428 0 -2.0 1e-06 
0.0 -1.2427 0 -2.0 1e-06 
0.0 -1.2426 0 -2.0 1e-06 
0.0 -1.2425 0 -2.0 1e-06 
0.0 -1.2424 0 -2.0 1e-06 
0.0 -1.2423 0 -2.0 1e-06 
0.0 -1.2422 0 -2.0 1e-06 
0.0 -1.2421 0 -2.0 1e-06 
0.0 -1.242 0 -2.0 1e-06 
0.0 -1.2419 0 -2.0 1e-06 
0.0 -1.2418 0 -2.0 1e-06 
0.0 -1.2417 0 -2.0 1e-06 
0.0 -1.2416 0 -2.0 1e-06 
0.0 -1.2415 0 -2.0 1e-06 
0.0 -1.2414 0 -2.0 1e-06 
0.0 -1.2413 0 -2.0 1e-06 
0.0 -1.2412 0 -2.0 1e-06 
0.0 -1.2411 0 -2.0 1e-06 
0.0 -1.241 0 -2.0 1e-06 
0.0 -1.2409 0 -2.0 1e-06 
0.0 -1.2408 0 -2.0 1e-06 
0.0 -1.2407 0 -2.0 1e-06 
0.0 -1.2406 0 -2.0 1e-06 
0.0 -1.2405 0 -2.0 1e-06 
0.0 -1.2404 0 -2.0 1e-06 
0.0 -1.2403 0 -2.0 1e-06 
0.0 -1.2402 0 -2.0 1e-06 
0.0 -1.2401 0 -2.0 1e-06 
0.0 -1.24 0 -2.0 1e-06 
0.0 -1.2399 0 -2.0 1e-06 
0.0 -1.2398 0 -2.0 1e-06 
0.0 -1.2397 0 -2.0 1e-06 
0.0 -1.2396 0 -2.0 1e-06 
0.0 -1.2395 0 -2.0 1e-06 
0.0 -1.2394 0 -2.0 1e-06 
0.0 -1.2393 0 -2.0 1e-06 
0.0 -1.2392 0 -2.0 1e-06 
0.0 -1.2391 0 -2.0 1e-06 
0.0 -1.239 0 -2.0 1e-06 
0.0 -1.2389 0 -2.0 1e-06 
0.0 -1.2388 0 -2.0 1e-06 
0.0 -1.2387 0 -2.0 1e-06 
0.0 -1.2386 0 -2.0 1e-06 
0.0 -1.2385 0 -2.0 1e-06 
0.0 -1.2384 0 -2.0 1e-06 
0.0 -1.2383 0 -2.0 1e-06 
0.0 -1.2382 0 -2.0 1e-06 
0.0 -1.2381 0 -2.0 1e-06 
0.0 -1.238 0 -2.0 1e-06 
0.0 -1.2379 0 -2.0 1e-06 
0.0 -1.2378 0 -2.0 1e-06 
0.0 -1.2377 0 -2.0 1e-06 
0.0 -1.2376 0 -2.0 1e-06 
0.0 -1.2375 0 -2.0 1e-06 
0.0 -1.2374 0 -2.0 1e-06 
0.0 -1.2373 0 -2.0 1e-06 
0.0 -1.2372 0 -2.0 1e-06 
0.0 -1.2371 0 -2.0 1e-06 
0.0 -1.237 0 -2.0 1e-06 
0.0 -1.2369 0 -2.0 1e-06 
0.0 -1.2368 0 -2.0 1e-06 
0.0 -1.2367 0 -2.0 1e-06 
0.0 -1.2366 0 -2.0 1e-06 
0.0 -1.2365 0 -2.0 1e-06 
0.0 -1.2364 0 -2.0 1e-06 
0.0 -1.2363 0 -2.0 1e-06 
0.0 -1.2362 0 -2.0 1e-06 
0.0 -1.2361 0 -2.0 1e-06 
0.0 -1.236 0 -2.0 1e-06 
0.0 -1.2359 0 -2.0 1e-06 
0.0 -1.2358 0 -2.0 1e-06 
0.0 -1.2357 0 -2.0 1e-06 
0.0 -1.2356 0 -2.0 1e-06 
0.0 -1.2355 0 -2.0 1e-06 
0.0 -1.2354 0 -2.0 1e-06 
0.0 -1.2353 0 -2.0 1e-06 
0.0 -1.2352 0 -2.0 1e-06 
0.0 -1.2351 0 -2.0 1e-06 
0.0 -1.235 0 -2.0 1e-06 
0.0 -1.2349 0 -2.0 1e-06 
0.0 -1.2348 0 -2.0 1e-06 
0.0 -1.2347 0 -2.0 1e-06 
0.0 -1.2346 0 -2.0 1e-06 
0.0 -1.2345 0 -2.0 1e-06 
0.0 -1.2344 0 -2.0 1e-06 
0.0 -1.2343 0 -2.0 1e-06 
0.0 -1.2342 0 -2.0 1e-06 
0.0 -1.2341 0 -2.0 1e-06 
0.0 -1.234 0 -2.0 1e-06 
0.0 -1.2339 0 -2.0 1e-06 
0.0 -1.2338 0 -2.0 1e-06 
0.0 -1.2337 0 -2.0 1e-06 
0.0 -1.2336 0 -2.0 1e-06 
0.0 -1.2335 0 -2.0 1e-06 
0.0 -1.2334 0 -2.0 1e-06 
0.0 -1.2333 0 -2.0 1e-06 
0.0 -1.2332 0 -2.0 1e-06 
0.0 -1.2331 0 -2.0 1e-06 
0.0 -1.233 0 -2.0 1e-06 
0.0 -1.2329 0 -2.0 1e-06 
0.0 -1.2328 0 -2.0 1e-06 
0.0 -1.2327 0 -2.0 1e-06 
0.0 -1.2326 0 -2.0 1e-06 
0.0 -1.2325 0 -2.0 1e-06 
0.0 -1.2324 0 -2.0 1e-06 
0.0 -1.2323 0 -2.0 1e-06 
0.0 -1.2322 0 -2.0 1e-06 
0.0 -1.2321 0 -2.0 1e-06 
0.0 -1.232 0 -2.0 1e-06 
0.0 -1.2319 0 -2.0 1e-06 
0.0 -1.2318 0 -2.0 1e-06 
0.0 -1.2317 0 -2.0 1e-06 
0.0 -1.2316 0 -2.0 1e-06 
0.0 -1.2315 0 -2.0 1e-06 
0.0 -1.2314 0 -2.0 1e-06 
0.0 -1.2313 0 -2.0 1e-06 
0.0 -1.2312 0 -2.0 1e-06 
0.0 -1.2311 0 -2.0 1e-06 
0.0 -1.231 0 -2.0 1e-06 
0.0 -1.2309 0 -2.0 1e-06 
0.0 -1.2308 0 -2.0 1e-06 
0.0 -1.2307 0 -2.0 1e-06 
0.0 -1.2306 0 -2.0 1e-06 
0.0 -1.2305 0 -2.0 1e-06 
0.0 -1.2304 0 -2.0 1e-06 
0.0 -1.2303 0 -2.0 1e-06 
0.0 -1.2302 0 -2.0 1e-06 
0.0 -1.2301 0 -2.0 1e-06 
0.0 -1.23 0 -2.0 1e-06 
0.0 -1.2299 0 -2.0 1e-06 
0.0 -1.2298 0 -2.0 1e-06 
0.0 -1.2297 0 -2.0 1e-06 
0.0 -1.2296 0 -2.0 1e-06 
0.0 -1.2295 0 -2.0 1e-06 
0.0 -1.2294 0 -2.0 1e-06 
0.0 -1.2293 0 -2.0 1e-06 
0.0 -1.2292 0 -2.0 1e-06 
0.0 -1.2291 0 -2.0 1e-06 
0.0 -1.229 0 -2.0 1e-06 
0.0 -1.2289 0 -2.0 1e-06 
0.0 -1.2288 0 -2.0 1e-06 
0.0 -1.2287 0 -2.0 1e-06 
0.0 -1.2286 0 -2.0 1e-06 
0.0 -1.2285 0 -2.0 1e-06 
0.0 -1.2284 0 -2.0 1e-06 
0.0 -1.2283 0 -2.0 1e-06 
0.0 -1.2282 0 -2.0 1e-06 
0.0 -1.2281 0 -2.0 1e-06 
0.0 -1.228 0 -2.0 1e-06 
0.0 -1.2279 0 -2.0 1e-06 
0.0 -1.2278 0 -2.0 1e-06 
0.0 -1.2277 0 -2.0 1e-06 
0.0 -1.2276 0 -2.0 1e-06 
0.0 -1.2275 0 -2.0 1e-06 
0.0 -1.2274 0 -2.0 1e-06 
0.0 -1.2273 0 -2.0 1e-06 
0.0 -1.2272 0 -2.0 1e-06 
0.0 -1.2271 0 -2.0 1e-06 
0.0 -1.227 0 -2.0 1e-06 
0.0 -1.2269 0 -2.0 1e-06 
0.0 -1.2268 0 -2.0 1e-06 
0.0 -1.2267 0 -2.0 1e-06 
0.0 -1.2266 0 -2.0 1e-06 
0.0 -1.2265 0 -2.0 1e-06 
0.0 -1.2264 0 -2.0 1e-06 
0.0 -1.2263 0 -2.0 1e-06 
0.0 -1.2262 0 -2.0 1e-06 
0.0 -1.2261 0 -2.0 1e-06 
0.0 -1.226 0 -2.0 1e-06 
0.0 -1.2259 0 -2.0 1e-06 
0.0 -1.2258 0 -2.0 1e-06 
0.0 -1.2257 0 -2.0 1e-06 
0.0 -1.2256 0 -2.0 1e-06 
0.0 -1.2255 0 -2.0 1e-06 
0.0 -1.2254 0 -2.0 1e-06 
0.0 -1.2253 0 -2.0 1e-06 
0.0 -1.2252 0 -2.0 1e-06 
0.0 -1.2251 0 -2.0 1e-06 
0.0 -1.225 0 -2.0 1e-06 
0.0 -1.2249 0 -2.0 1e-06 
0.0 -1.2248 0 -2.0 1e-06 
0.0 -1.2247 0 -2.0 1e-06 
0.0 -1.2246 0 -2.0 1e-06 
0.0 -1.2245 0 -2.0 1e-06 
0.0 -1.2244 0 -2.0 1e-06 
0.0 -1.2243 0 -2.0 1e-06 
0.0 -1.2242 0 -2.0 1e-06 
0.0 -1.2241 0 -2.0 1e-06 
0.0 -1.224 0 -2.0 1e-06 
0.0 -1.2239 0 -2.0 1e-06 
0.0 -1.2238 0 -2.0 1e-06 
0.0 -1.2237 0 -2.0 1e-06 
0.0 -1.2236 0 -2.0 1e-06 
0.0 -1.2235 0 -2.0 1e-06 
0.0 -1.2234 0 -2.0 1e-06 
0.0 -1.2233 0 -2.0 1e-06 
0.0 -1.2232 0 -2.0 1e-06 
0.0 -1.2231 0 -2.0 1e-06 
0.0 -1.223 0 -2.0 1e-06 
0.0 -1.2229 0 -2.0 1e-06 
0.0 -1.2228 0 -2.0 1e-06 
0.0 -1.2227 0 -2.0 1e-06 
0.0 -1.2226 0 -2.0 1e-06 
0.0 -1.2225 0 -2.0 1e-06 
0.0 -1.2224 0 -2.0 1e-06 
0.0 -1.2223 0 -2.0 1e-06 
0.0 -1.2222 0 -2.0 1e-06 
0.0 -1.2221 0 -2.0 1e-06 
0.0 -1.222 0 -2.0 1e-06 
0.0 -1.2219 0 -2.0 1e-06 
0.0 -1.2218 0 -2.0 1e-06 
0.0 -1.2217 0 -2.0 1e-06 
0.0 -1.2216 0 -2.0 1e-06 
0.0 -1.2215 0 -2.0 1e-06 
0.0 -1.2214 0 -2.0 1e-06 
0.0 -1.2213 0 -2.0 1e-06 
0.0 -1.2212 0 -2.0 1e-06 
0.0 -1.2211 0 -2.0 1e-06 
0.0 -1.221 0 -2.0 1e-06 
0.0 -1.2209 0 -2.0 1e-06 
0.0 -1.2208 0 -2.0 1e-06 
0.0 -1.2207 0 -2.0 1e-06 
0.0 -1.2206 0 -2.0 1e-06 
0.0 -1.2205 0 -2.0 1e-06 
0.0 -1.2204 0 -2.0 1e-06 
0.0 -1.2203 0 -2.0 1e-06 
0.0 -1.2202 0 -2.0 1e-06 
0.0 -1.2201 0 -2.0 1e-06 
0.0 -1.22 0 -2.0 1e-06 
0.0 -1.2199 0 -2.0 1e-06 
0.0 -1.2198 0 -2.0 1e-06 
0.0 -1.2197 0 -2.0 1e-06 
0.0 -1.2196 0 -2.0 1e-06 
0.0 -1.2195 0 -2.0 1e-06 
0.0 -1.2194 0 -2.0 1e-06 
0.0 -1.2193 0 -2.0 1e-06 
0.0 -1.2192 0 -2.0 1e-06 
0.0 -1.2191 0 -2.0 1e-06 
0.0 -1.219 0 -2.0 1e-06 
0.0 -1.2189 0 -2.0 1e-06 
0.0 -1.2188 0 -2.0 1e-06 
0.0 -1.2187 0 -2.0 1e-06 
0.0 -1.2186 0 -2.0 1e-06 
0.0 -1.2185 0 -2.0 1e-06 
0.0 -1.2184 0 -2.0 1e-06 
0.0 -1.2183 0 -2.0 1e-06 
0.0 -1.2182 0 -2.0 1e-06 
0.0 -1.2181 0 -2.0 1e-06 
0.0 -1.218 0 -2.0 1e-06 
0.0 -1.2179 0 -2.0 1e-06 
0.0 -1.2178 0 -2.0 1e-06 
0.0 -1.2177 0 -2.0 1e-06 
0.0 -1.2176 0 -2.0 1e-06 
0.0 -1.2175 0 -2.0 1e-06 
0.0 -1.2174 0 -2.0 1e-06 
0.0 -1.2173 0 -2.0 1e-06 
0.0 -1.2172 0 -2.0 1e-06 
0.0 -1.2171 0 -2.0 1e-06 
0.0 -1.217 0 -2.0 1e-06 
0.0 -1.2169 0 -2.0 1e-06 
0.0 -1.2168 0 -2.0 1e-06 
0.0 -1.2167 0 -2.0 1e-06 
0.0 -1.2166 0 -2.0 1e-06 
0.0 -1.2165 0 -2.0 1e-06 
0.0 -1.2164 0 -2.0 1e-06 
0.0 -1.2163 0 -2.0 1e-06 
0.0 -1.2162 0 -2.0 1e-06 
0.0 -1.2161 0 -2.0 1e-06 
0.0 -1.216 0 -2.0 1e-06 
0.0 -1.2159 0 -2.0 1e-06 
0.0 -1.2158 0 -2.0 1e-06 
0.0 -1.2157 0 -2.0 1e-06 
0.0 -1.2156 0 -2.0 1e-06 
0.0 -1.2155 0 -2.0 1e-06 
0.0 -1.2154 0 -2.0 1e-06 
0.0 -1.2153 0 -2.0 1e-06 
0.0 -1.2152 0 -2.0 1e-06 
0.0 -1.2151 0 -2.0 1e-06 
0.0 -1.215 0 -2.0 1e-06 
0.0 -1.2149 0 -2.0 1e-06 
0.0 -1.2148 0 -2.0 1e-06 
0.0 -1.2147 0 -2.0 1e-06 
0.0 -1.2146 0 -2.0 1e-06 
0.0 -1.2145 0 -2.0 1e-06 
0.0 -1.2144 0 -2.0 1e-06 
0.0 -1.2143 0 -2.0 1e-06 
0.0 -1.2142 0 -2.0 1e-06 
0.0 -1.2141 0 -2.0 1e-06 
0.0 -1.214 0 -2.0 1e-06 
0.0 -1.2139 0 -2.0 1e-06 
0.0 -1.2138 0 -2.0 1e-06 
0.0 -1.2137 0 -2.0 1e-06 
0.0 -1.2136 0 -2.0 1e-06 
0.0 -1.2135 0 -2.0 1e-06 
0.0 -1.2134 0 -2.0 1e-06 
0.0 -1.2133 0 -2.0 1e-06 
0.0 -1.2132 0 -2.0 1e-06 
0.0 -1.2131 0 -2.0 1e-06 
0.0 -1.213 0 -2.0 1e-06 
0.0 -1.2129 0 -2.0 1e-06 
0.0 -1.2128 0 -2.0 1e-06 
0.0 -1.2127 0 -2.0 1e-06 
0.0 -1.2126 0 -2.0 1e-06 
0.0 -1.2125 0 -2.0 1e-06 
0.0 -1.2124 0 -2.0 1e-06 
0.0 -1.2123 0 -2.0 1e-06 
0.0 -1.2122 0 -2.0 1e-06 
0.0 -1.2121 0 -2.0 1e-06 
0.0 -1.212 0 -2.0 1e-06 
0.0 -1.2119 0 -2.0 1e-06 
0.0 -1.2118 0 -2.0 1e-06 
0.0 -1.2117 0 -2.0 1e-06 
0.0 -1.2116 0 -2.0 1e-06 
0.0 -1.2115 0 -2.0 1e-06 
0.0 -1.2114 0 -2.0 1e-06 
0.0 -1.2113 0 -2.0 1e-06 
0.0 -1.2112 0 -2.0 1e-06 
0.0 -1.2111 0 -2.0 1e-06 
0.0 -1.211 0 -2.0 1e-06 
0.0 -1.2109 0 -2.0 1e-06 
0.0 -1.2108 0 -2.0 1e-06 
0.0 -1.2107 0 -2.0 1e-06 
0.0 -1.2106 0 -2.0 1e-06 
0.0 -1.2105 0 -2.0 1e-06 
0.0 -1.2104 0 -2.0 1e-06 
0.0 -1.2103 0 -2.0 1e-06 
0.0 -1.2102 0 -2.0 1e-06 
0.0 -1.2101 0 -2.0 1e-06 
0.0 -1.21 0 -2.0 1e-06 
0.0 -1.2099 0 -2.0 1e-06 
0.0 -1.2098 0 -2.0 1e-06 
0.0 -1.2097 0 -2.0 1e-06 
0.0 -1.2096 0 -2.0 1e-06 
0.0 -1.2095 0 -2.0 1e-06 
0.0 -1.2094 0 -2.0 1e-06 
0.0 -1.2093 0 -2.0 1e-06 
0.0 -1.2092 0 -2.0 1e-06 
0.0 -1.2091 0 -2.0 1e-06 
0.0 -1.209 0 -2.0 1e-06 
0.0 -1.2089 0 -2.0 1e-06 
0.0 -1.2088 0 -2.0 1e-06 
0.0 -1.2087 0 -2.0 1e-06 
0.0 -1.2086 0 -2.0 1e-06 
0.0 -1.2085 0 -2.0 1e-06 
0.0 -1.2084 0 -2.0 1e-06 
0.0 -1.2083 0 -2.0 1e-06 
0.0 -1.2082 0 -2.0 1e-06 
0.0 -1.2081 0 -2.0 1e-06 
0.0 -1.208 0 -2.0 1e-06 
0.0 -1.2079 0 -2.0 1e-06 
0.0 -1.2078 0 -2.0 1e-06 
0.0 -1.2077 0 -2.0 1e-06 
0.0 -1.2076 0 -2.0 1e-06 
0.0 -1.2075 0 -2.0 1e-06 
0.0 -1.2074 0 -2.0 1e-06 
0.0 -1.2073 0 -2.0 1e-06 
0.0 -1.2072 0 -2.0 1e-06 
0.0 -1.2071 0 -2.0 1e-06 
0.0 -1.207 0 -2.0 1e-06 
0.0 -1.2069 0 -2.0 1e-06 
0.0 -1.2068 0 -2.0 1e-06 
0.0 -1.2067 0 -2.0 1e-06 
0.0 -1.2066 0 -2.0 1e-06 
0.0 -1.2065 0 -2.0 1e-06 
0.0 -1.2064 0 -2.0 1e-06 
0.0 -1.2063 0 -2.0 1e-06 
0.0 -1.2062 0 -2.0 1e-06 
0.0 -1.2061 0 -2.0 1e-06 
0.0 -1.206 0 -2.0 1e-06 
0.0 -1.2059 0 -2.0 1e-06 
0.0 -1.2058 0 -2.0 1e-06 
0.0 -1.2057 0 -2.0 1e-06 
0.0 -1.2056 0 -2.0 1e-06 
0.0 -1.2055 0 -2.0 1e-06 
0.0 -1.2054 0 -2.0 1e-06 
0.0 -1.2053 0 -2.0 1e-06 
0.0 -1.2052 0 -2.0 1e-06 
0.0 -1.2051 0 -2.0 1e-06 
0.0 -1.205 0 -2.0 1e-06 
0.0 -1.2049 0 -2.0 1e-06 
0.0 -1.2048 0 -2.0 1e-06 
0.0 -1.2047 0 -2.0 1e-06 
0.0 -1.2046 0 -2.0 1e-06 
0.0 -1.2045 0 -2.0 1e-06 
0.0 -1.2044 0 -2.0 1e-06 
0.0 -1.2043 0 -2.0 1e-06 
0.0 -1.2042 0 -2.0 1e-06 
0.0 -1.2041 0 -2.0 1e-06 
0.0 -1.204 0 -2.0 1e-06 
0.0 -1.2039 0 -2.0 1e-06 
0.0 -1.2038 0 -2.0 1e-06 
0.0 -1.2037 0 -2.0 1e-06 
0.0 -1.2036 0 -2.0 1e-06 
0.0 -1.2035 0 -2.0 1e-06 
0.0 -1.2034 0 -2.0 1e-06 
0.0 -1.2033 0 -2.0 1e-06 
0.0 -1.2032 0 -2.0 1e-06 
0.0 -1.2031 0 -2.0 1e-06 
0.0 -1.203 0 -2.0 1e-06 
0.0 -1.2029 0 -2.0 1e-06 
0.0 -1.2028 0 -2.0 1e-06 
0.0 -1.2027 0 -2.0 1e-06 
0.0 -1.2026 0 -2.0 1e-06 
0.0 -1.2025 0 -2.0 1e-06 
0.0 -1.2024 0 -2.0 1e-06 
0.0 -1.2023 0 -2.0 1e-06 
0.0 -1.2022 0 -2.0 1e-06 
0.0 -1.2021 0 -2.0 1e-06 
0.0 -1.202 0 -2.0 1e-06 
0.0 -1.2019 0 -2.0 1e-06 
0.0 -1.2018 0 -2.0 1e-06 
0.0 -1.2017 0 -2.0 1e-06 
0.0 -1.2016 0 -2.0 1e-06 
0.0 -1.2015 0 -2.0 1e-06 
0.0 -1.2014 0 -2.0 1e-06 
0.0 -1.2013 0 -2.0 1e-06 
0.0 -1.2012 0 -2.0 1e-06 
0.0 -1.2011 0 -2.0 1e-06 
0.0 -1.201 0 -2.0 1e-06 
0.0 -1.2009 0 -2.0 1e-06 
0.0 -1.2008 0 -2.0 1e-06 
0.0 -1.2007 0 -2.0 1e-06 
0.0 -1.2006 0 -2.0 1e-06 
0.0 -1.2005 0 -2.0 1e-06 
0.0 -1.2004 0 -2.0 1e-06 
0.0 -1.2003 0 -2.0 1e-06 
0.0 -1.2002 0 -2.0 1e-06 
0.0 -1.2001 0 -2.0 1e-06 
0.0 -1.2 0 -2.0 1e-06 
0.0 -1.1999 0 -2.0 1e-06 
0.0 -1.1998 0 -2.0 1e-06 
0.0 -1.1997 0 -2.0 1e-06 
0.0 -1.1996 0 -2.0 1e-06 
0.0 -1.1995 0 -2.0 1e-06 
0.0 -1.1994 0 -2.0 1e-06 
0.0 -1.1993 0 -2.0 1e-06 
0.0 -1.1992 0 -2.0 1e-06 
0.0 -1.1991 0 -2.0 1e-06 
0.0 -1.199 0 -2.0 1e-06 
0.0 -1.1989 0 -2.0 1e-06 
0.0 -1.1988 0 -2.0 1e-06 
0.0 -1.1987 0 -2.0 1e-06 
0.0 -1.1986 0 -2.0 1e-06 
0.0 -1.1985 0 -2.0 1e-06 
0.0 -1.1984 0 -2.0 1e-06 
0.0 -1.1983 0 -2.0 1e-06 
0.0 -1.1982 0 -2.0 1e-06 
0.0 -1.1981 0 -2.0 1e-06 
0.0 -1.198 0 -2.0 1e-06 
0.0 -1.1979 0 -2.0 1e-06 
0.0 -1.1978 0 -2.0 1e-06 
0.0 -1.1977 0 -2.0 1e-06 
0.0 -1.1976 0 -2.0 1e-06 
0.0 -1.1975 0 -2.0 1e-06 
0.0 -1.1974 0 -2.0 1e-06 
0.0 -1.1973 0 -2.0 1e-06 
0.0 -1.1972 0 -2.0 1e-06 
0.0 -1.1971 0 -2.0 1e-06 
0.0 -1.197 0 -2.0 1e-06 
0.0 -1.1969 0 -2.0 1e-06 
0.0 -1.1968 0 -2.0 1e-06 
0.0 -1.1967 0 -2.0 1e-06 
0.0 -1.1966 0 -2.0 1e-06 
0.0 -1.1965 0 -2.0 1e-06 
0.0 -1.1964 0 -2.0 1e-06 
0.0 -1.1963 0 -2.0 1e-06 
0.0 -1.1962 0 -2.0 1e-06 
0.0 -1.1961 0 -2.0 1e-06 
0.0 -1.196 0 -2.0 1e-06 
0.0 -1.1959 0 -2.0 1e-06 
0.0 -1.1958 0 -2.0 1e-06 
0.0 -1.1957 0 -2.0 1e-06 
0.0 -1.1956 0 -2.0 1e-06 
0.0 -1.1955 0 -2.0 1e-06 
0.0 -1.1954 0 -2.0 1e-06 
0.0 -1.1953 0 -2.0 1e-06 
0.0 -1.1952 0 -2.0 1e-06 
0.0 -1.1951 0 -2.0 1e-06 
0.0 -1.195 0 -2.0 1e-06 
0.0 -1.1949 0 -2.0 1e-06 
0.0 -1.1948 0 -2.0 1e-06 
0.0 -1.1947 0 -2.0 1e-06 
0.0 -1.1946 0 -2.0 1e-06 
0.0 -1.1945 0 -2.0 1e-06 
0.0 -1.1944 0 -2.0 1e-06 
0.0 -1.1943 0 -2.0 1e-06 
0.0 -1.1942 0 -2.0 1e-06 
0.0 -1.1941 0 -2.0 1e-06 
0.0 -1.194 0 -2.0 1e-06 
0.0 -1.1939 0 -2.0 1e-06 
0.0 -1.1938 0 -2.0 1e-06 
0.0 -1.1937 0 -2.0 1e-06 
0.0 -1.1936 0 -2.0 1e-06 
0.0 -1.1935 0 -2.0 1e-06 
0.0 -1.1934 0 -2.0 1e-06 
0.0 -1.1933 0 -2.0 1e-06 
0.0 -1.1932 0 -2.0 1e-06 
0.0 -1.1931 0 -2.0 1e-06 
0.0 -1.193 0 -2.0 1e-06 
0.0 -1.1929 0 -2.0 1e-06 
0.0 -1.1928 0 -2.0 1e-06 
0.0 -1.1927 0 -2.0 1e-06 
0.0 -1.1926 0 -2.0 1e-06 
0.0 -1.1925 0 -2.0 1e-06 
0.0 -1.1924 0 -2.0 1e-06 
0.0 -1.1923 0 -2.0 1e-06 
0.0 -1.1922 0 -2.0 1e-06 
0.0 -1.1921 0 -2.0 1e-06 
0.0 -1.192 0 -2.0 1e-06 
0.0 -1.1919 0 -2.0 1e-06 
0.0 -1.1918 0 -2.0 1e-06 
0.0 -1.1917 0 -2.0 1e-06 
0.0 -1.1916 0 -2.0 1e-06 
0.0 -1.1915 0 -2.0 1e-06 
0.0 -1.1914 0 -2.0 1e-06 
0.0 -1.1913 0 -2.0 1e-06 
0.0 -1.1912 0 -2.0 1e-06 
0.0 -1.1911 0 -2.0 1e-06 
0.0 -1.191 0 -2.0 1e-06 
0.0 -1.1909 0 -2.0 1e-06 
0.0 -1.1908 0 -2.0 1e-06 
0.0 -1.1907 0 -2.0 1e-06 
0.0 -1.1906 0 -2.0 1e-06 
0.0 -1.1905 0 -2.0 1e-06 
0.0 -1.1904 0 -2.0 1e-06 
0.0 -1.1903 0 -2.0 1e-06 
0.0 -1.1902 0 -2.0 1e-06 
0.0 -1.1901 0 -2.0 1e-06 
0.0 -1.19 0 -2.0 1e-06 
0.0 -1.1899 0 -2.0 1e-06 
0.0 -1.1898 0 -2.0 1e-06 
0.0 -1.1897 0 -2.0 1e-06 
0.0 -1.1896 0 -2.0 1e-06 
0.0 -1.1895 0 -2.0 1e-06 
0.0 -1.1894 0 -2.0 1e-06 
0.0 -1.1893 0 -2.0 1e-06 
0.0 -1.1892 0 -2.0 1e-06 
0.0 -1.1891 0 -2.0 1e-06 
0.0 -1.189 0 -2.0 1e-06 
0.0 -1.1889 0 -2.0 1e-06 
0.0 -1.1888 0 -2.0 1e-06 
0.0 -1.1887 0 -2.0 1e-06 
0.0 -1.1886 0 -2.0 1e-06 
0.0 -1.1885 0 -2.0 1e-06 
0.0 -1.1884 0 -2.0 1e-06 
0.0 -1.1883 0 -2.0 1e-06 
0.0 -1.1882 0 -2.0 1e-06 
0.0 -1.1881 0 -2.0 1e-06 
0.0 -1.188 0 -2.0 1e-06 
0.0 -1.1879 0 -2.0 1e-06 
0.0 -1.1878 0 -2.0 1e-06 
0.0 -1.1877 0 -2.0 1e-06 
0.0 -1.1876 0 -2.0 1e-06 
0.0 -1.1875 0 -2.0 1e-06 
0.0 -1.1874 0 -2.0 1e-06 
0.0 -1.1873 0 -2.0 1e-06 
0.0 -1.1872 0 -2.0 1e-06 
0.0 -1.1871 0 -2.0 1e-06 
0.0 -1.187 0 -2.0 1e-06 
0.0 -1.1869 0 -2.0 1e-06 
0.0 -1.1868 0 -2.0 1e-06 
0.0 -1.1867 0 -2.0 1e-06 
0.0 -1.1866 0 -2.0 1e-06 
0.0 -1.1865 0 -2.0 1e-06 
0.0 -1.1864 0 -2.0 1e-06 
0.0 -1.1863 0 -2.0 1e-06 
0.0 -1.1862 0 -2.0 1e-06 
0.0 -1.1861 0 -2.0 1e-06 
0.0 -1.186 0 -2.0 1e-06 
0.0 -1.1859 0 -2.0 1e-06 
0.0 -1.1858 0 -2.0 1e-06 
0.0 -1.1857 0 -2.0 1e-06 
0.0 -1.1856 0 -2.0 1e-06 
0.0 -1.1855 0 -2.0 1e-06 
0.0 -1.1854 0 -2.0 1e-06 
0.0 -1.1853 0 -2.0 1e-06 
0.0 -1.1852 0 -2.0 1e-06 
0.0 -1.1851 0 -2.0 1e-06 
0.0 -1.185 0 -2.0 1e-06 
0.0 -1.1849 0 -2.0 1e-06 
0.0 -1.1848 0 -2.0 1e-06 
0.0 -1.1847 0 -2.0 1e-06 
0.0 -1.1846 0 -2.0 1e-06 
0.0 -1.1845 0 -2.0 1e-06 
0.0 -1.1844 0 -2.0 1e-06 
0.0 -1.1843 0 -2.0 1e-06 
0.0 -1.1842 0 -2.0 1e-06 
0.0 -1.1841 0 -2.0 1e-06 
0.0 -1.184 0 -2.0 1e-06 
0.0 -1.1839 0 -2.0 1e-06 
0.0 -1.1838 0 -2.0 1e-06 
0.0 -1.1837 0 -2.0 1e-06 
0.0 -1.1836 0 -2.0 1e-06 
0.0 -1.1835 0 -2.0 1e-06 
0.0 -1.1834 0 -2.0 1e-06 
0.0 -1.1833 0 -2.0 1e-06 
0.0 -1.1832 0 -2.0 1e-06 
0.0 -1.1831 0 -2.0 1e-06 
0.0 -1.183 0 -2.0 1e-06 
0.0 -1.1829 0 -2.0 1e-06 
0.0 -1.1828 0 -2.0 1e-06 
0.0 -1.1827 0 -2.0 1e-06 
0.0 -1.1826 0 -2.0 1e-06 
0.0 -1.1825 0 -2.0 1e-06 
0.0 -1.1824 0 -2.0 1e-06 
0.0 -1.1823 0 -2.0 1e-06 
0.0 -1.1822 0 -2.0 1e-06 
0.0 -1.1821 0 -2.0 1e-06 
0.0 -1.182 0 -2.0 1e-06 
0.0 -1.1819 0 -2.0 1e-06 
0.0 -1.1818 0 -2.0 1e-06 
0.0 -1.1817 0 -2.0 1e-06 
0.0 -1.1816 0 -2.0 1e-06 
0.0 -1.1815 0 -2.0 1e-06 
0.0 -1.1814 0 -2.0 1e-06 
0.0 -1.1813 0 -2.0 1e-06 
0.0 -1.1812 0 -2.0 1e-06 
0.0 -1.1811 0 -2.0 1e-06 
0.0 -1.181 0 -2.0 1e-06 
0.0 -1.1809 0 -2.0 1e-06 
0.0 -1.1808 0 -2.0 1e-06 
0.0 -1.1807 0 -2.0 1e-06 
0.0 -1.1806 0 -2.0 1e-06 
0.0 -1.1805 0 -2.0 1e-06 
0.0 -1.1804 0 -2.0 1e-06 
0.0 -1.1803 0 -2.0 1e-06 
0.0 -1.1802 0 -2.0 1e-06 
0.0 -1.1801 0 -2.0 1e-06 
0.0 -1.18 0 -2.0 1e-06 
0.0 -1.1799 0 -2.0 1e-06 
0.0 -1.1798 0 -2.0 1e-06 
0.0 -1.1797 0 -2.0 1e-06 
0.0 -1.1796 0 -2.0 1e-06 
0.0 -1.1795 0 -2.0 1e-06 
0.0 -1.1794 0 -2.0 1e-06 
0.0 -1.1793 0 -2.0 1e-06 
0.0 -1.1792 0 -2.0 1e-06 
0.0 -1.1791 0 -2.0 1e-06 
0.0 -1.179 0 -2.0 1e-06 
0.0 -1.1789 0 -2.0 1e-06 
0.0 -1.1788 0 -2.0 1e-06 
0.0 -1.1787 0 -2.0 1e-06 
0.0 -1.1786 0 -2.0 1e-06 
0.0 -1.1785 0 -2.0 1e-06 
0.0 -1.1784 0 -2.0 1e-06 
0.0 -1.1783 0 -2.0 1e-06 
0.0 -1.1782 0 -2.0 1e-06 
0.0 -1.1781 0 -2.0 1e-06 
0.0 -1.178 0 -2.0 1e-06 
0.0 -1.1779 0 -2.0 1e-06 
0.0 -1.1778 0 -2.0 1e-06 
0.0 -1.1777 0 -2.0 1e-06 
0.0 -1.1776 0 -2.0 1e-06 
0.0 -1.1775 0 -2.0 1e-06 
0.0 -1.1774 0 -2.0 1e-06 
0.0 -1.1773 0 -2.0 1e-06 
0.0 -1.1772 0 -2.0 1e-06 
0.0 -1.1771 0 -2.0 1e-06 
0.0 -1.177 0 -2.0 1e-06 
0.0 -1.1769 0 -2.0 1e-06 
0.0 -1.1768 0 -2.0 1e-06 
0.0 -1.1767 0 -2.0 1e-06 
0.0 -1.1766 0 -2.0 1e-06 
0.0 -1.1765 0 -2.0 1e-06 
0.0 -1.1764 0 -2.0 1e-06 
0.0 -1.1763 0 -2.0 1e-06 
0.0 -1.1762 0 -2.0 1e-06 
0.0 -1.1761 0 -2.0 1e-06 
0.0 -1.176 0 -2.0 1e-06 
0.0 -1.1759 0 -2.0 1e-06 
0.0 -1.1758 0 -2.0 1e-06 
0.0 -1.1757 0 -2.0 1e-06 
0.0 -1.1756 0 -2.0 1e-06 
0.0 -1.1755 0 -2.0 1e-06 
0.0 -1.1754 0 -2.0 1e-06 
0.0 -1.1753 0 -2.0 1e-06 
0.0 -1.1752 0 -2.0 1e-06 
0.0 -1.1751 0 -2.0 1e-06 
0.0 -1.175 0 -2.0 1e-06 
0.0 -1.1749 0 -2.0 1e-06 
0.0 -1.1748 0 -2.0 1e-06 
0.0 -1.1747 0 -2.0 1e-06 
0.0 -1.1746 0 -2.0 1e-06 
0.0 -1.1745 0 -2.0 1e-06 
0.0 -1.1744 0 -2.0 1e-06 
0.0 -1.1743 0 -2.0 1e-06 
0.0 -1.1742 0 -2.0 1e-06 
0.0 -1.1741 0 -2.0 1e-06 
0.0 -1.174 0 -2.0 1e-06 
0.0 -1.1739 0 -2.0 1e-06 
0.0 -1.1738 0 -2.0 1e-06 
0.0 -1.1737 0 -2.0 1e-06 
0.0 -1.1736 0 -2.0 1e-06 
0.0 -1.1735 0 -2.0 1e-06 
0.0 -1.1734 0 -2.0 1e-06 
0.0 -1.1733 0 -2.0 1e-06 
0.0 -1.1732 0 -2.0 1e-06 
0.0 -1.1731 0 -2.0 1e-06 
0.0 -1.173 0 -2.0 1e-06 
0.0 -1.1729 0 -2.0 1e-06 
0.0 -1.1728 0 -2.0 1e-06 
0.0 -1.1727 0 -2.0 1e-06 
0.0 -1.1726 0 -2.0 1e-06 
0.0 -1.1725 0 -2.0 1e-06 
0.0 -1.1724 0 -2.0 1e-06 
0.0 -1.1723 0 -2.0 1e-06 
0.0 -1.1722 0 -2.0 1e-06 
0.0 -1.1721 0 -2.0 1e-06 
0.0 -1.172 0 -2.0 1e-06 
0.0 -1.1719 0 -2.0 1e-06 
0.0 -1.1718 0 -2.0 1e-06 
0.0 -1.1717 0 -2.0 1e-06 
0.0 -1.1716 0 -2.0 1e-06 
0.0 -1.1715 0 -2.0 1e-06 
0.0 -1.1714 0 -2.0 1e-06 
0.0 -1.1713 0 -2.0 1e-06 
0.0 -1.1712 0 -2.0 1e-06 
0.0 -1.1711 0 -2.0 1e-06 
0.0 -1.171 0 -2.0 1e-06 
0.0 -1.1709 0 -2.0 1e-06 
0.0 -1.1708 0 -2.0 1e-06 
0.0 -1.1707 0 -2.0 1e-06 
0.0 -1.1706 0 -2.0 1e-06 
0.0 -1.1705 0 -2.0 1e-06 
0.0 -1.1704 0 -2.0 1e-06 
0.0 -1.1703 0 -2.0 1e-06 
0.0 -1.1702 0 -2.0 1e-06 
0.0 -1.1701 0 -2.0 1e-06 
0.0 -1.17 0 -2.0 1e-06 
0.0 -1.1699 0 -2.0 1e-06 
0.0 -1.1698 0 -2.0 1e-06 
0.0 -1.1697 0 -2.0 1e-06 
0.0 -1.1696 0 -2.0 1e-06 
0.0 -1.1695 0 -2.0 1e-06 
0.0 -1.1694 0 -2.0 1e-06 
0.0 -1.1693 0 -2.0 1e-06 
0.0 -1.1692 0 -2.0 1e-06 
0.0 -1.1691 0 -2.0 1e-06 
0.0 -1.169 0 -2.0 1e-06 
0.0 -1.1689 0 -2.0 1e-06 
0.0 -1.1688 0 -2.0 1e-06 
0.0 -1.1687 0 -2.0 1e-06 
0.0 -1.1686 0 -2.0 1e-06 
0.0 -1.1685 0 -2.0 1e-06 
0.0 -1.1684 0 -2.0 1e-06 
0.0 -1.1683 0 -2.0 1e-06 
0.0 -1.1682 0 -2.0 1e-06 
0.0 -1.1681 0 -2.0 1e-06 
0.0 -1.168 0 -2.0 1e-06 
0.0 -1.1679 0 -2.0 1e-06 
0.0 -1.1678 0 -2.0 1e-06 
0.0 -1.1677 0 -2.0 1e-06 
0.0 -1.1676 0 -2.0 1e-06 
0.0 -1.1675 0 -2.0 1e-06 
0.0 -1.1674 0 -2.0 1e-06 
0.0 -1.1673 0 -2.0 1e-06 
0.0 -1.1672 0 -2.0 1e-06 
0.0 -1.1671 0 -2.0 1e-06 
0.0 -1.167 0 -2.0 1e-06 
0.0 -1.1669 0 -2.0 1e-06 
0.0 -1.1668 0 -2.0 1e-06 
0.0 -1.1667 0 -2.0 1e-06 
0.0 -1.1666 0 -2.0 1e-06 
0.0 -1.1665 0 -2.0 1e-06 
0.0 -1.1664 0 -2.0 1e-06 
0.0 -1.1663 0 -2.0 1e-06 
0.0 -1.1662 0 -2.0 1e-06 
0.0 -1.1661 0 -2.0 1e-06 
0.0 -1.166 0 -2.0 1e-06 
0.0 -1.1659 0 -2.0 1e-06 
0.0 -1.1658 0 -2.0 1e-06 
0.0 -1.1657 0 -2.0 1e-06 
0.0 -1.1656 0 -2.0 1e-06 
0.0 -1.1655 0 -2.0 1e-06 
0.0 -1.1654 0 -2.0 1e-06 
0.0 -1.1653 0 -2.0 1e-06 
0.0 -1.1652 0 -2.0 1e-06 
0.0 -1.1651 0 -2.0 1e-06 
0.0 -1.165 0 -2.0 1e-06 
0.0 -1.1649 0 -2.0 1e-06 
0.0 -1.1648 0 -2.0 1e-06 
0.0 -1.1647 0 -2.0 1e-06 
0.0 -1.1646 0 -2.0 1e-06 
0.0 -1.1645 0 -2.0 1e-06 
0.0 -1.1644 0 -2.0 1e-06 
0.0 -1.1643 0 -2.0 1e-06 
0.0 -1.1642 0 -2.0 1e-06 
0.0 -1.1641 0 -2.0 1e-06 
0.0 -1.164 0 -2.0 1e-06 
0.0 -1.1639 0 -2.0 1e-06 
0.0 -1.1638 0 -2.0 1e-06 
0.0 -1.1637 0 -2.0 1e-06 
0.0 -1.1636 0 -2.0 1e-06 
0.0 -1.1635 0 -2.0 1e-06 
0.0 -1.1634 0 -2.0 1e-06 
0.0 -1.1633 0 -2.0 1e-06 
0.0 -1.1632 0 -2.0 1e-06 
0.0 -1.1631 0 -2.0 1e-06 
0.0 -1.163 0 -2.0 1e-06 
0.0 -1.1629 0 -2.0 1e-06 
0.0 -1.1628 0 -2.0 1e-06 
0.0 -1.1627 0 -2.0 1e-06 
0.0 -1.1626 0 -2.0 1e-06 
0.0 -1.1625 0 -2.0 1e-06 
0.0 -1.1624 0 -2.0 1e-06 
0.0 -1.1623 0 -2.0 1e-06 
0.0 -1.1622 0 -2.0 1e-06 
0.0 -1.1621 0 -2.0 1e-06 
0.0 -1.162 0 -2.0 1e-06 
0.0 -1.1619 0 -2.0 1e-06 
0.0 -1.1618 0 -2.0 1e-06 
0.0 -1.1617 0 -2.0 1e-06 
0.0 -1.1616 0 -2.0 1e-06 
0.0 -1.1615 0 -2.0 1e-06 
0.0 -1.1614 0 -2.0 1e-06 
0.0 -1.1613 0 -2.0 1e-06 
0.0 -1.1612 0 -2.0 1e-06 
0.0 -1.1611 0 -2.0 1e-06 
0.0 -1.161 0 -2.0 1e-06 
0.0 -1.1609 0 -2.0 1e-06 
0.0 -1.1608 0 -2.0 1e-06 
0.0 -1.1607 0 -2.0 1e-06 
0.0 -1.1606 0 -2.0 1e-06 
0.0 -1.1605 0 -2.0 1e-06 
0.0 -1.1604 0 -2.0 1e-06 
0.0 -1.1603 0 -2.0 1e-06 
0.0 -1.1602 0 -2.0 1e-06 
0.0 -1.1601 0 -2.0 1e-06 
0.0 -1.16 0 -2.0 1e-06 
0.0 -1.1599 0 -2.0 1e-06 
0.0 -1.1598 0 -2.0 1e-06 
0.0 -1.1597 0 -2.0 1e-06 
0.0 -1.1596 0 -2.0 1e-06 
0.0 -1.1595 0 -2.0 1e-06 
0.0 -1.1594 0 -2.0 1e-06 
0.0 -1.1593 0 -2.0 1e-06 
0.0 -1.1592 0 -2.0 1e-06 
0.0 -1.1591 0 -2.0 1e-06 
0.0 -1.159 0 -2.0 1e-06 
0.0 -1.1589 0 -2.0 1e-06 
0.0 -1.1588 0 -2.0 1e-06 
0.0 -1.1587 0 -2.0 1e-06 
0.0 -1.1586 0 -2.0 1e-06 
0.0 -1.1585 0 -2.0 1e-06 
0.0 -1.1584 0 -2.0 1e-06 
0.0 -1.1583 0 -2.0 1e-06 
0.0 -1.1582 0 -2.0 1e-06 
0.0 -1.1581 0 -2.0 1e-06 
0.0 -1.158 0 -2.0 1e-06 
0.0 -1.1579 0 -2.0 1e-06 
0.0 -1.1578 0 -2.0 1e-06 
0.0 -1.1577 0 -2.0 1e-06 
0.0 -1.1576 0 -2.0 1e-06 
0.0 -1.1575 0 -2.0 1e-06 
0.0 -1.1574 0 -2.0 1e-06 
0.0 -1.1573 0 -2.0 1e-06 
0.0 -1.1572 0 -2.0 1e-06 
0.0 -1.1571 0 -2.0 1e-06 
0.0 -1.157 0 -2.0 1e-06 
0.0 -1.1569 0 -2.0 1e-06 
0.0 -1.1568 0 -2.0 1e-06 
0.0 -1.1567 0 -2.0 1e-06 
0.0 -1.1566 0 -2.0 1e-06 
0.0 -1.1565 0 -2.0 1e-06 
0.0 -1.1564 0 -2.0 1e-06 
0.0 -1.1563 0 -2.0 1e-06 
0.0 -1.1562 0 -2.0 1e-06 
0.0 -1.1561 0 -2.0 1e-06 
0.0 -1.156 0 -2.0 1e-06 
0.0 -1.1559 0 -2.0 1e-06 
0.0 -1.1558 0 -2.0 1e-06 
0.0 -1.1557 0 -2.0 1e-06 
0.0 -1.1556 0 -2.0 1e-06 
0.0 -1.1555 0 -2.0 1e-06 
0.0 -1.1554 0 -2.0 1e-06 
0.0 -1.1553 0 -2.0 1e-06 
0.0 -1.1552 0 -2.0 1e-06 
0.0 -1.1551 0 -2.0 1e-06 
0.0 -1.155 0 -2.0 1e-06 
0.0 -1.1549 0 -2.0 1e-06 
0.0 -1.1548 0 -2.0 1e-06 
0.0 -1.1547 0 -2.0 1e-06 
0.0 -1.1546 0 -2.0 1e-06 
0.0 -1.1545 0 -2.0 1e-06 
0.0 -1.1544 0 -2.0 1e-06 
0.0 -1.1543 0 -2.0 1e-06 
0.0 -1.1542 0 -2.0 1e-06 
0.0 -1.1541 0 -2.0 1e-06 
0.0 -1.154 0 -2.0 1e-06 
0.0 -1.1539 0 -2.0 1e-06 
0.0 -1.1538 0 -2.0 1e-06 
0.0 -1.1537 0 -2.0 1e-06 
0.0 -1.1536 0 -2.0 1e-06 
0.0 -1.1535 0 -2.0 1e-06 
0.0 -1.1534 0 -2.0 1e-06 
0.0 -1.1533 0 -2.0 1e-06 
0.0 -1.1532 0 -2.0 1e-06 
0.0 -1.1531 0 -2.0 1e-06 
0.0 -1.153 0 -2.0 1e-06 
0.0 -1.1529 0 -2.0 1e-06 
0.0 -1.1528 0 -2.0 1e-06 
0.0 -1.1527 0 -2.0 1e-06 
0.0 -1.1526 0 -2.0 1e-06 
0.0 -1.1525 0 -2.0 1e-06 
0.0 -1.1524 0 -2.0 1e-06 
0.0 -1.1523 0 -2.0 1e-06 
0.0 -1.1522 0 -2.0 1e-06 
0.0 -1.1521 0 -2.0 1e-06 
0.0 -1.152 0 -2.0 1e-06 
0.0 -1.1519 0 -2.0 1e-06 
0.0 -1.1518 0 -2.0 1e-06 
0.0 -1.1517 0 -2.0 1e-06 
0.0 -1.1516 0 -2.0 1e-06 
0.0 -1.1515 0 -2.0 1e-06 
0.0 -1.1514 0 -2.0 1e-06 
0.0 -1.1513 0 -2.0 1e-06 
0.0 -1.1512 0 -2.0 1e-06 
0.0 -1.1511 0 -2.0 1e-06 
0.0 -1.151 0 -2.0 1e-06 
0.0 -1.1509 0 -2.0 1e-06 
0.0 -1.1508 0 -2.0 1e-06 
0.0 -1.1507 0 -2.0 1e-06 
0.0 -1.1506 0 -2.0 1e-06 
0.0 -1.1505 0 -2.0 1e-06 
0.0 -1.1504 0 -2.0 1e-06 
0.0 -1.1503 0 -2.0 1e-06 
0.0 -1.1502 0 -2.0 1e-06 
0.0 -1.1501 0 -2.0 1e-06 
0.0 -1.15 0 -2.0 1e-06 
0.0 -1.1499 0 -2.0 1e-06 
0.0 -1.1498 0 -2.0 1e-06 
0.0 -1.1497 0 -2.0 1e-06 
0.0 -1.1496 0 -2.0 1e-06 
0.0 -1.1495 0 -2.0 1e-06 
0.0 -1.1494 0 -2.0 1e-06 
0.0 -1.1493 0 -2.0 1e-06 
0.0 -1.1492 0 -2.0 1e-06 
0.0 -1.1491 0 -2.0 1e-06 
0.0 -1.149 0 -2.0 1e-06 
0.0 -1.1489 0 -2.0 1e-06 
0.0 -1.1488 0 -2.0 1e-06 
0.0 -1.1487 0 -2.0 1e-06 
0.0 -1.1486 0 -2.0 1e-06 
0.0 -1.1485 0 -2.0 1e-06 
0.0 -1.1484 0 -2.0 1e-06 
0.0 -1.1483 0 -2.0 1e-06 
0.0 -1.1482 0 -2.0 1e-06 
0.0 -1.1481 0 -2.0 1e-06 
0.0 -1.148 0 -2.0 1e-06 
0.0 -1.1479 0 -2.0 1e-06 
0.0 -1.1478 0 -2.0 1e-06 
0.0 -1.1477 0 -2.0 1e-06 
0.0 -1.1476 0 -2.0 1e-06 
0.0 -1.1475 0 -2.0 1e-06 
0.0 -1.1474 0 -2.0 1e-06 
0.0 -1.1473 0 -2.0 1e-06 
0.0 -1.1472 0 -2.0 1e-06 
0.0 -1.1471 0 -2.0 1e-06 
0.0 -1.147 0 -2.0 1e-06 
0.0 -1.1469 0 -2.0 1e-06 
0.0 -1.1468 0 -2.0 1e-06 
0.0 -1.1467 0 -2.0 1e-06 
0.0 -1.1466 0 -2.0 1e-06 
0.0 -1.1465 0 -2.0 1e-06 
0.0 -1.1464 0 -2.0 1e-06 
0.0 -1.1463 0 -2.0 1e-06 
0.0 -1.1462 0 -2.0 1e-06 
0.0 -1.1461 0 -2.0 1e-06 
0.0 -1.146 0 -2.0 1e-06 
0.0 -1.1459 0 -2.0 1e-06 
0.0 -1.1458 0 -2.0 1e-06 
0.0 -1.1457 0 -2.0 1e-06 
0.0 -1.1456 0 -2.0 1e-06 
0.0 -1.1455 0 -2.0 1e-06 
0.0 -1.1454 0 -2.0 1e-06 
0.0 -1.1453 0 -2.0 1e-06 
0.0 -1.1452 0 -2.0 1e-06 
0.0 -1.1451 0 -2.0 1e-06 
0.0 -1.145 0 -2.0 1e-06 
0.0 -1.1449 0 -2.0 1e-06 
0.0 -1.1448 0 -2.0 1e-06 
0.0 -1.1447 0 -2.0 1e-06 
0.0 -1.1446 0 -2.0 1e-06 
0.0 -1.1445 0 -2.0 1e-06 
0.0 -1.1444 0 -2.0 1e-06 
0.0 -1.1443 0 -2.0 1e-06 
0.0 -1.1442 0 -2.0 1e-06 
0.0 -1.1441 0 -2.0 1e-06 
0.0 -1.144 0 -2.0 1e-06 
0.0 -1.1439 0 -2.0 1e-06 
0.0 -1.1438 0 -2.0 1e-06 
0.0 -1.1437 0 -2.0 1e-06 
0.0 -1.1436 0 -2.0 1e-06 
0.0 -1.1435 0 -2.0 1e-06 
0.0 -1.1434 0 -2.0 1e-06 
0.0 -1.1433 0 -2.0 1e-06 
0.0 -1.1432 0 -2.0 1e-06 
0.0 -1.1431 0 -2.0 1e-06 
0.0 -1.143 0 -2.0 1e-06 
0.0 -1.1429 0 -2.0 1e-06 
0.0 -1.1428 0 -2.0 1e-06 
0.0 -1.1427 0 -2.0 1e-06 
0.0 -1.1426 0 -2.0 1e-06 
0.0 -1.1425 0 -2.0 1e-06 
0.0 -1.1424 0 -2.0 1e-06 
0.0 -1.1423 0 -2.0 1e-06 
0.0 -1.1422 0 -2.0 1e-06 
0.0 -1.1421 0 -2.0 1e-06 
0.0 -1.142 0 -2.0 1e-06 
0.0 -1.1419 0 -2.0 1e-06 
0.0 -1.1418 0 -2.0 1e-06 
0.0 -1.1417 0 -2.0 1e-06 
0.0 -1.1416 0 -2.0 1e-06 
0.0 -1.1415 0 -2.0 1e-06 
0.0 -1.1414 0 -2.0 1e-06 
0.0 -1.1413 0 -2.0 1e-06 
0.0 -1.1412 0 -2.0 1e-06 
0.0 -1.1411 0 -2.0 1e-06 
0.0 -1.141 0 -2.0 1e-06 
0.0 -1.1409 0 -2.0 1e-06 
0.0 -1.1408 0 -2.0 1e-06 
0.0 -1.1407 0 -2.0 1e-06 
0.0 -1.1406 0 -2.0 1e-06 
0.0 -1.1405 0 -2.0 1e-06 
0.0 -1.1404 0 -2.0 1e-06 
0.0 -1.1403 0 -2.0 1e-06 
0.0 -1.1402 0 -2.0 1e-06 
0.0 -1.1401 0 -2.0 1e-06 
0.0 -1.14 0 -2.0 1e-06 
0.0 -1.1399 0 -2.0 1e-06 
0.0 -1.1398 0 -2.0 1e-06 
0.0 -1.1397 0 -2.0 1e-06 
0.0 -1.1396 0 -2.0 1e-06 
0.0 -1.1395 0 -2.0 1e-06 
0.0 -1.1394 0 -2.0 1e-06 
0.0 -1.1393 0 -2.0 1e-06 
0.0 -1.1392 0 -2.0 1e-06 
0.0 -1.1391 0 -2.0 1e-06 
0.0 -1.139 0 -2.0 1e-06 
0.0 -1.1389 0 -2.0 1e-06 
0.0 -1.1388 0 -2.0 1e-06 
0.0 -1.1387 0 -2.0 1e-06 
0.0 -1.1386 0 -2.0 1e-06 
0.0 -1.1385 0 -2.0 1e-06 
0.0 -1.1384 0 -2.0 1e-06 
0.0 -1.1383 0 -2.0 1e-06 
0.0 -1.1382 0 -2.0 1e-06 
0.0 -1.1381 0 -2.0 1e-06 
0.0 -1.138 0 -2.0 1e-06 
0.0 -1.1379 0 -2.0 1e-06 
0.0 -1.1378 0 -2.0 1e-06 
0.0 -1.1377 0 -2.0 1e-06 
0.0 -1.1376 0 -2.0 1e-06 
0.0 -1.1375 0 -2.0 1e-06 
0.0 -1.1374 0 -2.0 1e-06 
0.0 -1.1373 0 -2.0 1e-06 
0.0 -1.1372 0 -2.0 1e-06 
0.0 -1.1371 0 -2.0 1e-06 
0.0 -1.137 0 -2.0 1e-06 
0.0 -1.1369 0 -2.0 1e-06 
0.0 -1.1368 0 -2.0 1e-06 
0.0 -1.1367 0 -2.0 1e-06 
0.0 -1.1366 0 -2.0 1e-06 
0.0 -1.1365 0 -2.0 1e-06 
0.0 -1.1364 0 -2.0 1e-06 
0.0 -1.1363 0 -2.0 1e-06 
0.0 -1.1362 0 -2.0 1e-06 
0.0 -1.1361 0 -2.0 1e-06 
0.0 -1.136 0 -2.0 1e-06 
0.0 -1.1359 0 -2.0 1e-06 
0.0 -1.1358 0 -2.0 1e-06 
0.0 -1.1357 0 -2.0 1e-06 
0.0 -1.1356 0 -2.0 1e-06 
0.0 -1.1355 0 -2.0 1e-06 
0.0 -1.1354 0 -2.0 1e-06 
0.0 -1.1353 0 -2.0 1e-06 
0.0 -1.1352 0 -2.0 1e-06 
0.0 -1.1351 0 -2.0 1e-06 
0.0 -1.135 0 -2.0 1e-06 
0.0 -1.1349 0 -2.0 1e-06 
0.0 -1.1348 0 -2.0 1e-06 
0.0 -1.1347 0 -2.0 1e-06 
0.0 -1.1346 0 -2.0 1e-06 
0.0 -1.1345 0 -2.0 1e-06 
0.0 -1.1344 0 -2.0 1e-06 
0.0 -1.1343 0 -2.0 1e-06 
0.0 -1.1342 0 -2.0 1e-06 
0.0 -1.1341 0 -2.0 1e-06 
0.0 -1.134 0 -2.0 1e-06 
0.0 -1.1339 0 -2.0 1e-06 
0.0 -1.1338 0 -2.0 1e-06 
0.0 -1.1337 0 -2.0 1e-06 
0.0 -1.1336 0 -2.0 1e-06 
0.0 -1.1335 0 -2.0 1e-06 
0.0 -1.1334 0 -2.0 1e-06 
0.0 -1.1333 0 -2.0 1e-06 
0.0 -1.1332 0 -2.0 1e-06 
0.0 -1.1331 0 -2.0 1e-06 
0.0 -1.133 0 -2.0 1e-06 
0.0 -1.1329 0 -2.0 1e-06 
0.0 -1.1328 0 -2.0 1e-06 
0.0 -1.1327 0 -2.0 1e-06 
0.0 -1.1326 0 -2.0 1e-06 
0.0 -1.1325 0 -2.0 1e-06 
0.0 -1.1324 0 -2.0 1e-06 
0.0 -1.1323 0 -2.0 1e-06 
0.0 -1.1322 0 -2.0 1e-06 
0.0 -1.1321 0 -2.0 1e-06 
0.0 -1.132 0 -2.0 1e-06 
0.0 -1.1319 0 -2.0 1e-06 
0.0 -1.1318 0 -2.0 1e-06 
0.0 -1.1317 0 -2.0 1e-06 
0.0 -1.1316 0 -2.0 1e-06 
0.0 -1.1315 0 -2.0 1e-06 
0.0 -1.1314 0 -2.0 1e-06 
0.0 -1.1313 0 -2.0 1e-06 
0.0 -1.1312 0 -2.0 1e-06 
0.0 -1.1311 0 -2.0 1e-06 
0.0 -1.131 0 -2.0 1e-06 
0.0 -1.1309 0 -2.0 1e-06 
0.0 -1.1308 0 -2.0 1e-06 
0.0 -1.1307 0 -2.0 1e-06 
0.0 -1.1306 0 -2.0 1e-06 
0.0 -1.1305 0 -2.0 1e-06 
0.0 -1.1304 0 -2.0 1e-06 
0.0 -1.1303 0 -2.0 1e-06 
0.0 -1.1302 0 -2.0 1e-06 
0.0 -1.1301 0 -2.0 1e-06 
0.0 -1.13 0 -2.0 1e-06 
0.0 -1.1299 0 -2.0 1e-06 
0.0 -1.1298 0 -2.0 1e-06 
0.0 -1.1297 0 -2.0 1e-06 
0.0 -1.1296 0 -2.0 1e-06 
0.0 -1.1295 0 -2.0 1e-06 
0.0 -1.1294 0 -2.0 1e-06 
0.0 -1.1293 0 -2.0 1e-06 
0.0 -1.1292 0 -2.0 1e-06 
0.0 -1.1291 0 -2.0 1e-06 
0.0 -1.129 0 -2.0 1e-06 
0.0 -1.1289 0 -2.0 1e-06 
0.0 -1.1288 0 -2.0 1e-06 
0.0 -1.1287 0 -2.0 1e-06 
0.0 -1.1286 0 -2.0 1e-06 
0.0 -1.1285 0 -2.0 1e-06 
0.0 -1.1284 0 -2.0 1e-06 
0.0 -1.1283 0 -2.0 1e-06 
0.0 -1.1282 0 -2.0 1e-06 
0.0 -1.1281 0 -2.0 1e-06 
0.0 -1.128 0 -2.0 1e-06 
0.0 -1.1279 0 -2.0 1e-06 
0.0 -1.1278 0 -2.0 1e-06 
0.0 -1.1277 0 -2.0 1e-06 
0.0 -1.1276 0 -2.0 1e-06 
0.0 -1.1275 0 -2.0 1e-06 
0.0 -1.1274 0 -2.0 1e-06 
0.0 -1.1273 0 -2.0 1e-06 
0.0 -1.1272 0 -2.0 1e-06 
0.0 -1.1271 0 -2.0 1e-06 
0.0 -1.127 0 -2.0 1e-06 
0.0 -1.1269 0 -2.0 1e-06 
0.0 -1.1268 0 -2.0 1e-06 
0.0 -1.1267 0 -2.0 1e-06 
0.0 -1.1266 0 -2.0 1e-06 
0.0 -1.1265 0 -2.0 1e-06 
0.0 -1.1264 0 -2.0 1e-06 
0.0 -1.1263 0 -2.0 1e-06 
0.0 -1.1262 0 -2.0 1e-06 
0.0 -1.1261 0 -2.0 1e-06 
0.0 -1.126 0 -2.0 1e-06 
0.0 -1.1259 0 -2.0 1e-06 
0.0 -1.1258 0 -2.0 1e-06 
0.0 -1.1257 0 -2.0 1e-06 
0.0 -1.1256 0 -2.0 1e-06 
0.0 -1.1255 0 -2.0 1e-06 
0.0 -1.1254 0 -2.0 1e-06 
0.0 -1.1253 0 -2.0 1e-06 
0.0 -1.1252 0 -2.0 1e-06 
0.0 -1.1251 0 -2.0 1e-06 
0.0 -1.125 0 -2.0 1e-06 
0.0 -1.1249 0 -2.0 1e-06 
0.0 -1.1248 0 -2.0 1e-06 
0.0 -1.1247 0 -2.0 1e-06 
0.0 -1.1246 0 -2.0 1e-06 
0.0 -1.1245 0 -2.0 1e-06 
0.0 -1.1244 0 -2.0 1e-06 
0.0 -1.1243 0 -2.0 1e-06 
0.0 -1.1242 0 -2.0 1e-06 
0.0 -1.1241 0 -2.0 1e-06 
0.0 -1.124 0 -2.0 1e-06 
0.0 -1.1239 0 -2.0 1e-06 
0.0 -1.1238 0 -2.0 1e-06 
0.0 -1.1237 0 -2.0 1e-06 
0.0 -1.1236 0 -2.0 1e-06 
0.0 -1.1235 0 -2.0 1e-06 
0.0 -1.1234 0 -2.0 1e-06 
0.0 -1.1233 0 -2.0 1e-06 
0.0 -1.1232 0 -2.0 1e-06 
0.0 -1.1231 0 -2.0 1e-06 
0.0 -1.123 0 -2.0 1e-06 
0.0 -1.1229 0 -2.0 1e-06 
0.0 -1.1228 0 -2.0 1e-06 
0.0 -1.1227 0 -2.0 1e-06 
0.0 -1.1226 0 -2.0 1e-06 
0.0 -1.1225 0 -2.0 1e-06 
0.0 -1.1224 0 -2.0 1e-06 
0.0 -1.1223 0 -2.0 1e-06 
0.0 -1.1222 0 -2.0 1e-06 
0.0 -1.1221 0 -2.0 1e-06 
0.0 -1.122 0 -2.0 1e-06 
0.0 -1.1219 0 -2.0 1e-06 
0.0 -1.1218 0 -2.0 1e-06 
0.0 -1.1217 0 -2.0 1e-06 
0.0 -1.1216 0 -2.0 1e-06 
0.0 -1.1215 0 -2.0 1e-06 
0.0 -1.1214 0 -2.0 1e-06 
0.0 -1.1213 0 -2.0 1e-06 
0.0 -1.1212 0 -2.0 1e-06 
0.0 -1.1211 0 -2.0 1e-06 
0.0 -1.121 0 -2.0 1e-06 
0.0 -1.1209 0 -2.0 1e-06 
0.0 -1.1208 0 -2.0 1e-06 
0.0 -1.1207 0 -2.0 1e-06 
0.0 -1.1206 0 -2.0 1e-06 
0.0 -1.1205 0 -2.0 1e-06 
0.0 -1.1204 0 -2.0 1e-06 
0.0 -1.1203 0 -2.0 1e-06 
0.0 -1.1202 0 -2.0 1e-06 
0.0 -1.1201 0 -2.0 1e-06 
0.0 -1.12 0 -2.0 1e-06 
0.0 -1.1199 0 -2.0 1e-06 
0.0 -1.1198 0 -2.0 1e-06 
0.0 -1.1197 0 -2.0 1e-06 
0.0 -1.1196 0 -2.0 1e-06 
0.0 -1.1195 0 -2.0 1e-06 
0.0 -1.1194 0 -2.0 1e-06 
0.0 -1.1193 0 -2.0 1e-06 
0.0 -1.1192 0 -2.0 1e-06 
0.0 -1.1191 0 -2.0 1e-06 
0.0 -1.119 0 -2.0 1e-06 
0.0 -1.1189 0 -2.0 1e-06 
0.0 -1.1188 0 -2.0 1e-06 
0.0 -1.1187 0 -2.0 1e-06 
0.0 -1.1186 0 -2.0 1e-06 
0.0 -1.1185 0 -2.0 1e-06 
0.0 -1.1184 0 -2.0 1e-06 
0.0 -1.1183 0 -2.0 1e-06 
0.0 -1.1182 0 -2.0 1e-06 
0.0 -1.1181 0 -2.0 1e-06 
0.0 -1.118 0 -2.0 1e-06 
0.0 -1.1179 0 -2.0 1e-06 
0.0 -1.1178 0 -2.0 1e-06 
0.0 -1.1177 0 -2.0 1e-06 
0.0 -1.1176 0 -2.0 1e-06 
0.0 -1.1175 0 -2.0 1e-06 
0.0 -1.1174 0 -2.0 1e-06 
0.0 -1.1173 0 -2.0 1e-06 
0.0 -1.1172 0 -2.0 1e-06 
0.0 -1.1171 0 -2.0 1e-06 
0.0 -1.117 0 -2.0 1e-06 
0.0 -1.1169 0 -2.0 1e-06 
0.0 -1.1168 0 -2.0 1e-06 
0.0 -1.1167 0 -2.0 1e-06 
0.0 -1.1166 0 -2.0 1e-06 
0.0 -1.1165 0 -2.0 1e-06 
0.0 -1.1164 0 -2.0 1e-06 
0.0 -1.1163 0 -2.0 1e-06 
0.0 -1.1162 0 -2.0 1e-06 
0.0 -1.1161 0 -2.0 1e-06 
0.0 -1.116 0 -2.0 1e-06 
0.0 -1.1159 0 -2.0 1e-06 
0.0 -1.1158 0 -2.0 1e-06 
0.0 -1.1157 0 -2.0 1e-06 
0.0 -1.1156 0 -2.0 1e-06 
0.0 -1.1155 0 -2.0 1e-06 
0.0 -1.1154 0 -2.0 1e-06 
0.0 -1.1153 0 -2.0 1e-06 
0.0 -1.1152 0 -2.0 1e-06 
0.0 -1.1151 0 -2.0 1e-06 
0.0 -1.115 0 -2.0 1e-06 
0.0 -1.1149 0 -2.0 1e-06 
0.0 -1.1148 0 -2.0 1e-06 
0.0 -1.1147 0 -2.0 1e-06 
0.0 -1.1146 0 -2.0 1e-06 
0.0 -1.1145 0 -2.0 1e-06 
0.0 -1.1144 0 -2.0 1e-06 
0.0 -1.1143 0 -2.0 1e-06 
0.0 -1.1142 0 -2.0 1e-06 
0.0 -1.1141 0 -2.0 1e-06 
0.0 -1.114 0 -2.0 1e-06 
0.0 -1.1139 0 -2.0 1e-06 
0.0 -1.1138 0 -2.0 1e-06 
0.0 -1.1137 0 -2.0 1e-06 
0.0 -1.1136 0 -2.0 1e-06 
0.0 -1.1135 0 -2.0 1e-06 
0.0 -1.1134 0 -2.0 1e-06 
0.0 -1.1133 0 -2.0 1e-06 
0.0 -1.1132 0 -2.0 1e-06 
0.0 -1.1131 0 -2.0 1e-06 
0.0 -1.113 0 -2.0 1e-06 
0.0 -1.1129 0 -2.0 1e-06 
0.0 -1.1128 0 -2.0 1e-06 
0.0 -1.1127 0 -2.0 1e-06 
0.0 -1.1126 0 -2.0 1e-06 
0.0 -1.1125 0 -2.0 1e-06 
0.0 -1.1124 0 -2.0 1e-06 
0.0 -1.1123 0 -2.0 1e-06 
0.0 -1.1122 0 -2.0 1e-06 
0.0 -1.1121 0 -2.0 1e-06 
0.0 -1.112 0 -2.0 1e-06 
0.0 -1.1119 0 -2.0 1e-06 
0.0 -1.1118 0 -2.0 1e-06 
0.0 -1.1117 0 -2.0 1e-06 
0.0 -1.1116 0 -2.0 1e-06 
0.0 -1.1115 0 -2.0 1e-06 
0.0 -1.1114 0 -2.0 1e-06 
0.0 -1.1113 0 -2.0 1e-06 
0.0 -1.1112 0 -2.0 1e-06 
0.0 -1.1111 0 -2.0 1e-06 
0.0 -1.111 0 -2.0 1e-06 
0.0 -1.1109 0 -2.0 1e-06 
0.0 -1.1108 0 -2.0 1e-06 
0.0 -1.1107 0 -2.0 1e-06 
0.0 -1.1106 0 -2.0 1e-06 
0.0 -1.1105 0 -2.0 1e-06 
0.0 -1.1104 0 -2.0 1e-06 
0.0 -1.1103 0 -2.0 1e-06 
0.0 -1.1102 0 -2.0 1e-06 
0.0 -1.1101 0 -2.0 1e-06 
0.0 -1.11 0 -2.0 1e-06 
0.0 -1.1099 0 -2.0 1e-06 
0.0 -1.1098 0 -2.0 1e-06 
0.0 -1.1097 0 -2.0 1e-06 
0.0 -1.1096 0 -2.0 1e-06 
0.0 -1.1095 0 -2.0 1e-06 
0.0 -1.1094 0 -2.0 1e-06 
0.0 -1.1093 0 -2.0 1e-06 
0.0 -1.1092 0 -2.0 1e-06 
0.0 -1.1091 0 -2.0 1e-06 
0.0 -1.109 0 -2.0 1e-06 
0.0 -1.1089 0 -2.0 1e-06 
0.0 -1.1088 0 -2.0 1e-06 
0.0 -1.1087 0 -2.0 1e-06 
0.0 -1.1086 0 -2.0 1e-06 
0.0 -1.1085 0 -2.0 1e-06 
0.0 -1.1084 0 -2.0 1e-06 
0.0 -1.1083 0 -2.0 1e-06 
0.0 -1.1082 0 -2.0 1e-06 
0.0 -1.1081 0 -2.0 1e-06 
0.0 -1.108 0 -2.0 1e-06 
0.0 -1.1079 0 -2.0 1e-06 
0.0 -1.1078 0 -2.0 1e-06 
0.0 -1.1077 0 -2.0 1e-06 
0.0 -1.1076 0 -2.0 1e-06 
0.0 -1.1075 0 -2.0 1e-06 
0.0 -1.1074 0 -2.0 1e-06 
0.0 -1.1073 0 -2.0 1e-06 
0.0 -1.1072 0 -2.0 1e-06 
0.0 -1.1071 0 -2.0 1e-06 
0.0 -1.107 0 -2.0 1e-06 
0.0 -1.1069 0 -2.0 1e-06 
0.0 -1.1068 0 -2.0 1e-06 
0.0 -1.1067 0 -2.0 1e-06 
0.0 -1.1066 0 -2.0 1e-06 
0.0 -1.1065 0 -2.0 1e-06 
0.0 -1.1064 0 -2.0 1e-06 
0.0 -1.1063 0 -2.0 1e-06 
0.0 -1.1062 0 -2.0 1e-06 
0.0 -1.1061 0 -2.0 1e-06 
0.0 -1.106 0 -2.0 1e-06 
0.0 -1.1059 0 -2.0 1e-06 
0.0 -1.1058 0 -2.0 1e-06 
0.0 -1.1057 0 -2.0 1e-06 
0.0 -1.1056 0 -2.0 1e-06 
0.0 -1.1055 0 -2.0 1e-06 
0.0 -1.1054 0 -2.0 1e-06 
0.0 -1.1053 0 -2.0 1e-06 
0.0 -1.1052 0 -2.0 1e-06 
0.0 -1.1051 0 -2.0 1e-06 
0.0 -1.105 0 -2.0 1e-06 
0.0 -1.1049 0 -2.0 1e-06 
0.0 -1.1048 0 -2.0 1e-06 
0.0 -1.1047 0 -2.0 1e-06 
0.0 -1.1046 0 -2.0 1e-06 
0.0 -1.1045 0 -2.0 1e-06 
0.0 -1.1044 0 -2.0 1e-06 
0.0 -1.1043 0 -2.0 1e-06 
0.0 -1.1042 0 -2.0 1e-06 
0.0 -1.1041 0 -2.0 1e-06 
0.0 -1.104 0 -2.0 1e-06 
0.0 -1.1039 0 -2.0 1e-06 
0.0 -1.1038 0 -2.0 1e-06 
0.0 -1.1037 0 -2.0 1e-06 
0.0 -1.1036 0 -2.0 1e-06 
0.0 -1.1035 0 -2.0 1e-06 
0.0 -1.1034 0 -2.0 1e-06 
0.0 -1.1033 0 -2.0 1e-06 
0.0 -1.1032 0 -2.0 1e-06 
0.0 -1.1031 0 -2.0 1e-06 
0.0 -1.103 0 -2.0 1e-06 
0.0 -1.1029 0 -2.0 1e-06 
0.0 -1.1028 0 -2.0 1e-06 
0.0 -1.1027 0 -2.0 1e-06 
0.0 -1.1026 0 -2.0 1e-06 
0.0 -1.1025 0 -2.0 1e-06 
0.0 -1.1024 0 -2.0 1e-06 
0.0 -1.1023 0 -2.0 1e-06 
0.0 -1.1022 0 -2.0 1e-06 
0.0 -1.1021 0 -2.0 1e-06 
0.0 -1.102 0 -2.0 1e-06 
0.0 -1.1019 0 -2.0 1e-06 
0.0 -1.1018 0 -2.0 1e-06 
0.0 -1.1017 0 -2.0 1e-06 
0.0 -1.1016 0 -2.0 1e-06 
0.0 -1.1015 0 -2.0 1e-06 
0.0 -1.1014 0 -2.0 1e-06 
0.0 -1.1013 0 -2.0 1e-06 
0.0 -1.1012 0 -2.0 1e-06 
0.0 -1.1011 0 -2.0 1e-06 
0.0 -1.101 0 -2.0 1e-06 
0.0 -1.1009 0 -2.0 1e-06 
0.0 -1.1008 0 -2.0 1e-06 
0.0 -1.1007 0 -2.0 1e-06 
0.0 -1.1006 0 -2.0 1e-06 
0.0 -1.1005 0 -2.0 1e-06 
0.0 -1.1004 0 -2.0 1e-06 
0.0 -1.1003 0 -2.0 1e-06 
0.0 -1.1002 0 -2.0 1e-06 
0.0 -1.1001 0 -2.0 1e-06 
0.0 -1.1 0 -2.0 1e-06 
0.0 -1.0999 0 -2.0 1e-06 
0.0 -1.0998 0 -2.0 1e-06 
0.0 -1.0997 0 -2.0 1e-06 
0.0 -1.0996 0 -2.0 1e-06 
0.0 -1.0995 0 -2.0 1e-06 
0.0 -1.0994 0 -2.0 1e-06 
0.0 -1.0993 0 -2.0 1e-06 
0.0 -1.0992 0 -2.0 1e-06 
0.0 -1.0991 0 -2.0 1e-06 
0.0 -1.099 0 -2.0 1e-06 
0.0 -1.0989 0 -2.0 1e-06 
0.0 -1.0988 0 -2.0 1e-06 
0.0 -1.0987 0 -2.0 1e-06 
0.0 -1.0986 0 -2.0 1e-06 
0.0 -1.0985 0 -2.0 1e-06 
0.0 -1.0984 0 -2.0 1e-06 
0.0 -1.0983 0 -2.0 1e-06 
0.0 -1.0982 0 -2.0 1e-06 
0.0 -1.0981 0 -2.0 1e-06 
0.0 -1.098 0 -2.0 1e-06 
0.0 -1.0979 0 -2.0 1e-06 
0.0 -1.0978 0 -2.0 1e-06 
0.0 -1.0977 0 -2.0 1e-06 
0.0 -1.0976 0 -2.0 1e-06 
0.0 -1.0975 0 -2.0 1e-06 
0.0 -1.0974 0 -2.0 1e-06 
0.0 -1.0973 0 -2.0 1e-06 
0.0 -1.0972 0 -2.0 1e-06 
0.0 -1.0971 0 -2.0 1e-06 
0.0 -1.097 0 -2.0 1e-06 
0.0 -1.0969 0 -2.0 1e-06 
0.0 -1.0968 0 -2.0 1e-06 
0.0 -1.0967 0 -2.0 1e-06 
0.0 -1.0966 0 -2.0 1e-06 
0.0 -1.0965 0 -2.0 1e-06 
0.0 -1.0964 0 -2.0 1e-06 
0.0 -1.0963 0 -2.0 1e-06 
0.0 -1.0962 0 -2.0 1e-06 
0.0 -1.0961 0 -2.0 1e-06 
0.0 -1.096 0 -2.0 1e-06 
0.0 -1.0959 0 -2.0 1e-06 
0.0 -1.0958 0 -2.0 1e-06 
0.0 -1.0957 0 -2.0 1e-06 
0.0 -1.0956 0 -2.0 1e-06 
0.0 -1.0955 0 -2.0 1e-06 
0.0 -1.0954 0 -2.0 1e-06 
0.0 -1.0953 0 -2.0 1e-06 
0.0 -1.0952 0 -2.0 1e-06 
0.0 -1.0951 0 -2.0 1e-06 
0.0 -1.095 0 -2.0 1e-06 
0.0 -1.0949 0 -2.0 1e-06 
0.0 -1.0948 0 -2.0 1e-06 
0.0 -1.0947 0 -2.0 1e-06 
0.0 -1.0946 0 -2.0 1e-06 
0.0 -1.0945 0 -2.0 1e-06 
0.0 -1.0944 0 -2.0 1e-06 
0.0 -1.0943 0 -2.0 1e-06 
0.0 -1.0942 0 -2.0 1e-06 
0.0 -1.0941 0 -2.0 1e-06 
0.0 -1.094 0 -2.0 1e-06 
0.0 -1.0939 0 -2.0 1e-06 
0.0 -1.0938 0 -2.0 1e-06 
0.0 -1.0937 0 -2.0 1e-06 
0.0 -1.0936 0 -2.0 1e-06 
0.0 -1.0935 0 -2.0 1e-06 
0.0 -1.0934 0 -2.0 1e-06 
0.0 -1.0933 0 -2.0 1e-06 
0.0 -1.0932 0 -2.0 1e-06 
0.0 -1.0931 0 -2.0 1e-06 
0.0 -1.093 0 -2.0 1e-06 
0.0 -1.0929 0 -2.0 1e-06 
0.0 -1.0928 0 -2.0 1e-06 
0.0 -1.0927 0 -2.0 1e-06 
0.0 -1.0926 0 -2.0 1e-06 
0.0 -1.0925 0 -2.0 1e-06 
0.0 -1.0924 0 -2.0 1e-06 
0.0 -1.0923 0 -2.0 1e-06 
0.0 -1.0922 0 -2.0 1e-06 
0.0 -1.0921 0 -2.0 1e-06 
0.0 -1.092 0 -2.0 1e-06 
0.0 -1.0919 0 -2.0 1e-06 
0.0 -1.0918 0 -2.0 1e-06 
0.0 -1.0917 0 -2.0 1e-06 
0.0 -1.0916 0 -2.0 1e-06 
0.0 -1.0915 0 -2.0 1e-06 
0.0 -1.0914 0 -2.0 1e-06 
0.0 -1.0913 0 -2.0 1e-06 
0.0 -1.0912 0 -2.0 1e-06 
0.0 -1.0911 0 -2.0 1e-06 
0.0 -1.091 0 -2.0 1e-06 
0.0 -1.0909 0 -2.0 1e-06 
0.0 -1.0908 0 -2.0 1e-06 
0.0 -1.0907 0 -2.0 1e-06 
0.0 -1.0906 0 -2.0 1e-06 
0.0 -1.0905 0 -2.0 1e-06 
0.0 -1.0904 0 -2.0 1e-06 
0.0 -1.0903 0 -2.0 1e-06 
0.0 -1.0902 0 -2.0 1e-06 
0.0 -1.0901 0 -2.0 1e-06 
0.0 -1.09 0 -2.0 1e-06 
0.0 -1.0899 0 -2.0 1e-06 
0.0 -1.0898 0 -2.0 1e-06 
0.0 -1.0897 0 -2.0 1e-06 
0.0 -1.0896 0 -2.0 1e-06 
0.0 -1.0895 0 -2.0 1e-06 
0.0 -1.0894 0 -2.0 1e-06 
0.0 -1.0893 0 -2.0 1e-06 
0.0 -1.0892 0 -2.0 1e-06 
0.0 -1.0891 0 -2.0 1e-06 
0.0 -1.089 0 -2.0 1e-06 
0.0 -1.0889 0 -2.0 1e-06 
0.0 -1.0888 0 -2.0 1e-06 
0.0 -1.0887 0 -2.0 1e-06 
0.0 -1.0886 0 -2.0 1e-06 
0.0 -1.0885 0 -2.0 1e-06 
0.0 -1.0884 0 -2.0 1e-06 
0.0 -1.0883 0 -2.0 1e-06 
0.0 -1.0882 0 -2.0 1e-06 
0.0 -1.0881 0 -2.0 1e-06 
0.0 -1.088 0 -2.0 1e-06 
0.0 -1.0879 0 -2.0 1e-06 
0.0 -1.0878 0 -2.0 1e-06 
0.0 -1.0877 0 -2.0 1e-06 
0.0 -1.0876 0 -2.0 1e-06 
0.0 -1.0875 0 -2.0 1e-06 
0.0 -1.0874 0 -2.0 1e-06 
0.0 -1.0873 0 -2.0 1e-06 
0.0 -1.0872 0 -2.0 1e-06 
0.0 -1.0871 0 -2.0 1e-06 
0.0 -1.087 0 -2.0 1e-06 
0.0 -1.0869 0 -2.0 1e-06 
0.0 -1.0868 0 -2.0 1e-06 
0.0 -1.0867 0 -2.0 1e-06 
0.0 -1.0866 0 -2.0 1e-06 
0.0 -1.0865 0 -2.0 1e-06 
0.0 -1.0864 0 -2.0 1e-06 
0.0 -1.0863 0 -2.0 1e-06 
0.0 -1.0862 0 -2.0 1e-06 
0.0 -1.0861 0 -2.0 1e-06 
0.0 -1.086 0 -2.0 1e-06 
0.0 -1.0859 0 -2.0 1e-06 
0.0 -1.0858 0 -2.0 1e-06 
0.0 -1.0857 0 -2.0 1e-06 
0.0 -1.0856 0 -2.0 1e-06 
0.0 -1.0855 0 -2.0 1e-06 
0.0 -1.0854 0 -2.0 1e-06 
0.0 -1.0853 0 -2.0 1e-06 
0.0 -1.0852 0 -2.0 1e-06 
0.0 -1.0851 0 -2.0 1e-06 
0.0 -1.085 0 -2.0 1e-06 
0.0 -1.0849 0 -2.0 1e-06 
0.0 -1.0848 0 -2.0 1e-06 
0.0 -1.0847 0 -2.0 1e-06 
0.0 -1.0846 0 -2.0 1e-06 
0.0 -1.0845 0 -2.0 1e-06 
0.0 -1.0844 0 -2.0 1e-06 
0.0 -1.0843 0 -2.0 1e-06 
0.0 -1.0842 0 -2.0 1e-06 
0.0 -1.0841 0 -2.0 1e-06 
0.0 -1.084 0 -2.0 1e-06 
0.0 -1.0839 0 -2.0 1e-06 
0.0 -1.0838 0 -2.0 1e-06 
0.0 -1.0837 0 -2.0 1e-06 
0.0 -1.0836 0 -2.0 1e-06 
0.0 -1.0835 0 -2.0 1e-06 
0.0 -1.0834 0 -2.0 1e-06 
0.0 -1.0833 0 -2.0 1e-06 
0.0 -1.0832 0 -2.0 1e-06 
0.0 -1.0831 0 -2.0 1e-06 
0.0 -1.083 0 -2.0 1e-06 
0.0 -1.0829 0 -2.0 1e-06 
0.0 -1.0828 0 -2.0 1e-06 
0.0 -1.0827 0 -2.0 1e-06 
0.0 -1.0826 0 -2.0 1e-06 
0.0 -1.0825 0 -2.0 1e-06 
0.0 -1.0824 0 -2.0 1e-06 
0.0 -1.0823 0 -2.0 1e-06 
0.0 -1.0822 0 -2.0 1e-06 
0.0 -1.0821 0 -2.0 1e-06 
0.0 -1.082 0 -2.0 1e-06 
0.0 -1.0819 0 -2.0 1e-06 
0.0 -1.0818 0 -2.0 1e-06 
0.0 -1.0817 0 -2.0 1e-06 
0.0 -1.0816 0 -2.0 1e-06 
0.0 -1.0815 0 -2.0 1e-06 
0.0 -1.0814 0 -2.0 1e-06 
0.0 -1.0813 0 -2.0 1e-06 
0.0 -1.0812 0 -2.0 1e-06 
0.0 -1.0811 0 -2.0 1e-06 
0.0 -1.081 0 -2.0 1e-06 
0.0 -1.0809 0 -2.0 1e-06 
0.0 -1.0808 0 -2.0 1e-06 
0.0 -1.0807 0 -2.0 1e-06 
0.0 -1.0806 0 -2.0 1e-06 
0.0 -1.0805 0 -2.0 1e-06 
0.0 -1.0804 0 -2.0 1e-06 
0.0 -1.0803 0 -2.0 1e-06 
0.0 -1.0802 0 -2.0 1e-06 
0.0 -1.0801 0 -2.0 1e-06 
0.0 -1.08 0 -2.0 1e-06 
0.0 -1.0799 0 -2.0 1e-06 
0.0 -1.0798 0 -2.0 1e-06 
0.0 -1.0797 0 -2.0 1e-06 
0.0 -1.0796 0 -2.0 1e-06 
0.0 -1.0795 0 -2.0 1e-06 
0.0 -1.0794 0 -2.0 1e-06 
0.0 -1.0793 0 -2.0 1e-06 
0.0 -1.0792 0 -2.0 1e-06 
0.0 -1.0791 0 -2.0 1e-06 
0.0 -1.079 0 -2.0 1e-06 
0.0 -1.0789 0 -2.0 1e-06 
0.0 -1.0788 0 -2.0 1e-06 
0.0 -1.0787 0 -2.0 1e-06 
0.0 -1.0786 0 -2.0 1e-06 
0.0 -1.0785 0 -2.0 1e-06 
0.0 -1.0784 0 -2.0 1e-06 
0.0 -1.0783 0 -2.0 1e-06 
0.0 -1.0782 0 -2.0 1e-06 
0.0 -1.0781 0 -2.0 1e-06 
0.0 -1.078 0 -2.0 1e-06 
0.0 -1.0779 0 -2.0 1e-06 
0.0 -1.0778 0 -2.0 1e-06 
0.0 -1.0777 0 -2.0 1e-06 
0.0 -1.0776 0 -2.0 1e-06 
0.0 -1.0775 0 -2.0 1e-06 
0.0 -1.0774 0 -2.0 1e-06 
0.0 -1.0773 0 -2.0 1e-06 
0.0 -1.0772 0 -2.0 1e-06 
0.0 -1.0771 0 -2.0 1e-06 
0.0 -1.077 0 -2.0 1e-06 
0.0 -1.0769 0 -2.0 1e-06 
0.0 -1.0768 0 -2.0 1e-06 
0.0 -1.0767 0 -2.0 1e-06 
0.0 -1.0766 0 -2.0 1e-06 
0.0 -1.0765 0 -2.0 1e-06 
0.0 -1.0764 0 -2.0 1e-06 
0.0 -1.0763 0 -2.0 1e-06 
0.0 -1.0762 0 -2.0 1e-06 
0.0 -1.0761 0 -2.0 1e-06 
0.0 -1.076 0 -2.0 1e-06 
0.0 -1.0759 0 -2.0 1e-06 
0.0 -1.0758 0 -2.0 1e-06 
0.0 -1.0757 0 -2.0 1e-06 
0.0 -1.0756 0 -2.0 1e-06 
0.0 -1.0755 0 -2.0 1e-06 
0.0 -1.0754 0 -2.0 1e-06 
0.0 -1.0753 0 -2.0 1e-06 
0.0 -1.0752 0 -2.0 1e-06 
0.0 -1.0751 0 -2.0 1e-06 
0.0 -1.075 0 -2.0 1e-06 
0.0 -1.0749 0 -2.0 1e-06 
0.0 -1.0748 0 -2.0 1e-06 
0.0 -1.0747 0 -2.0 1e-06 
0.0 -1.0746 0 -2.0 1e-06 
0.0 -1.0745 0 -2.0 1e-06 
0.0 -1.0744 0 -2.0 1e-06 
0.0 -1.0743 0 -2.0 1e-06 
0.0 -1.0742 0 -2.0 1e-06 
0.0 -1.0741 0 -2.0 1e-06 
0.0 -1.074 0 -2.0 1e-06 
0.0 -1.0739 0 -2.0 1e-06 
0.0 -1.0738 0 -2.0 1e-06 
0.0 -1.0737 0 -2.0 1e-06 
0.0 -1.0736 0 -2.0 1e-06 
0.0 -1.0735 0 -2.0 1e-06 
0.0 -1.0734 0 -2.0 1e-06 
0.0 -1.0733 0 -2.0 1e-06 
0.0 -1.0732 0 -2.0 1e-06 
0.0 -1.0731 0 -2.0 1e-06 
0.0 -1.073 0 -2.0 1e-06 
0.0 -1.0729 0 -2.0 1e-06 
0.0 -1.0728 0 -2.0 1e-06 
0.0 -1.0727 0 -2.0 1e-06 
0.0 -1.0726 0 -2.0 1e-06 
0.0 -1.0725 0 -2.0 1e-06 
0.0 -1.0724 0 -2.0 1e-06 
0.0 -1.0723 0 -2.0 1e-06 
0.0 -1.0722 0 -2.0 1e-06 
0.0 -1.0721 0 -2.0 1e-06 
0.0 -1.072 0 -2.0 1e-06 
0.0 -1.0719 0 -2.0 1e-06 
0.0 -1.0718 0 -2.0 1e-06 
0.0 -1.0717 0 -2.0 1e-06 
0.0 -1.0716 0 -2.0 1e-06 
0.0 -1.0715 0 -2.0 1e-06 
0.0 -1.0714 0 -2.0 1e-06 
0.0 -1.0713 0 -2.0 1e-06 
0.0 -1.0712 0 -2.0 1e-06 
0.0 -1.0711 0 -2.0 1e-06 
0.0 -1.071 0 -2.0 1e-06 
0.0 -1.0709 0 -2.0 1e-06 
0.0 -1.0708 0 -2.0 1e-06 
0.0 -1.0707 0 -2.0 1e-06 
0.0 -1.0706 0 -2.0 1e-06 
0.0 -1.0705 0 -2.0 1e-06 
0.0 -1.0704 0 -2.0 1e-06 
0.0 -1.0703 0 -2.0 1e-06 
0.0 -1.0702 0 -2.0 1e-06 
0.0 -1.0701 0 -2.0 1e-06 
0.0 -1.07 0 -2.0 1e-06 
0.0 -1.0699 0 -2.0 1e-06 
0.0 -1.0698 0 -2.0 1e-06 
0.0 -1.0697 0 -2.0 1e-06 
0.0 -1.0696 0 -2.0 1e-06 
0.0 -1.0695 0 -2.0 1e-06 
0.0 -1.0694 0 -2.0 1e-06 
0.0 -1.0693 0 -2.0 1e-06 
0.0 -1.0692 0 -2.0 1e-06 
0.0 -1.0691 0 -2.0 1e-06 
0.0 -1.069 0 -2.0 1e-06 
0.0 -1.0689 0 -2.0 1e-06 
0.0 -1.0688 0 -2.0 1e-06 
0.0 -1.0687 0 -2.0 1e-06 
0.0 -1.0686 0 -2.0 1e-06 
0.0 -1.0685 0 -2.0 1e-06 
0.0 -1.0684 0 -2.0 1e-06 
0.0 -1.0683 0 -2.0 1e-06 
0.0 -1.0682 0 -2.0 1e-06 
0.0 -1.0681 0 -2.0 1e-06 
0.0 -1.068 0 -2.0 1e-06 
0.0 -1.0679 0 -2.0 1e-06 
0.0 -1.0678 0 -2.0 1e-06 
0.0 -1.0677 0 -2.0 1e-06 
0.0 -1.0676 0 -2.0 1e-06 
0.0 -1.0675 0 -2.0 1e-06 
0.0 -1.0674 0 -2.0 1e-06 
0.0 -1.0673 0 -2.0 1e-06 
0.0 -1.0672 0 -2.0 1e-06 
0.0 -1.0671 0 -2.0 1e-06 
0.0 -1.067 0 -2.0 1e-06 
0.0 -1.0669 0 -2.0 1e-06 
0.0 -1.0668 0 -2.0 1e-06 
0.0 -1.0667 0 -2.0 1e-06 
0.0 -1.0666 0 -2.0 1e-06 
0.0 -1.0665 0 -2.0 1e-06 
0.0 -1.0664 0 -2.0 1e-06 
0.0 -1.0663 0 -2.0 1e-06 
0.0 -1.0662 0 -2.0 1e-06 
0.0 -1.0661 0 -2.0 1e-06 
0.0 -1.066 0 -2.0 1e-06 
0.0 -1.0659 0 -2.0 1e-06 
0.0 -1.0658 0 -2.0 1e-06 
0.0 -1.0657 0 -2.0 1e-06 
0.0 -1.0656 0 -2.0 1e-06 
0.0 -1.0655 0 -2.0 1e-06 
0.0 -1.0654 0 -2.0 1e-06 
0.0 -1.0653 0 -2.0 1e-06 
0.0 -1.0652 0 -2.0 1e-06 
0.0 -1.0651 0 -2.0 1e-06 
0.0 -1.065 0 -2.0 1e-06 
0.0 -1.0649 0 -2.0 1e-06 
0.0 -1.0648 0 -2.0 1e-06 
0.0 -1.0647 0 -2.0 1e-06 
0.0 -1.0646 0 -2.0 1e-06 
0.0 -1.0645 0 -2.0 1e-06 
0.0 -1.0644 0 -2.0 1e-06 
0.0 -1.0643 0 -2.0 1e-06 
0.0 -1.0642 0 -2.0 1e-06 
0.0 -1.0641 0 -2.0 1e-06 
0.0 -1.064 0 -2.0 1e-06 
0.0 -1.0639 0 -2.0 1e-06 
0.0 -1.0638 0 -2.0 1e-06 
0.0 -1.0637 0 -2.0 1e-06 
0.0 -1.0636 0 -2.0 1e-06 
0.0 -1.0635 0 -2.0 1e-06 
0.0 -1.0634 0 -2.0 1e-06 
0.0 -1.0633 0 -2.0 1e-06 
0.0 -1.0632 0 -2.0 1e-06 
0.0 -1.0631 0 -2.0 1e-06 
0.0 -1.063 0 -2.0 1e-06 
0.0 -1.0629 0 -2.0 1e-06 
0.0 -1.0628 0 -2.0 1e-06 
0.0 -1.0627 0 -2.0 1e-06 
0.0 -1.0626 0 -2.0 1e-06 
0.0 -1.0625 0 -2.0 1e-06 
0.0 -1.0624 0 -2.0 1e-06 
0.0 -1.0623 0 -2.0 1e-06 
0.0 -1.0622 0 -2.0 1e-06 
0.0 -1.0621 0 -2.0 1e-06 
0.0 -1.062 0 -2.0 1e-06 
0.0 -1.0619 0 -2.0 1e-06 
0.0 -1.0618 0 -2.0 1e-06 
0.0 -1.0617 0 -2.0 1e-06 
0.0 -1.0616 0 -2.0 1e-06 
0.0 -1.0615 0 -2.0 1e-06 
0.0 -1.0614 0 -2.0 1e-06 
0.0 -1.0613 0 -2.0 1e-06 
0.0 -1.0612 0 -2.0 1e-06 
0.0 -1.0611 0 -2.0 1e-06 
0.0 -1.061 0 -2.0 1e-06 
0.0 -1.0609 0 -2.0 1e-06 
0.0 -1.0608 0 -2.0 1e-06 
0.0 -1.0607 0 -2.0 1e-06 
0.0 -1.0606 0 -2.0 1e-06 
0.0 -1.0605 0 -2.0 1e-06 
0.0 -1.0604 0 -2.0 1e-06 
0.0 -1.0603 0 -2.0 1e-06 
0.0 -1.0602 0 -2.0 1e-06 
0.0 -1.0601 0 -2.0 1e-06 
0.0 -1.06 0 -2.0 1e-06 
0.0 -1.0599 0 -2.0 1e-06 
0.0 -1.0598 0 -2.0 1e-06 
0.0 -1.0597 0 -2.0 1e-06 
0.0 -1.0596 0 -2.0 1e-06 
0.0 -1.0595 0 -2.0 1e-06 
0.0 -1.0594 0 -2.0 1e-06 
0.0 -1.0593 0 -2.0 1e-06 
0.0 -1.0592 0 -2.0 1e-06 
0.0 -1.0591 0 -2.0 1e-06 
0.0 -1.059 0 -2.0 1e-06 
0.0 -1.0589 0 -2.0 1e-06 
0.0 -1.0588 0 -2.0 1e-06 
0.0 -1.0587 0 -2.0 1e-06 
0.0 -1.0586 0 -2.0 1e-06 
0.0 -1.0585 0 -2.0 1e-06 
0.0 -1.0584 0 -2.0 1e-06 
0.0 -1.0583 0 -2.0 1e-06 
0.0 -1.0582 0 -2.0 1e-06 
0.0 -1.0581 0 -2.0 1e-06 
0.0 -1.058 0 -2.0 1e-06 
0.0 -1.0579 0 -2.0 1e-06 
0.0 -1.0578 0 -2.0 1e-06 
0.0 -1.0577 0 -2.0 1e-06 
0.0 -1.0576 0 -2.0 1e-06 
0.0 -1.0575 0 -2.0 1e-06 
0.0 -1.0574 0 -2.0 1e-06 
0.0 -1.0573 0 -2.0 1e-06 
0.0 -1.0572 0 -2.0 1e-06 
0.0 -1.0571 0 -2.0 1e-06 
0.0 -1.057 0 -2.0 1e-06 
0.0 -1.0569 0 -2.0 1e-06 
0.0 -1.0568 0 -2.0 1e-06 
0.0 -1.0567 0 -2.0 1e-06 
0.0 -1.0566 0 -2.0 1e-06 
0.0 -1.0565 0 -2.0 1e-06 
0.0 -1.0564 0 -2.0 1e-06 
0.0 -1.0563 0 -2.0 1e-06 
0.0 -1.0562 0 -2.0 1e-06 
0.0 -1.0561 0 -2.0 1e-06 
0.0 -1.056 0 -2.0 1e-06 
0.0 -1.0559 0 -2.0 1e-06 
0.0 -1.0558 0 -2.0 1e-06 
0.0 -1.0557 0 -2.0 1e-06 
0.0 -1.0556 0 -2.0 1e-06 
0.0 -1.0555 0 -2.0 1e-06 
0.0 -1.0554 0 -2.0 1e-06 
0.0 -1.0553 0 -2.0 1e-06 
0.0 -1.0552 0 -2.0 1e-06 
0.0 -1.0551 0 -2.0 1e-06 
0.0 -1.055 0 -2.0 1e-06 
0.0 -1.0549 0 -2.0 1e-06 
0.0 -1.0548 0 -2.0 1e-06 
0.0 -1.0547 0 -2.0 1e-06 
0.0 -1.0546 0 -2.0 1e-06 
0.0 -1.0545 0 -2.0 1e-06 
0.0 -1.0544 0 -2.0 1e-06 
0.0 -1.0543 0 -2.0 1e-06 
0.0 -1.0542 0 -2.0 1e-06 
0.0 -1.0541 0 -2.0 1e-06 
0.0 -1.054 0 -2.0 1e-06 
0.0 -1.0539 0 -2.0 1e-06 
0.0 -1.0538 0 -2.0 1e-06 
0.0 -1.0537 0 -2.0 1e-06 
0.0 -1.0536 0 -2.0 1e-06 
0.0 -1.0535 0 -2.0 1e-06 
0.0 -1.0534 0 -2.0 1e-06 
0.0 -1.0533 0 -2.0 1e-06 
0.0 -1.0532 0 -2.0 1e-06 
0.0 -1.0531 0 -2.0 1e-06 
0.0 -1.053 0 -2.0 1e-06 
0.0 -1.0529 0 -2.0 1e-06 
0.0 -1.0528 0 -2.0 1e-06 
0.0 -1.0527 0 -2.0 1e-06 
0.0 -1.0526 0 -2.0 1e-06 
0.0 -1.0525 0 -2.0 1e-06 
0.0 -1.0524 0 -2.0 1e-06 
0.0 -1.0523 0 -2.0 1e-06 
0.0 -1.0522 0 -2.0 1e-06 
0.0 -1.0521 0 -2.0 1e-06 
0.0 -1.052 0 -2.0 1e-06 
0.0 -1.0519 0 -2.0 1e-06 
0.0 -1.0518 0 -2.0 1e-06 
0.0 -1.0517 0 -2.0 1e-06 
0.0 -1.0516 0 -2.0 1e-06 
0.0 -1.0515 0 -2.0 1e-06 
0.0 -1.0514 0 -2.0 1e-06 
0.0 -1.0513 0 -2.0 1e-06 
0.0 -1.0512 0 -2.0 1e-06 
0.0 -1.0511 0 -2.0 1e-06 
0.0 -1.051 0 -2.0 1e-06 
0.0 -1.0509 0 -2.0 1e-06 
0.0 -1.0508 0 -2.0 1e-06 
0.0 -1.0507 0 -2.0 1e-06 
0.0 -1.0506 0 -2.0 1e-06 
0.0 -1.0505 0 -2.0 1e-06 
0.0 -1.0504 0 -2.0 1e-06 
0.0 -1.0503 0 -2.0 1e-06 
0.0 -1.0502 0 -2.0 1e-06 
0.0 -1.0501 0 -2.0 1e-06 
0.0 -1.05 0 -2.0 1e-06 
0.0 -1.0499 0 -2.0 1e-06 
0.0 -1.0498 0 -2.0 1e-06 
0.0 -1.0497 0 -2.0 1e-06 
0.0 -1.0496 0 -2.0 1e-06 
0.0 -1.0495 0 -2.0 1e-06 
0.0 -1.0494 0 -2.0 1e-06 
0.0 -1.0493 0 -2.0 1e-06 
0.0 -1.0492 0 -2.0 1e-06 
0.0 -1.0491 0 -2.0 1e-06 
0.0 -1.049 0 -2.0 1e-06 
0.0 -1.0489 0 -2.0 1e-06 
0.0 -1.0488 0 -2.0 1e-06 
0.0 -1.0487 0 -2.0 1e-06 
0.0 -1.0486 0 -2.0 1e-06 
0.0 -1.0485 0 -2.0 1e-06 
0.0 -1.0484 0 -2.0 1e-06 
0.0 -1.0483 0 -2.0 1e-06 
0.0 -1.0482 0 -2.0 1e-06 
0.0 -1.0481 0 -2.0 1e-06 
0.0 -1.048 0 -2.0 1e-06 
0.0 -1.0479 0 -2.0 1e-06 
0.0 -1.0478 0 -2.0 1e-06 
0.0 -1.0477 0 -2.0 1e-06 
0.0 -1.0476 0 -2.0 1e-06 
0.0 -1.0475 0 -2.0 1e-06 
0.0 -1.0474 0 -2.0 1e-06 
0.0 -1.0473 0 -2.0 1e-06 
0.0 -1.0472 0 -2.0 1e-06 
0.0 -1.0471 0 -2.0 1e-06 
0.0 -1.047 0 -2.0 1e-06 
0.0 -1.0469 0 -2.0 1e-06 
0.0 -1.0468 0 -2.0 1e-06 
0.0 -1.0467 0 -2.0 1e-06 
0.0 -1.0466 0 -2.0 1e-06 
0.0 -1.0465 0 -2.0 1e-06 
0.0 -1.0464 0 -2.0 1e-06 
0.0 -1.0463 0 -2.0 1e-06 
0.0 -1.0462 0 -2.0 1e-06 
0.0 -1.0461 0 -2.0 1e-06 
0.0 -1.046 0 -2.0 1e-06 
0.0 -1.0459 0 -2.0 1e-06 
0.0 -1.0458 0 -2.0 1e-06 
0.0 -1.0457 0 -2.0 1e-06 
0.0 -1.0456 0 -2.0 1e-06 
0.0 -1.0455 0 -2.0 1e-06 
0.0 -1.0454 0 -2.0 1e-06 
0.0 -1.0453 0 -2.0 1e-06 
0.0 -1.0452 0 -2.0 1e-06 
0.0 -1.0451 0 -2.0 1e-06 
0.0 -1.045 0 -2.0 1e-06 
0.0 -1.0449 0 -2.0 1e-06 
0.0 -1.0448 0 -2.0 1e-06 
0.0 -1.0447 0 -2.0 1e-06 
0.0 -1.0446 0 -2.0 1e-06 
0.0 -1.0445 0 -2.0 1e-06 
0.0 -1.0444 0 -2.0 1e-06 
0.0 -1.0443 0 -2.0 1e-06 
0.0 -1.0442 0 -2.0 1e-06 
0.0 -1.0441 0 -2.0 1e-06 
0.0 -1.044 0 -2.0 1e-06 
0.0 -1.0439 0 -2.0 1e-06 
0.0 -1.0438 0 -2.0 1e-06 
0.0 -1.0437 0 -2.0 1e-06 
0.0 -1.0436 0 -2.0 1e-06 
0.0 -1.0435 0 -2.0 1e-06 
0.0 -1.0434 0 -2.0 1e-06 
0.0 -1.0433 0 -2.0 1e-06 
0.0 -1.0432 0 -2.0 1e-06 
0.0 -1.0431 0 -2.0 1e-06 
0.0 -1.043 0 -2.0 1e-06 
0.0 -1.0429 0 -2.0 1e-06 
0.0 -1.0428 0 -2.0 1e-06 
0.0 -1.0427 0 -2.0 1e-06 
0.0 -1.0426 0 -2.0 1e-06 
0.0 -1.0425 0 -2.0 1e-06 
0.0 -1.0424 0 -2.0 1e-06 
0.0 -1.0423 0 -2.0 1e-06 
0.0 -1.0422 0 -2.0 1e-06 
0.0 -1.0421 0 -2.0 1e-06 
0.0 -1.042 0 -2.0 1e-06 
0.0 -1.0419 0 -2.0 1e-06 
0.0 -1.0418 0 -2.0 1e-06 
0.0 -1.0417 0 -2.0 1e-06 
0.0 -1.0416 0 -2.0 1e-06 
0.0 -1.0415 0 -2.0 1e-06 
0.0 -1.0414 0 -2.0 1e-06 
0.0 -1.0413 0 -2.0 1e-06 
0.0 -1.0412 0 -2.0 1e-06 
0.0 -1.0411 0 -2.0 1e-06 
0.0 -1.041 0 -2.0 1e-06 
0.0 -1.0409 0 -2.0 1e-06 
0.0 -1.0408 0 -2.0 1e-06 
0.0 -1.0407 0 -2.0 1e-06 
0.0 -1.0406 0 -2.0 1e-06 
0.0 -1.0405 0 -2.0 1e-06 
0.0 -1.0404 0 -2.0 1e-06 
0.0 -1.0403 0 -2.0 1e-06 
0.0 -1.0402 0 -2.0 1e-06 
0.0 -1.0401 0 -2.0 1e-06 
0.0 -1.04 0 -2.0 1e-06 
0.0 -1.0399 0 -2.0 1e-06 
0.0 -1.0398 0 -2.0 1e-06 
0.0 -1.0397 0 -2.0 1e-06 
0.0 -1.0396 0 -2.0 1e-06 
0.0 -1.0395 0 -2.0 1e-06 
0.0 -1.0394 0 -2.0 1e-06 
0.0 -1.0393 0 -2.0 1e-06 
0.0 -1.0392 0 -2.0 1e-06 
0.0 -1.0391 0 -2.0 1e-06 
0.0 -1.039 0 -2.0 1e-06 
0.0 -1.0389 0 -2.0 1e-06 
0.0 -1.0388 0 -2.0 1e-06 
0.0 -1.0387 0 -2.0 1e-06 
0.0 -1.0386 0 -2.0 1e-06 
0.0 -1.0385 0 -2.0 1e-06 
0.0 -1.0384 0 -2.0 1e-06 
0.0 -1.0383 0 -2.0 1e-06 
0.0 -1.0382 0 -2.0 1e-06 
0.0 -1.0381 0 -2.0 1e-06 
0.0 -1.038 0 -2.0 1e-06 
0.0 -1.0379 0 -2.0 1e-06 
0.0 -1.0378 0 -2.0 1e-06 
0.0 -1.0377 0 -2.0 1e-06 
0.0 -1.0376 0 -2.0 1e-06 
0.0 -1.0375 0 -2.0 1e-06 
0.0 -1.0374 0 -2.0 1e-06 
0.0 -1.0373 0 -2.0 1e-06 
0.0 -1.0372 0 -2.0 1e-06 
0.0 -1.0371 0 -2.0 1e-06 
0.0 -1.037 0 -2.0 1e-06 
0.0 -1.0369 0 -2.0 1e-06 
0.0 -1.0368 0 -2.0 1e-06 
0.0 -1.0367 0 -2.0 1e-06 
0.0 -1.0366 0 -2.0 1e-06 
0.0 -1.0365 0 -2.0 1e-06 
0.0 -1.0364 0 -2.0 1e-06 
0.0 -1.0363 0 -2.0 1e-06 
0.0 -1.0362 0 -2.0 1e-06 
0.0 -1.0361 0 -2.0 1e-06 
0.0 -1.036 0 -2.0 1e-06 
0.0 -1.0359 0 -2.0 1e-06 
0.0 -1.0358 0 -2.0 1e-06 
0.0 -1.0357 0 -2.0 1e-06 
0.0 -1.0356 0 -2.0 1e-06 
0.0 -1.0355 0 -2.0 1e-06 
0.0 -1.0354 0 -2.0 1e-06 
0.0 -1.0353 0 -2.0 1e-06 
0.0 -1.0352 0 -2.0 1e-06 
0.0 -1.0351 0 -2.0 1e-06 
0.0 -1.035 0 -2.0 1e-06 
0.0 -1.0349 0 -2.0 1e-06 
0.0 -1.0348 0 -2.0 1e-06 
0.0 -1.0347 0 -2.0 1e-06 
0.0 -1.0346 0 -2.0 1e-06 
0.0 -1.0345 0 -2.0 1e-06 
0.0 -1.0344 0 -2.0 1e-06 
0.0 -1.0343 0 -2.0 1e-06 
0.0 -1.0342 0 -2.0 1e-06 
0.0 -1.0341 0 -2.0 1e-06 
0.0 -1.034 0 -2.0 1e-06 
0.0 -1.0339 0 -2.0 1e-06 
0.0 -1.0338 0 -2.0 1e-06 
0.0 -1.0337 0 -2.0 1e-06 
0.0 -1.0336 0 -2.0 1e-06 
0.0 -1.0335 0 -2.0 1e-06 
0.0 -1.0334 0 -2.0 1e-06 
0.0 -1.0333 0 -2.0 1e-06 
0.0 -1.0332 0 -2.0 1e-06 
0.0 -1.0331 0 -2.0 1e-06 
0.0 -1.033 0 -2.0 1e-06 
0.0 -1.0329 0 -2.0 1e-06 
0.0 -1.0328 0 -2.0 1e-06 
0.0 -1.0327 0 -2.0 1e-06 
0.0 -1.0326 0 -2.0 1e-06 
0.0 -1.0325 0 -2.0 1e-06 
0.0 -1.0324 0 -2.0 1e-06 
0.0 -1.0323 0 -2.0 1e-06 
0.0 -1.0322 0 -2.0 1e-06 
0.0 -1.0321 0 -2.0 1e-06 
0.0 -1.032 0 -2.0 1e-06 
0.0 -1.0319 0 -2.0 1e-06 
0.0 -1.0318 0 -2.0 1e-06 
0.0 -1.0317 0 -2.0 1e-06 
0.0 -1.0316 0 -2.0 1e-06 
0.0 -1.0315 0 -2.0 1e-06 
0.0 -1.0314 0 -2.0 1e-06 
0.0 -1.0313 0 -2.0 1e-06 
0.0 -1.0312 0 -2.0 1e-06 
0.0 -1.0311 0 -2.0 1e-06 
0.0 -1.031 0 -2.0 1e-06 
0.0 -1.0309 0 -2.0 1e-06 
0.0 -1.0308 0 -2.0 1e-06 
0.0 -1.0307 0 -2.0 1e-06 
0.0 -1.0306 0 -2.0 1e-06 
0.0 -1.0305 0 -2.0 1e-06 
0.0 -1.0304 0 -2.0 1e-06 
0.0 -1.0303 0 -2.0 1e-06 
0.0 -1.0302 0 -2.0 1e-06 
0.0 -1.0301 0 -2.0 1e-06 
0.0 -1.03 0 -2.0 1e-06 
0.0 -1.0299 0 -2.0 1e-06 
0.0 -1.0298 0 -2.0 1e-06 
0.0 -1.0297 0 -2.0 1e-06 
0.0 -1.0296 0 -2.0 1e-06 
0.0 -1.0295 0 -2.0 1e-06 
0.0 -1.0294 0 -2.0 1e-06 
0.0 -1.0293 0 -2.0 1e-06 
0.0 -1.0292 0 -2.0 1e-06 
0.0 -1.0291 0 -2.0 1e-06 
0.0 -1.029 0 -2.0 1e-06 
0.0 -1.0289 0 -2.0 1e-06 
0.0 -1.0288 0 -2.0 1e-06 
0.0 -1.0287 0 -2.0 1e-06 
0.0 -1.0286 0 -2.0 1e-06 
0.0 -1.0285 0 -2.0 1e-06 
0.0 -1.0284 0 -2.0 1e-06 
0.0 -1.0283 0 -2.0 1e-06 
0.0 -1.0282 0 -2.0 1e-06 
0.0 -1.0281 0 -2.0 1e-06 
0.0 -1.028 0 -2.0 1e-06 
0.0 -1.0279 0 -2.0 1e-06 
0.0 -1.0278 0 -2.0 1e-06 
0.0 -1.0277 0 -2.0 1e-06 
0.0 -1.0276 0 -2.0 1e-06 
0.0 -1.0275 0 -2.0 1e-06 
0.0 -1.0274 0 -2.0 1e-06 
0.0 -1.0273 0 -2.0 1e-06 
0.0 -1.0272 0 -2.0 1e-06 
0.0 -1.0271 0 -2.0 1e-06 
0.0 -1.027 0 -2.0 1e-06 
0.0 -1.0269 0 -2.0 1e-06 
0.0 -1.0268 0 -2.0 1e-06 
0.0 -1.0267 0 -2.0 1e-06 
0.0 -1.0266 0 -2.0 1e-06 
0.0 -1.0265 0 -2.0 1e-06 
0.0 -1.0264 0 -2.0 1e-06 
0.0 -1.0263 0 -2.0 1e-06 
0.0 -1.0262 0 -2.0 1e-06 
0.0 -1.0261 0 -2.0 1e-06 
0.0 -1.026 0 -2.0 1e-06 
0.0 -1.0259 0 -2.0 1e-06 
0.0 -1.0258 0 -2.0 1e-06 
0.0 -1.0257 0 -2.0 1e-06 
0.0 -1.0256 0 -2.0 1e-06 
0.0 -1.0255 0 -2.0 1e-06 
0.0 -1.0254 0 -2.0 1e-06 
0.0 -1.0253 0 -2.0 1e-06 
0.0 -1.0252 0 -2.0 1e-06 
0.0 -1.0251 0 -2.0 1e-06 
0.0 -1.025 0 -2.0 1e-06 
0.0 -1.0249 0 -2.0 1e-06 
0.0 -1.0248 0 -2.0 1e-06 
0.0 -1.0247 0 -2.0 1e-06 
0.0 -1.0246 0 -2.0 1e-06 
0.0 -1.0245 0 -2.0 1e-06 
0.0 -1.0244 0 -2.0 1e-06 
0.0 -1.0243 0 -2.0 1e-06 
0.0 -1.0242 0 -2.0 1e-06 
0.0 -1.0241 0 -2.0 1e-06 
0.0 -1.024 0 -2.0 1e-06 
0.0 -1.0239 0 -2.0 1e-06 
0.0 -1.0238 0 -2.0 1e-06 
0.0 -1.0237 0 -2.0 1e-06 
0.0 -1.0236 0 -2.0 1e-06 
0.0 -1.0235 0 -2.0 1e-06 
0.0 -1.0234 0 -2.0 1e-06 
0.0 -1.0233 0 -2.0 1e-06 
0.0 -1.0232 0 -2.0 1e-06 
0.0 -1.0231 0 -2.0 1e-06 
0.0 -1.023 0 -2.0 1e-06 
0.0 -1.0229 0 -2.0 1e-06 
0.0 -1.0228 0 -2.0 1e-06 
0.0 -1.0227 0 -2.0 1e-06 
0.0 -1.0226 0 -2.0 1e-06 
0.0 -1.0225 0 -2.0 1e-06 
0.0 -1.0224 0 -2.0 1e-06 
0.0 -1.0223 0 -2.0 1e-06 
0.0 -1.0222 0 -2.0 1e-06 
0.0 -1.0221 0 -2.0 1e-06 
0.0 -1.022 0 -2.0 1e-06 
0.0 -1.0219 0 -2.0 1e-06 
0.0 -1.0218 0 -2.0 1e-06 
0.0 -1.0217 0 -2.0 1e-06 
0.0 -1.0216 0 -2.0 1e-06 
0.0 -1.0215 0 -2.0 1e-06 
0.0 -1.0214 0 -2.0 1e-06 
0.0 -1.0213 0 -2.0 1e-06 
0.0 -1.0212 0 -2.0 1e-06 
0.0 -1.0211 0 -2.0 1e-06 
0.0 -1.021 0 -2.0 1e-06 
0.0 -1.0209 0 -2.0 1e-06 
0.0 -1.0208 0 -2.0 1e-06 
0.0 -1.0207 0 -2.0 1e-06 
0.0 -1.0206 0 -2.0 1e-06 
0.0 -1.0205 0 -2.0 1e-06 
0.0 -1.0204 0 -2.0 1e-06 
0.0 -1.0203 0 -2.0 1e-06 
0.0 -1.0202 0 -2.0 1e-06 
0.0 -1.0201 0 -2.0 1e-06 
0.0 -1.02 0 -2.0 1e-06 
0.0 -1.0199 0 -2.0 1e-06 
0.0 -1.0198 0 -2.0 1e-06 
0.0 -1.0197 0 -2.0 1e-06 
0.0 -1.0196 0 -2.0 1e-06 
0.0 -1.0195 0 -2.0 1e-06 
0.0 -1.0194 0 -2.0 1e-06 
0.0 -1.0193 0 -2.0 1e-06 
0.0 -1.0192 0 -2.0 1e-06 
0.0 -1.0191 0 -2.0 1e-06 
0.0 -1.019 0 -2.0 1e-06 
0.0 -1.0189 0 -2.0 1e-06 
0.0 -1.0188 0 -2.0 1e-06 
0.0 -1.0187 0 -2.0 1e-06 
0.0 -1.0186 0 -2.0 1e-06 
0.0 -1.0185 0 -2.0 1e-06 
0.0 -1.0184 0 -2.0 1e-06 
0.0 -1.0183 0 -2.0 1e-06 
0.0 -1.0182 0 -2.0 1e-06 
0.0 -1.0181 0 -2.0 1e-06 
0.0 -1.018 0 -2.0 1e-06 
0.0 -1.0179 0 -2.0 1e-06 
0.0 -1.0178 0 -2.0 1e-06 
0.0 -1.0177 0 -2.0 1e-06 
0.0 -1.0176 0 -2.0 1e-06 
0.0 -1.0175 0 -2.0 1e-06 
0.0 -1.0174 0 -2.0 1e-06 
0.0 -1.0173 0 -2.0 1e-06 
0.0 -1.0172 0 -2.0 1e-06 
0.0 -1.0171 0 -2.0 1e-06 
0.0 -1.017 0 -2.0 1e-06 
0.0 -1.0169 0 -2.0 1e-06 
0.0 -1.0168 0 -2.0 1e-06 
0.0 -1.0167 0 -2.0 1e-06 
0.0 -1.0166 0 -2.0 1e-06 
0.0 -1.0165 0 -2.0 1e-06 
0.0 -1.0164 0 -2.0 1e-06 
0.0 -1.0163 0 -2.0 1e-06 
0.0 -1.0162 0 -2.0 1e-06 
0.0 -1.0161 0 -2.0 1e-06 
0.0 -1.016 0 -2.0 1e-06 
0.0 -1.0159 0 -2.0 1e-06 
0.0 -1.0158 0 -2.0 1e-06 
0.0 -1.0157 0 -2.0 1e-06 
0.0 -1.0156 0 -2.0 1e-06 
0.0 -1.0155 0 -2.0 1e-06 
0.0 -1.0154 0 -2.0 1e-06 
0.0 -1.0153 0 -2.0 1e-06 
0.0 -1.0152 0 -2.0 1e-06 
0.0 -1.0151 0 -2.0 1e-06 
0.0 -1.015 0 -2.0 1e-06 
0.0 -1.0149 0 -2.0 1e-06 
0.0 -1.0148 0 -2.0 1e-06 
0.0 -1.0147 0 -2.0 1e-06 
0.0 -1.0146 0 -2.0 1e-06 
0.0 -1.0145 0 -2.0 1e-06 
0.0 -1.0144 0 -2.0 1e-06 
0.0 -1.0143 0 -2.0 1e-06 
0.0 -1.0142 0 -2.0 1e-06 
0.0 -1.0141 0 -2.0 1e-06 
0.0 -1.014 0 -2.0 1e-06 
0.0 -1.0139 0 -2.0 1e-06 
0.0 -1.0138 0 -2.0 1e-06 
0.0 -1.0137 0 -2.0 1e-06 
0.0 -1.0136 0 -2.0 1e-06 
0.0 -1.0135 0 -2.0 1e-06 
0.0 -1.0134 0 -2.0 1e-06 
0.0 -1.0133 0 -2.0 1e-06 
0.0 -1.0132 0 -2.0 1e-06 
0.0 -1.0131 0 -2.0 1e-06 
0.0 -1.013 0 -2.0 1e-06 
0.0 -1.0129 0 -2.0 1e-06 
0.0 -1.0128 0 -2.0 1e-06 
0.0 -1.0127 0 -2.0 1e-06 
0.0 -1.0126 0 -2.0 1e-06 
0.0 -1.0125 0 -2.0 1e-06 
0.0 -1.0124 0 -2.0 1e-06 
0.0 -1.0123 0 -2.0 1e-06 
0.0 -1.0122 0 -2.0 1e-06 
0.0 -1.0121 0 -2.0 1e-06 
0.0 -1.012 0 -2.0 1e-06 
0.0 -1.0119 0 -2.0 1e-06 
0.0 -1.0118 0 -2.0 1e-06 
0.0 -1.0117 0 -2.0 1e-06 
0.0 -1.0116 0 -2.0 1e-06 
0.0 -1.0115 0 -2.0 1e-06 
0.0 -1.0114 0 -2.0 1e-06 
0.0 -1.0113 0 -2.0 1e-06 
0.0 -1.0112 0 -2.0 1e-06 
0.0 -1.0111 0 -2.0 1e-06 
0.0 -1.011 0 -2.0 1e-06 
0.0 -1.0109 0 -2.0 1e-06 
0.0 -1.0108 0 -2.0 1e-06 
0.0 -1.0107 0 -2.0 1e-06 
0.0 -1.0106 0 -2.0 1e-06 
0.0 -1.0105 0 -2.0 1e-06 
0.0 -1.0104 0 -2.0 1e-06 
0.0 -1.0103 0 -2.0 1e-06 
0.0 -1.0102 0 -2.0 1e-06 
0.0 -1.0101 0 -2.0 1e-06 
0.0 -1.01 0 -2.0 1e-06 
0.0 -1.0099 0 -2.0 1e-06 
0.0 -1.0098 0 -2.0 1e-06 
0.0 -1.0097 0 -2.0 1e-06 
0.0 -1.0096 0 -2.0 1e-06 
0.0 -1.0095 0 -2.0 1e-06 
0.0 -1.0094 0 -2.0 1e-06 
0.0 -1.0093 0 -2.0 1e-06 
0.0 -1.0092 0 -2.0 1e-06 
0.0 -1.0091 0 -2.0 1e-06 
0.0 -1.009 0 -2.0 1e-06 
0.0 -1.0089 0 -2.0 1e-06 
0.0 -1.0088 0 -2.0 1e-06 
0.0 -1.0087 0 -2.0 1e-06 
0.0 -1.0086 0 -2.0 1e-06 
0.0 -1.0085 0 -2.0 1e-06 
0.0 -1.0084 0 -2.0 1e-06 
0.0 -1.0083 0 -2.0 1e-06 
0.0 -1.0082 0 -2.0 1e-06 
0.0 -1.0081 0 -2.0 1e-06 
0.0 -1.008 0 -2.0 1e-06 
0.0 -1.0079 0 -2.0 1e-06 
0.0 -1.0078 0 -2.0 1e-06 
0.0 -1.0077 0 -2.0 1e-06 
0.0 -1.0076 0 -2.0 1e-06 
0.0 -1.0075 0 -2.0 1e-06 
0.0 -1.0074 0 -2.0 1e-06 
0.0 -1.0073 0 -2.0 1e-06 
0.0 -1.0072 0 -2.0 1e-06 
0.0 -1.0071 0 -2.0 1e-06 
0.0 -1.007 0 -2.0 1e-06 
0.0 -1.0069 0 -2.0 1e-06 
0.0 -1.0068 0 -2.0 1e-06 
0.0 -1.0067 0 -2.0 1e-06 
0.0 -1.0066 0 -2.0 1e-06 
0.0 -1.0065 0 -2.0 1e-06 
0.0 -1.0064 0 -2.0 1e-06 
0.0 -1.0063 0 -2.0 1e-06 
0.0 -1.0062 0 -2.0 1e-06 
0.0 -1.0061 0 -2.0 1e-06 
0.0 -1.006 0 -2.0 1e-06 
0.0 -1.0059 0 -2.0 1e-06 
0.0 -1.0058 0 -2.0 1e-06 
0.0 -1.0057 0 -2.0 1e-06 
0.0 -1.0056 0 -2.0 1e-06 
0.0 -1.0055 0 -2.0 1e-06 
0.0 -1.0054 0 -2.0 1e-06 
0.0 -1.0053 0 -2.0 1e-06 
0.0 -1.0052 0 -2.0 1e-06 
0.0 -1.0051 0 -2.0 1e-06 
0.0 -1.005 0 -2.0 1e-06 
0.0 -1.0049 0 -2.0 1e-06 
0.0 -1.0048 0 -2.0 1e-06 
0.0 -1.0047 0 -2.0 1e-06 
0.0 -1.0046 0 -2.0 1e-06 
0.0 -1.0045 0 -2.0 1e-06 
0.0 -1.0044 0 -2.0 1e-06 
0.0 -1.0043 0 -2.0 1e-06 
0.0 -1.0042 0 -2.0 1e-06 
0.0 -1.0041 0 -2.0 1e-06 
0.0 -1.004 0 -2.0 1e-06 
0.0 -1.0039 0 -2.0 1e-06 
0.0 -1.0038 0 -2.0 1e-06 
0.0 -1.0037 0 -2.0 1e-06 
0.0 -1.0036 0 -2.0 1e-06 
0.0 -1.0035 0 -2.0 1e-06 
0.0 -1.0034 0 -2.0 1e-06 
0.0 -1.0033 0 -2.0 1e-06 
0.0 -1.0032 0 -2.0 1e-06 
0.0 -1.0031 0 -2.0 1e-06 
0.0 -1.003 0 -2.0 1e-06 
0.0 -1.0029 0 -2.0 1e-06 
0.0 -1.0028 0 -2.0 1e-06 
0.0 -1.0027 0 -2.0 1e-06 
0.0 -1.0026 0 -2.0 1e-06 
0.0 -1.0025 0 -2.0 1e-06 
0.0 -1.0024 0 -2.0 1e-06 
0.0 -1.0023 0 -2.0 1e-06 
0.0 -1.0022 0 -2.0 1e-06 
0.0 -1.0021 0 -2.0 1e-06 
0.0 -1.002 0 -2.0 1e-06 
0.0 -1.0019 0 -2.0 1e-06 
0.0 -1.0018 0 -2.0 1e-06 
0.0 -1.0017 0 -2.0 1e-06 
0.0 -1.0016 0 -2.0 1e-06 
0.0 -1.0015 0 -2.0 1e-06 
0.0 -1.0014 0 -2.0 1e-06 
0.0 -1.0013 0 -2.0 1e-06 
0.0 -1.0012 0 -2.0 1e-06 
0.0 -1.0011 0 -2.0 1e-06 
0.0 -1.001 0 -2.0 1e-06 
0.0 -1.0009 0 -2.0 1e-06 
0.0 -1.0008 0 -2.0 1e-06 
0.0 -1.0007 0 -2.0 1e-06 
0.0 -1.0006 0 -2.0 1e-06 
0.0 -1.0005 0 -2.0 1e-06 
0.0 -1.0004 0 -2.0 1e-06 
0.0 -1.0003 0 -2.0 1e-06 
0.0 -1.0002 0 -2.0 1e-06 
0.0 -1.0001 0 -2.0 1e-06 
0.0 -1.0 0 -2.0 1e-06 
0.0 -0.9999 0 -2.0 1e-06 
0.0 -0.9998 0 -2.0 1e-06 
0.0 -0.9997 0 -2.0 1e-06 
0.0 -0.9996 0 -2.0 1e-06 
0.0 -0.9995 0 -2.0 1e-06 
0.0 -0.9994 0 -2.0 1e-06 
0.0 -0.9993 0 -2.0 1e-06 
0.0 -0.9992 0 -2.0 1e-06 
0.0 -0.9991 0 -2.0 1e-06 
0.0 -0.999 0 -2.0 1e-06 
0.0 -0.9989 0 -2.0 1e-06 
0.0 -0.9988 0 -2.0 1e-06 
0.0 -0.9987 0 -2.0 1e-06 
0.0 -0.9986 0 -2.0 1e-06 
0.0 -0.9985 0 -2.0 1e-06 
0.0 -0.9984 0 -2.0 1e-06 
0.0 -0.9983 0 -2.0 1e-06 
0.0 -0.9982 0 -2.0 1e-06 
0.0 -0.9981 0 -2.0 1e-06 
0.0 -0.998 0 -2.0 1e-06 
0.0 -0.9979 0 -2.0 1e-06 
0.0 -0.9978 0 -2.0 1e-06 
0.0 -0.9977 0 -2.0 1e-06 
0.0 -0.9976 0 -2.0 1e-06 
0.0 -0.9975 0 -2.0 1e-06 
0.0 -0.9974 0 -2.0 1e-06 
0.0 -0.9973 0 -2.0 1e-06 
0.0 -0.9972 0 -2.0 1e-06 
0.0 -0.9971 0 -2.0 1e-06 
0.0 -0.997 0 -2.0 1e-06 
0.0 -0.9969 0 -2.0 1e-06 
0.0 -0.9968 0 -2.0 1e-06 
0.0 -0.9967 0 -2.0 1e-06 
0.0 -0.9966 0 -2.0 1e-06 
0.0 -0.9965 0 -2.0 1e-06 
0.0 -0.9964 0 -2.0 1e-06 
0.0 -0.9963 0 -2.0 1e-06 
0.0 -0.9962 0 -2.0 1e-06 
0.0 -0.9961 0 -2.0 1e-06 
0.0 -0.996 0 -2.0 1e-06 
0.0 -0.9959 0 -2.0 1e-06 
0.0 -0.9958 0 -2.0 1e-06 
0.0 -0.9957 0 -2.0 1e-06 
0.0 -0.9956 0 -2.0 1e-06 
0.0 -0.9955 0 -2.0 1e-06 
0.0 -0.9954 0 -2.0 1e-06 
0.0 -0.9953 0 -2.0 1e-06 
0.0 -0.9952 0 -2.0 1e-06 
0.0 -0.9951 0 -2.0 1e-06 
0.0 -0.995 0 -2.0 1e-06 
0.0 -0.9949 0 -2.0 1e-06 
0.0 -0.9948 0 -2.0 1e-06 
0.0 -0.9947 0 -2.0 1e-06 
0.0 -0.9946 0 -2.0 1e-06 
0.0 -0.9945 0 -2.0 1e-06 
0.0 -0.9944 0 -2.0 1e-06 
0.0 -0.9943 0 -2.0 1e-06 
0.0 -0.9942 0 -2.0 1e-06 
0.0 -0.9941 0 -2.0 1e-06 
0.0 -0.994 0 -2.0 1e-06 
0.0 -0.9939 0 -2.0 1e-06 
0.0 -0.9938 0 -2.0 1e-06 
0.0 -0.9937 0 -2.0 1e-06 
0.0 -0.9936 0 -2.0 1e-06 
0.0 -0.9935 0 -2.0 1e-06 
0.0 -0.9934 0 -2.0 1e-06 
0.0 -0.9933 0 -2.0 1e-06 
0.0 -0.9932 0 -2.0 1e-06 
0.0 -0.9931 0 -2.0 1e-06 
0.0 -0.993 0 -2.0 1e-06 
0.0 -0.9929 0 -2.0 1e-06 
0.0 -0.9928 0 -2.0 1e-06 
0.0 -0.9927 0 -2.0 1e-06 
0.0 -0.9926 0 -2.0 1e-06 
0.0 -0.9925 0 -2.0 1e-06 
0.0 -0.9924 0 -2.0 1e-06 
0.0 -0.9923 0 -2.0 1e-06 
0.0 -0.9922 0 -2.0 1e-06 
0.0 -0.9921 0 -2.0 1e-06 
0.0 -0.992 0 -2.0 1e-06 
0.0 -0.9919 0 -2.0 1e-06 
0.0 -0.9918 0 -2.0 1e-06 
0.0 -0.9917 0 -2.0 1e-06 
0.0 -0.9916 0 -2.0 1e-06 
0.0 -0.9915 0 -2.0 1e-06 
0.0 -0.9914 0 -2.0 1e-06 
0.0 -0.9913 0 -2.0 1e-06 
0.0 -0.9912 0 -2.0 1e-06 
0.0 -0.9911 0 -2.0 1e-06 
0.0 -0.991 0 -2.0 1e-06 
0.0 -0.9909 0 -2.0 1e-06 
0.0 -0.9908 0 -2.0 1e-06 
0.0 -0.9907 0 -2.0 1e-06 
0.0 -0.9906 0 -2.0 1e-06 
0.0 -0.9905 0 -2.0 1e-06 
0.0 -0.9904 0 -2.0 1e-06 
0.0 -0.9903 0 -2.0 1e-06 
0.0 -0.9902 0 -2.0 1e-06 
0.0 -0.9901 0 -2.0 1e-06 
0.0 -0.99 0 -2.0 1e-06 
0.0 -0.9899 0 -2.0 1e-06 
0.0 -0.9898 0 -2.0 1e-06 
0.0 -0.9897 0 -2.0 1e-06 
0.0 -0.9896 0 -2.0 1e-06 
0.0 -0.9895 0 -2.0 1e-06 
0.0 -0.9894 0 -2.0 1e-06 
0.0 -0.9893 0 -2.0 1e-06 
0.0 -0.9892 0 -2.0 1e-06 
0.0 -0.9891 0 -2.0 1e-06 
0.0 -0.989 0 -2.0 1e-06 
0.0 -0.9889 0 -2.0 1e-06 
0.0 -0.9888 0 -2.0 1e-06 
0.0 -0.9887 0 -2.0 1e-06 
0.0 -0.9886 0 -2.0 1e-06 
0.0 -0.9885 0 -2.0 1e-06 
0.0 -0.9884 0 -2.0 1e-06 
0.0 -0.9883 0 -2.0 1e-06 
0.0 -0.9882 0 -2.0 1e-06 
0.0 -0.9881 0 -2.0 1e-06 
0.0 -0.988 0 -2.0 1e-06 
0.0 -0.9879 0 -2.0 1e-06 
0.0 -0.9878 0 -2.0 1e-06 
0.0 -0.9877 0 -2.0 1e-06 
0.0 -0.9876 0 -2.0 1e-06 
0.0 -0.9875 0 -2.0 1e-06 
0.0 -0.9874 0 -2.0 1e-06 
0.0 -0.9873 0 -2.0 1e-06 
0.0 -0.9872 0 -2.0 1e-06 
0.0 -0.9871 0 -2.0 1e-06 
0.0 -0.987 0 -2.0 1e-06 
0.0 -0.9869 0 -2.0 1e-06 
0.0 -0.9868 0 -2.0 1e-06 
0.0 -0.9867 0 -2.0 1e-06 
0.0 -0.9866 0 -2.0 1e-06 
0.0 -0.9865 0 -2.0 1e-06 
0.0 -0.9864 0 -2.0 1e-06 
0.0 -0.9863 0 -2.0 1e-06 
0.0 -0.9862 0 -2.0 1e-06 
0.0 -0.9861 0 -2.0 1e-06 
0.0 -0.986 0 -2.0 1e-06 
0.0 -0.9859 0 -2.0 1e-06 
0.0 -0.9858 0 -2.0 1e-06 
0.0 -0.9857 0 -2.0 1e-06 
0.0 -0.9856 0 -2.0 1e-06 
0.0 -0.9855 0 -2.0 1e-06 
0.0 -0.9854 0 -2.0 1e-06 
0.0 -0.9853 0 -2.0 1e-06 
0.0 -0.9852 0 -2.0 1e-06 
0.0 -0.9851 0 -2.0 1e-06 
0.0 -0.985 0 -2.0 1e-06 
0.0 -0.9849 0 -2.0 1e-06 
0.0 -0.9848 0 -2.0 1e-06 
0.0 -0.9847 0 -2.0 1e-06 
0.0 -0.9846 0 -2.0 1e-06 
0.0 -0.9845 0 -2.0 1e-06 
0.0 -0.9844 0 -2.0 1e-06 
0.0 -0.9843 0 -2.0 1e-06 
0.0 -0.9842 0 -2.0 1e-06 
0.0 -0.9841 0 -2.0 1e-06 
0.0 -0.984 0 -2.0 1e-06 
0.0 -0.9839 0 -2.0 1e-06 
0.0 -0.9838 0 -2.0 1e-06 
0.0 -0.9837 0 -2.0 1e-06 
0.0 -0.9836 0 -2.0 1e-06 
0.0 -0.9835 0 -2.0 1e-06 
0.0 -0.9834 0 -2.0 1e-06 
0.0 -0.9833 0 -2.0 1e-06 
0.0 -0.9832 0 -2.0 1e-06 
0.0 -0.9831 0 -2.0 1e-06 
0.0 -0.983 0 -2.0 1e-06 
0.0 -0.9829 0 -2.0 1e-06 
0.0 -0.9828 0 -2.0 1e-06 
0.0 -0.9827 0 -2.0 1e-06 
0.0 -0.9826 0 -2.0 1e-06 
0.0 -0.9825 0 -2.0 1e-06 
0.0 -0.9824 0 -2.0 1e-06 
0.0 -0.9823 0 -2.0 1e-06 
0.0 -0.9822 0 -2.0 1e-06 
0.0 -0.9821 0 -2.0 1e-06 
0.0 -0.982 0 -2.0 1e-06 
0.0 -0.9819 0 -2.0 1e-06 
0.0 -0.9818 0 -2.0 1e-06 
0.0 -0.9817 0 -2.0 1e-06 
0.0 -0.9816 0 -2.0 1e-06 
0.0 -0.9815 0 -2.0 1e-06 
0.0 -0.9814 0 -2.0 1e-06 
0.0 -0.9813 0 -2.0 1e-06 
0.0 -0.9812 0 -2.0 1e-06 
0.0 -0.9811 0 -2.0 1e-06 
0.0 -0.981 0 -2.0 1e-06 
0.0 -0.9809 0 -2.0 1e-06 
0.0 -0.9808 0 -2.0 1e-06 
0.0 -0.9807 0 -2.0 1e-06 
0.0 -0.9806 0 -2.0 1e-06 
0.0 -0.9805 0 -2.0 1e-06 
0.0 -0.9804 0 -2.0 1e-06 
0.0 -0.9803 0 -2.0 1e-06 
0.0 -0.9802 0 -2.0 1e-06 
0.0 -0.9801 0 -2.0 1e-06 
0.0 -0.98 0 -2.0 1e-06 
0.0 -0.9799 0 -2.0 1e-06 
0.0 -0.9798 0 -2.0 1e-06 
0.0 -0.9797 0 -2.0 1e-06 
0.0 -0.9796 0 -2.0 1e-06 
0.0 -0.9795 0 -2.0 1e-06 
0.0 -0.9794 0 -2.0 1e-06 
0.0 -0.9793 0 -2.0 1e-06 
0.0 -0.9792 0 -2.0 1e-06 
0.0 -0.9791 0 -2.0 1e-06 
0.0 -0.979 0 -2.0 1e-06 
0.0 -0.9789 0 -2.0 1e-06 
0.0 -0.9788 0 -2.0 1e-06 
0.0 -0.9787 0 -2.0 1e-06 
0.0 -0.9786 0 -2.0 1e-06 
0.0 -0.9785 0 -2.0 1e-06 
0.0 -0.9784 0 -2.0 1e-06 
0.0 -0.9783 0 -2.0 1e-06 
0.0 -0.9782 0 -2.0 1e-06 
0.0 -0.9781 0 -2.0 1e-06 
0.0 -0.978 0 -2.0 1e-06 
0.0 -0.9779 0 -2.0 1e-06 
0.0 -0.9778 0 -2.0 1e-06 
0.0 -0.9777 0 -2.0 1e-06 
0.0 -0.9776 0 -2.0 1e-06 
0.0 -0.9775 0 -2.0 1e-06 
0.0 -0.9774 0 -2.0 1e-06 
0.0 -0.9773 0 -2.0 1e-06 
0.0 -0.9772 0 -2.0 1e-06 
0.0 -0.9771 0 -2.0 1e-06 
0.0 -0.977 0 -2.0 1e-06 
0.0 -0.9769 0 -2.0 1e-06 
0.0 -0.9768 0 -2.0 1e-06 
0.0 -0.9767 0 -2.0 1e-06 
0.0 -0.9766 0 -2.0 1e-06 
0.0 -0.9765 0 -2.0 1e-06 
0.0 -0.9764 0 -2.0 1e-06 
0.0 -0.9763 0 -2.0 1e-06 
0.0 -0.9762 0 -2.0 1e-06 
0.0 -0.9761 0 -2.0 1e-06 
0.0 -0.976 0 -2.0 1e-06 
0.0 -0.9759 0 -2.0 1e-06 
0.0 -0.9758 0 -2.0 1e-06 
0.0 -0.9757 0 -2.0 1e-06 
0.0 -0.9756 0 -2.0 1e-06 
0.0 -0.9755 0 -2.0 1e-06 
0.0 -0.9754 0 -2.0 1e-06 
0.0 -0.9753 0 -2.0 1e-06 
0.0 -0.9752 0 -2.0 1e-06 
0.0 -0.9751 0 -2.0 1e-06 
0.0 -0.975 0 -2.0 1e-06 
0.0 -0.9749 0 -2.0 1e-06 
0.0 -0.9748 0 -2.0 1e-06 
0.0 -0.9747 0 -2.0 1e-06 
0.0 -0.9746 0 -2.0 1e-06 
0.0 -0.9745 0 -2.0 1e-06 
0.0 -0.9744 0 -2.0 1e-06 
0.0 -0.9743 0 -2.0 1e-06 
0.0 -0.9742 0 -2.0 1e-06 
0.0 -0.9741 0 -2.0 1e-06 
0.0 -0.974 0 -2.0 1e-06 
0.0 -0.9739 0 -2.0 1e-06 
0.0 -0.9738 0 -2.0 1e-06 
0.0 -0.9737 0 -2.0 1e-06 
0.0 -0.9736 0 -2.0 1e-06 
0.0 -0.9735 0 -2.0 1e-06 
0.0 -0.9734 0 -2.0 1e-06 
0.0 -0.9733 0 -2.0 1e-06 
0.0 -0.9732 0 -2.0 1e-06 
0.0 -0.9731 0 -2.0 1e-06 
0.0 -0.973 0 -2.0 1e-06 
0.0 -0.9729 0 -2.0 1e-06 
0.0 -0.9728 0 -2.0 1e-06 
0.0 -0.9727 0 -2.0 1e-06 
0.0 -0.9726 0 -2.0 1e-06 
0.0 -0.9725 0 -2.0 1e-06 
0.0 -0.9724 0 -2.0 1e-06 
0.0 -0.9723 0 -2.0 1e-06 
0.0 -0.9722 0 -2.0 1e-06 
0.0 -0.9721 0 -2.0 1e-06 
0.0 -0.972 0 -2.0 1e-06 
0.0 -0.9719 0 -2.0 1e-06 
0.0 -0.9718 0 -2.0 1e-06 
0.0 -0.9717 0 -2.0 1e-06 
0.0 -0.9716 0 -2.0 1e-06 
0.0 -0.9715 0 -2.0 1e-06 
0.0 -0.9714 0 -2.0 1e-06 
0.0 -0.9713 0 -2.0 1e-06 
0.0 -0.9712 0 -2.0 1e-06 
0.0 -0.9711 0 -2.0 1e-06 
0.0 -0.971 0 -2.0 1e-06 
0.0 -0.9709 0 -2.0 1e-06 
0.0 -0.9708 0 -2.0 1e-06 
0.0 -0.9707 0 -2.0 1e-06 
0.0 -0.9706 0 -2.0 1e-06 
0.0 -0.9705 0 -2.0 1e-06 
0.0 -0.9704 0 -2.0 1e-06 
0.0 -0.9703 0 -2.0 1e-06 
0.0 -0.9702 0 -2.0 1e-06 
0.0 -0.9701 0 -2.0 1e-06 
0.0 -0.97 0 -2.0 1e-06 
0.0 -0.9699 0 -2.0 1e-06 
0.0 -0.9698 0 -2.0 1e-06 
0.0 -0.9697 0 -2.0 1e-06 
0.0 -0.9696 0 -2.0 1e-06 
0.0 -0.9695 0 -2.0 1e-06 
0.0 -0.9694 0 -2.0 1e-06 
0.0 -0.9693 0 -2.0 1e-06 
0.0 -0.9692 0 -2.0 1e-06 
0.0 -0.9691 0 -2.0 1e-06 
0.0 -0.969 0 -2.0 1e-06 
0.0 -0.9689 0 -2.0 1e-06 
0.0 -0.9688 0 -2.0 1e-06 
0.0 -0.9687 0 -2.0 1e-06 
0.0 -0.9686 0 -2.0 1e-06 
0.0 -0.9685 0 -2.0 1e-06 
0.0 -0.9684 0 -2.0 1e-06 
0.0 -0.9683 0 -2.0 1e-06 
0.0 -0.9682 0 -2.0 1e-06 
0.0 -0.9681 0 -2.0 1e-06 
0.0 -0.968 0 -2.0 1e-06 
0.0 -0.9679 0 -2.0 1e-06 
0.0 -0.9678 0 -2.0 1e-06 
0.0 -0.9677 0 -2.0 1e-06 
0.0 -0.9676 0 -2.0 1e-06 
0.0 -0.9675 0 -2.0 1e-06 
0.0 -0.9674 0 -2.0 1e-06 
0.0 -0.9673 0 -2.0 1e-06 
0.0 -0.9672 0 -2.0 1e-06 
0.0 -0.9671 0 -2.0 1e-06 
0.0 -0.967 0 -2.0 1e-06 
0.0 -0.9669 0 -2.0 1e-06 
0.0 -0.9668 0 -2.0 1e-06 
0.0 -0.9667 0 -2.0 1e-06 
0.0 -0.9666 0 -2.0 1e-06 
0.0 -0.9665 0 -2.0 1e-06 
0.0 -0.9664 0 -2.0 1e-06 
0.0 -0.9663 0 -2.0 1e-06 
0.0 -0.9662 0 -2.0 1e-06 
0.0 -0.9661 0 -2.0 1e-06 
0.0 -0.966 0 -2.0 1e-06 
0.0 -0.9659 0 -2.0 1e-06 
0.0 -0.9658 0 -2.0 1e-06 
0.0 -0.9657 0 -2.0 1e-06 
0.0 -0.9656 0 -2.0 1e-06 
0.0 -0.9655 0 -2.0 1e-06 
0.0 -0.9654 0 -2.0 1e-06 
0.0 -0.9653 0 -2.0 1e-06 
0.0 -0.9652 0 -2.0 1e-06 
0.0 -0.9651 0 -2.0 1e-06 
0.0 -0.965 0 -2.0 1e-06 
0.0 -0.9649 0 -2.0 1e-06 
0.0 -0.9648 0 -2.0 1e-06 
0.0 -0.9647 0 -2.0 1e-06 
0.0 -0.9646 0 -2.0 1e-06 
0.0 -0.9645 0 -2.0 1e-06 
0.0 -0.9644 0 -2.0 1e-06 
0.0 -0.9643 0 -2.0 1e-06 
0.0 -0.9642 0 -2.0 1e-06 
0.0 -0.9641 0 -2.0 1e-06 
0.0 -0.964 0 -2.0 1e-06 
0.0 -0.9639 0 -2.0 1e-06 
0.0 -0.9638 0 -2.0 1e-06 
0.0 -0.9637 0 -2.0 1e-06 
0.0 -0.9636 0 -2.0 1e-06 
0.0 -0.9635 0 -2.0 1e-06 
0.0 -0.9634 0 -2.0 1e-06 
0.0 -0.9633 0 -2.0 1e-06 
0.0 -0.9632 0 -2.0 1e-06 
0.0 -0.9631 0 -2.0 1e-06 
0.0 -0.963 0 -2.0 1e-06 
0.0 -0.9629 0 -2.0 1e-06 
0.0 -0.9628 0 -2.0 1e-06 
0.0 -0.9627 0 -2.0 1e-06 
0.0 -0.9626 0 -2.0 1e-06 
0.0 -0.9625 0 -2.0 1e-06 
0.0 -0.9624 0 -2.0 1e-06 
0.0 -0.9623 0 -2.0 1e-06 
0.0 -0.9622 0 -2.0 1e-06 
0.0 -0.9621 0 -2.0 1e-06 
0.0 -0.962 0 -2.0 1e-06 
0.0 -0.9619 0 -2.0 1e-06 
0.0 -0.9618 0 -2.0 1e-06 
0.0 -0.9617 0 -2.0 1e-06 
0.0 -0.9616 0 -2.0 1e-06 
0.0 -0.9615 0 -2.0 1e-06 
0.0 -0.9614 0 -2.0 1e-06 
0.0 -0.9613 0 -2.0 1e-06 
0.0 -0.9612 0 -2.0 1e-06 
0.0 -0.9611 0 -2.0 1e-06 
0.0 -0.961 0 -2.0 1e-06 
0.0 -0.9609 0 -2.0 1e-06 
0.0 -0.9608 0 -2.0 1e-06 
0.0 -0.9607 0 -2.0 1e-06 
0.0 -0.9606 0 -2.0 1e-06 
0.0 -0.9605 0 -2.0 1e-06 
0.0 -0.9604 0 -2.0 1e-06 
0.0 -0.9603 0 -2.0 1e-06 
0.0 -0.9602 0 -2.0 1e-06 
0.0 -0.9601 0 -2.0 1e-06 
0.0 -0.96 0 -2.0 1e-06 
0.0 -0.9599 0 -2.0 1e-06 
0.0 -0.9598 0 -2.0 1e-06 
0.0 -0.9597 0 -2.0 1e-06 
0.0 -0.9596 0 -2.0 1e-06 
0.0 -0.9595 0 -2.0 1e-06 
0.0 -0.9594 0 -2.0 1e-06 
0.0 -0.9593 0 -2.0 1e-06 
0.0 -0.9592 0 -2.0 1e-06 
0.0 -0.9591 0 -2.0 1e-06 
0.0 -0.959 0 -2.0 1e-06 
0.0 -0.9589 0 -2.0 1e-06 
0.0 -0.9588 0 -2.0 1e-06 
0.0 -0.9587 0 -2.0 1e-06 
0.0 -0.9586 0 -2.0 1e-06 
0.0 -0.9585 0 -2.0 1e-06 
0.0 -0.9584 0 -2.0 1e-06 
0.0 -0.9583 0 -2.0 1e-06 
0.0 -0.9582 0 -2.0 1e-06 
0.0 -0.9581 0 -2.0 1e-06 
0.0 -0.958 0 -2.0 1e-06 
0.0 -0.9579 0 -2.0 1e-06 
0.0 -0.9578 0 -2.0 1e-06 
0.0 -0.9577 0 -2.0 1e-06 
0.0 -0.9576 0 -2.0 1e-06 
0.0 -0.9575 0 -2.0 1e-06 
0.0 -0.9574 0 -2.0 1e-06 
0.0 -0.9573 0 -2.0 1e-06 
0.0 -0.9572 0 -2.0 1e-06 
0.0 -0.9571 0 -2.0 1e-06 
0.0 -0.957 0 -2.0 1e-06 
0.0 -0.9569 0 -2.0 1e-06 
0.0 -0.9568 0 -2.0 1e-06 
0.0 -0.9567 0 -2.0 1e-06 
0.0 -0.9566 0 -2.0 1e-06 
0.0 -0.9565 0 -2.0 1e-06 
0.0 -0.9564 0 -2.0 1e-06 
0.0 -0.9563 0 -2.0 1e-06 
0.0 -0.9562 0 -2.0 1e-06 
0.0 -0.9561 0 -2.0 1e-06 
0.0 -0.956 0 -2.0 1e-06 
0.0 -0.9559 0 -2.0 1e-06 
0.0 -0.9558 0 -2.0 1e-06 
0.0 -0.9557 0 -2.0 1e-06 
0.0 -0.9556 0 -2.0 1e-06 
0.0 -0.9555 0 -2.0 1e-06 
0.0 -0.9554 0 -2.0 1e-06 
0.0 -0.9553 0 -2.0 1e-06 
0.0 -0.9552 0 -2.0 1e-06 
0.0 -0.9551 0 -2.0 1e-06 
0.0 -0.955 0 -2.0 1e-06 
0.0 -0.9549 0 -2.0 1e-06 
0.0 -0.9548 0 -2.0 1e-06 
0.0 -0.9547 0 -2.0 1e-06 
0.0 -0.9546 0 -2.0 1e-06 
0.0 -0.9545 0 -2.0 1e-06 
0.0 -0.9544 0 -2.0 1e-06 
0.0 -0.9543 0 -2.0 1e-06 
0.0 -0.9542 0 -2.0 1e-06 
0.0 -0.9541 0 -2.0 1e-06 
0.0 -0.954 0 -2.0 1e-06 
0.0 -0.9539 0 -2.0 1e-06 
0.0 -0.9538 0 -2.0 1e-06 
0.0 -0.9537 0 -2.0 1e-06 
0.0 -0.9536 0 -2.0 1e-06 
0.0 -0.9535 0 -2.0 1e-06 
0.0 -0.9534 0 -2.0 1e-06 
0.0 -0.9533 0 -2.0 1e-06 
0.0 -0.9532 0 -2.0 1e-06 
0.0 -0.9531 0 -2.0 1e-06 
0.0 -0.953 0 -2.0 1e-06 
0.0 -0.9529 0 -2.0 1e-06 
0.0 -0.9528 0 -2.0 1e-06 
0.0 -0.9527 0 -2.0 1e-06 
0.0 -0.9526 0 -2.0 1e-06 
0.0 -0.9525 0 -2.0 1e-06 
0.0 -0.9524 0 -2.0 1e-06 
0.0 -0.9523 0 -2.0 1e-06 
0.0 -0.9522 0 -2.0 1e-06 
0.0 -0.9521 0 -2.0 1e-06 
0.0 -0.952 0 -2.0 1e-06 
0.0 -0.9519 0 -2.0 1e-06 
0.0 -0.9518 0 -2.0 1e-06 
0.0 -0.9517 0 -2.0 1e-06 
0.0 -0.9516 0 -2.0 1e-06 
0.0 -0.9515 0 -2.0 1e-06 
0.0 -0.9514 0 -2.0 1e-06 
0.0 -0.9513 0 -2.0 1e-06 
0.0 -0.9512 0 -2.0 1e-06 
0.0 -0.9511 0 -2.0 1e-06 
0.0 -0.951 0 -2.0 1e-06 
0.0 -0.9509 0 -2.0 1e-06 
0.0 -0.9508 0 -2.0 1e-06 
0.0 -0.9507 0 -2.0 1e-06 
0.0 -0.9506 0 -2.0 1e-06 
0.0 -0.9505 0 -2.0 1e-06 
0.0 -0.9504 0 -2.0 1e-06 
0.0 -0.9503 0 -2.0 1e-06 
0.0 -0.9502 0 -2.0 1e-06 
0.0 -0.9501 0 -2.0 1e-06 
0.0 -0.95 0 -2.0 1e-06 
0.0 -0.9499 0 -2.0 1e-06 
0.0 -0.9498 0 -2.0 1e-06 
0.0 -0.9497 0 -2.0 1e-06 
0.0 -0.9496 0 -2.0 1e-06 
0.0 -0.9495 0 -2.0 1e-06 
0.0 -0.9494 0 -2.0 1e-06 
0.0 -0.9493 0 -2.0 1e-06 
0.0 -0.9492 0 -2.0 1e-06 
0.0 -0.9491 0 -2.0 1e-06 
0.0 -0.949 0 -2.0 1e-06 
0.0 -0.9489 0 -2.0 1e-06 
0.0 -0.9488 0 -2.0 1e-06 
0.0 -0.9487 0 -2.0 1e-06 
0.0 -0.9486 0 -2.0 1e-06 
0.0 -0.9485 0 -2.0 1e-06 
0.0 -0.9484 0 -2.0 1e-06 
0.0 -0.9483 0 -2.0 1e-06 
0.0 -0.9482 0 -2.0 1e-06 
0.0 -0.9481 0 -2.0 1e-06 
0.0 -0.948 0 -2.0 1e-06 
0.0 -0.9479 0 -2.0 1e-06 
0.0 -0.9478 0 -2.0 1e-06 
0.0 -0.9477 0 -2.0 1e-06 
0.0 -0.9476 0 -2.0 1e-06 
0.0 -0.9475 0 -2.0 1e-06 
0.0 -0.9474 0 -2.0 1e-06 
0.0 -0.9473 0 -2.0 1e-06 
0.0 -0.9472 0 -2.0 1e-06 
0.0 -0.9471 0 -2.0 1e-06 
0.0 -0.947 0 -2.0 1e-06 
0.0 -0.9469 0 -2.0 1e-06 
0.0 -0.9468 0 -2.0 1e-06 
0.0 -0.9467 0 -2.0 1e-06 
0.0 -0.9466 0 -2.0 1e-06 
0.0 -0.9465 0 -2.0 1e-06 
0.0 -0.9464 0 -2.0 1e-06 
0.0 -0.9463 0 -2.0 1e-06 
0.0 -0.9462 0 -2.0 1e-06 
0.0 -0.9461 0 -2.0 1e-06 
0.0 -0.946 0 -2.0 1e-06 
0.0 -0.9459 0 -2.0 1e-06 
0.0 -0.9458 0 -2.0 1e-06 
0.0 -0.9457 0 -2.0 1e-06 
0.0 -0.9456 0 -2.0 1e-06 
0.0 -0.9455 0 -2.0 1e-06 
0.0 -0.9454 0 -2.0 1e-06 
0.0 -0.9453 0 -2.0 1e-06 
0.0 -0.9452 0 -2.0 1e-06 
0.0 -0.9451 0 -2.0 1e-06 
0.0 -0.945 0 -2.0 1e-06 
0.0 -0.9449 0 -2.0 1e-06 
0.0 -0.9448 0 -2.0 1e-06 
0.0 -0.9447 0 -2.0 1e-06 
0.0 -0.9446 0 -2.0 1e-06 
0.0 -0.9445 0 -2.0 1e-06 
0.0 -0.9444 0 -2.0 1e-06 
0.0 -0.9443 0 -2.0 1e-06 
0.0 -0.9442 0 -2.0 1e-06 
0.0 -0.9441 0 -2.0 1e-06 
0.0 -0.944 0 -2.0 1e-06 
0.0 -0.9439 0 -2.0 1e-06 
0.0 -0.9438 0 -2.0 1e-06 
0.0 -0.9437 0 -2.0 1e-06 
0.0 -0.9436 0 -2.0 1e-06 
0.0 -0.9435 0 -2.0 1e-06 
0.0 -0.9434 0 -2.0 1e-06 
0.0 -0.9433 0 -2.0 1e-06 
0.0 -0.9432 0 -2.0 1e-06 
0.0 -0.9431 0 -2.0 1e-06 
0.0 -0.943 0 -2.0 1e-06 
0.0 -0.9429 0 -2.0 1e-06 
0.0 -0.9428 0 -2.0 1e-06 
0.0 -0.9427 0 -2.0 1e-06 
0.0 -0.9426 0 -2.0 1e-06 
0.0 -0.9425 0 -2.0 1e-06 
0.0 -0.9424 0 -2.0 1e-06 
0.0 -0.9423 0 -2.0 1e-06 
0.0 -0.9422 0 -2.0 1e-06 
0.0 -0.9421 0 -2.0 1e-06 
0.0 -0.942 0 -2.0 1e-06 
0.0 -0.9419 0 -2.0 1e-06 
0.0 -0.9418 0 -2.0 1e-06 
0.0 -0.9417 0 -2.0 1e-06 
0.0 -0.9416 0 -2.0 1e-06 
0.0 -0.9415 0 -2.0 1e-06 
0.0 -0.9414 0 -2.0 1e-06 
0.0 -0.9413 0 -2.0 1e-06 
0.0 -0.9412 0 -2.0 1e-06 
0.0 -0.9411 0 -2.0 1e-06 
0.0 -0.941 0 -2.0 1e-06 
0.0 -0.9409 0 -2.0 1e-06 
0.0 -0.9408 0 -2.0 1e-06 
0.0 -0.9407 0 -2.0 1e-06 
0.0 -0.9406 0 -2.0 1e-06 
0.0 -0.9405 0 -2.0 1e-06 
0.0 -0.9404 0 -2.0 1e-06 
0.0 -0.9403 0 -2.0 1e-06 
0.0 -0.9402 0 -2.0 1e-06 
0.0 -0.9401 0 -2.0 1e-06 
0.0 -0.94 0 -2.0 1e-06 
0.0 -0.9399 0 -2.0 1e-06 
0.0 -0.9398 0 -2.0 1e-06 
0.0 -0.9397 0 -2.0 1e-06 
0.0 -0.9396 0 -2.0 1e-06 
0.0 -0.9395 0 -2.0 1e-06 
0.0 -0.9394 0 -2.0 1e-06 
0.0 -0.9393 0 -2.0 1e-06 
0.0 -0.9392 0 -2.0 1e-06 
0.0 -0.9391 0 -2.0 1e-06 
0.0 -0.939 0 -2.0 1e-06 
0.0 -0.9389 0 -2.0 1e-06 
0.0 -0.9388 0 -2.0 1e-06 
0.0 -0.9387 0 -2.0 1e-06 
0.0 -0.9386 0 -2.0 1e-06 
0.0 -0.9385 0 -2.0 1e-06 
0.0 -0.9384 0 -2.0 1e-06 
0.0 -0.9383 0 -2.0 1e-06 
0.0 -0.9382 0 -2.0 1e-06 
0.0 -0.9381 0 -2.0 1e-06 
0.0 -0.938 0 -2.0 1e-06 
0.0 -0.9379 0 -2.0 1e-06 
0.0 -0.9378 0 -2.0 1e-06 
0.0 -0.9377 0 -2.0 1e-06 
0.0 -0.9376 0 -2.0 1e-06 
0.0 -0.9375 0 -2.0 1e-06 
0.0 -0.9374 0 -2.0 1e-06 
0.0 -0.9373 0 -2.0 1e-06 
0.0 -0.9372 0 -2.0 1e-06 
0.0 -0.9371 0 -2.0 1e-06 
0.0 -0.937 0 -2.0 1e-06 
0.0 -0.9369 0 -2.0 1e-06 
0.0 -0.9368 0 -2.0 1e-06 
0.0 -0.9367 0 -2.0 1e-06 
0.0 -0.9366 0 -2.0 1e-06 
0.0 -0.9365 0 -2.0 1e-06 
0.0 -0.9364 0 -2.0 1e-06 
0.0 -0.9363 0 -2.0 1e-06 
0.0 -0.9362 0 -2.0 1e-06 
0.0 -0.9361 0 -2.0 1e-06 
0.0 -0.936 0 -2.0 1e-06 
0.0 -0.9359 0 -2.0 1e-06 
0.0 -0.9358 0 -2.0 1e-06 
0.0 -0.9357 0 -2.0 1e-06 
0.0 -0.9356 0 -2.0 1e-06 
0.0 -0.9355 0 -2.0 1e-06 
0.0 -0.9354 0 -2.0 1e-06 
0.0 -0.9353 0 -2.0 1e-06 
0.0 -0.9352 0 -2.0 1e-06 
0.0 -0.9351 0 -2.0 1e-06 
0.0 -0.935 0 -2.0 1e-06 
0.0 -0.9349 0 -2.0 1e-06 
0.0 -0.9348 0 -2.0 1e-06 
0.0 -0.9347 0 -2.0 1e-06 
0.0 -0.9346 0 -2.0 1e-06 
0.0 -0.9345 0 -2.0 1e-06 
0.0 -0.9344 0 -2.0 1e-06 
0.0 -0.9343 0 -2.0 1e-06 
0.0 -0.9342 0 -2.0 1e-06 
0.0 -0.9341 0 -2.0 1e-06 
0.0 -0.934 0 -2.0 1e-06 
0.0 -0.9339 0 -2.0 1e-06 
0.0 -0.9338 0 -2.0 1e-06 
0.0 -0.9337 0 -2.0 1e-06 
0.0 -0.9336 0 -2.0 1e-06 
0.0 -0.9335 0 -2.0 1e-06 
0.0 -0.9334 0 -2.0 1e-06 
0.0 -0.9333 0 -2.0 1e-06 
0.0 -0.9332 0 -2.0 1e-06 
0.0 -0.9331 0 -2.0 1e-06 
0.0 -0.933 0 -2.0 1e-06 
0.0 -0.9329 0 -2.0 1e-06 
0.0 -0.9328 0 -2.0 1e-06 
0.0 -0.9327 0 -2.0 1e-06 
0.0 -0.9326 0 -2.0 1e-06 
0.0 -0.9325 0 -2.0 1e-06 
0.0 -0.9324 0 -2.0 1e-06 
0.0 -0.9323 0 -2.0 1e-06 
0.0 -0.9322 0 -2.0 1e-06 
0.0 -0.9321 0 -2.0 1e-06 
0.0 -0.932 0 -2.0 1e-06 
0.0 -0.9319 0 -2.0 1e-06 
0.0 -0.9318 0 -2.0 1e-06 
0.0 -0.9317 0 -2.0 1e-06 
0.0 -0.9316 0 -2.0 1e-06 
0.0 -0.9315 0 -2.0 1e-06 
0.0 -0.9314 0 -2.0 1e-06 
0.0 -0.9313 0 -2.0 1e-06 
0.0 -0.9312 0 -2.0 1e-06 
0.0 -0.9311 0 -2.0 1e-06 
0.0 -0.931 0 -2.0 1e-06 
0.0 -0.9309 0 -2.0 1e-06 
0.0 -0.9308 0 -2.0 1e-06 
0.0 -0.9307 0 -2.0 1e-06 
0.0 -0.9306 0 -2.0 1e-06 
0.0 -0.9305 0 -2.0 1e-06 
0.0 -0.9304 0 -2.0 1e-06 
0.0 -0.9303 0 -2.0 1e-06 
0.0 -0.9302 0 -2.0 1e-06 
0.0 -0.9301 0 -2.0 1e-06 
0.0 -0.93 0 -2.0 1e-06 
0.0 -0.9299 0 -2.0 1e-06 
0.0 -0.9298 0 -2.0 1e-06 
0.0 -0.9297 0 -2.0 1e-06 
0.0 -0.9296 0 -2.0 1e-06 
0.0 -0.9295 0 -2.0 1e-06 
0.0 -0.9294 0 -2.0 1e-06 
0.0 -0.9293 0 -2.0 1e-06 
0.0 -0.9292 0 -2.0 1e-06 
0.0 -0.9291 0 -2.0 1e-06 
0.0 -0.929 0 -2.0 1e-06 
0.0 -0.9289 0 -2.0 1e-06 
0.0 -0.9288 0 -2.0 1e-06 
0.0 -0.9287 0 -2.0 1e-06 
0.0 -0.9286 0 -2.0 1e-06 
0.0 -0.9285 0 -2.0 1e-06 
0.0 -0.9284 0 -2.0 1e-06 
0.0 -0.9283 0 -2.0 1e-06 
0.0 -0.9282 0 -2.0 1e-06 
0.0 -0.9281 0 -2.0 1e-06 
0.0 -0.928 0 -2.0 1e-06 
0.0 -0.9279 0 -2.0 1e-06 
0.0 -0.9278 0 -2.0 1e-06 
0.0 -0.9277 0 -2.0 1e-06 
0.0 -0.9276 0 -2.0 1e-06 
0.0 -0.9275 0 -2.0 1e-06 
0.0 -0.9274 0 -2.0 1e-06 
0.0 -0.9273 0 -2.0 1e-06 
0.0 -0.9272 0 -2.0 1e-06 
0.0 -0.9271 0 -2.0 1e-06 
0.0 -0.927 0 -2.0 1e-06 
0.0 -0.9269 0 -2.0 1e-06 
0.0 -0.9268 0 -2.0 1e-06 
0.0 -0.9267 0 -2.0 1e-06 
0.0 -0.9266 0 -2.0 1e-06 
0.0 -0.9265 0 -2.0 1e-06 
0.0 -0.9264 0 -2.0 1e-06 
0.0 -0.9263 0 -2.0 1e-06 
0.0 -0.9262 0 -2.0 1e-06 
0.0 -0.9261 0 -2.0 1e-06 
0.0 -0.926 0 -2.0 1e-06 
0.0 -0.9259 0 -2.0 1e-06 
0.0 -0.9258 0 -2.0 1e-06 
0.0 -0.9257 0 -2.0 1e-06 
0.0 -0.9256 0 -2.0 1e-06 
0.0 -0.9255 0 -2.0 1e-06 
0.0 -0.9254 0 -2.0 1e-06 
0.0 -0.9253 0 -2.0 1e-06 
0.0 -0.9252 0 -2.0 1e-06 
0.0 -0.9251 0 -2.0 1e-06 
0.0 -0.925 0 -2.0 1e-06 
0.0 -0.9249 0 -2.0 1e-06 
0.0 -0.9248 0 -2.0 1e-06 
0.0 -0.9247 0 -2.0 1e-06 
0.0 -0.9246 0 -2.0 1e-06 
0.0 -0.9245 0 -2.0 1e-06 
0.0 -0.9244 0 -2.0 1e-06 
0.0 -0.9243 0 -2.0 1e-06 
0.0 -0.9242 0 -2.0 1e-06 
0.0 -0.9241 0 -2.0 1e-06 
0.0 -0.924 0 -2.0 1e-06 
0.0 -0.9239 0 -2.0 1e-06 
0.0 -0.9238 0 -2.0 1e-06 
0.0 -0.9237 0 -2.0 1e-06 
0.0 -0.9236 0 -2.0 1e-06 
0.0 -0.9235 0 -2.0 1e-06 
0.0 -0.9234 0 -2.0 1e-06 
0.0 -0.9233 0 -2.0 1e-06 
0.0 -0.9232 0 -2.0 1e-06 
0.0 -0.9231 0 -2.0 1e-06 
0.0 -0.923 0 -2.0 1e-06 
0.0 -0.9229 0 -2.0 1e-06 
0.0 -0.9228 0 -2.0 1e-06 
0.0 -0.9227 0 -2.0 1e-06 
0.0 -0.9226 0 -2.0 1e-06 
0.0 -0.9225 0 -2.0 1e-06 
0.0 -0.9224 0 -2.0 1e-06 
0.0 -0.9223 0 -2.0 1e-06 
0.0 -0.9222 0 -2.0 1e-06 
0.0 -0.9221 0 -2.0 1e-06 
0.0 -0.922 0 -2.0 1e-06 
0.0 -0.9219 0 -2.0 1e-06 
0.0 -0.9218 0 -2.0 1e-06 
0.0 -0.9217 0 -2.0 1e-06 
0.0 -0.9216 0 -2.0 1e-06 
0.0 -0.9215 0 -2.0 1e-06 
0.0 -0.9214 0 -2.0 1e-06 
0.0 -0.9213 0 -2.0 1e-06 
0.0 -0.9212 0 -2.0 1e-06 
0.0 -0.9211 0 -2.0 1e-06 
0.0 -0.921 0 -2.0 1e-06 
0.0 -0.9209 0 -2.0 1e-06 
0.0 -0.9208 0 -2.0 1e-06 
0.0 -0.9207 0 -2.0 1e-06 
0.0 -0.9206 0 -2.0 1e-06 
0.0 -0.9205 0 -2.0 1e-06 
0.0 -0.9204 0 -2.0 1e-06 
0.0 -0.9203 0 -2.0 1e-06 
0.0 -0.9202 0 -2.0 1e-06 
0.0 -0.9201 0 -2.0 1e-06 
0.0 -0.92 0 -2.0 1e-06 
0.0 -0.9199 0 -2.0 1e-06 
0.0 -0.9198 0 -2.0 1e-06 
0.0 -0.9197 0 -2.0 1e-06 
0.0 -0.9196 0 -2.0 1e-06 
0.0 -0.9195 0 -2.0 1e-06 
0.0 -0.9194 0 -2.0 1e-06 
0.0 -0.9193 0 -2.0 1e-06 
0.0 -0.9192 0 -2.0 1e-06 
0.0 -0.9191 0 -2.0 1e-06 
0.0 -0.919 0 -2.0 1e-06 
0.0 -0.9189 0 -2.0 1e-06 
0.0 -0.9188 0 -2.0 1e-06 
0.0 -0.9187 0 -2.0 1e-06 
0.0 -0.9186 0 -2.0 1e-06 
0.0 -0.9185 0 -2.0 1e-06 
0.0 -0.9184 0 -2.0 1e-06 
0.0 -0.9183 0 -2.0 1e-06 
0.0 -0.9182 0 -2.0 1e-06 
0.0 -0.9181 0 -2.0 1e-06 
0.0 -0.918 0 -2.0 1e-06 
0.0 -0.9179 0 -2.0 1e-06 
0.0 -0.9178 0 -2.0 1e-06 
0.0 -0.9177 0 -2.0 1e-06 
0.0 -0.9176 0 -2.0 1e-06 
0.0 -0.9175 0 -2.0 1e-06 
0.0 -0.9174 0 -2.0 1e-06 
0.0 -0.9173 0 -2.0 1e-06 
0.0 -0.9172 0 -2.0 1e-06 
0.0 -0.9171 0 -2.0 1e-06 
0.0 -0.917 0 -2.0 1e-06 
0.0 -0.9169 0 -2.0 1e-06 
0.0 -0.9168 0 -2.0 1e-06 
0.0 -0.9167 0 -2.0 1e-06 
0.0 -0.9166 0 -2.0 1e-06 
0.0 -0.9165 0 -2.0 1e-06 
0.0 -0.9164 0 -2.0 1e-06 
0.0 -0.9163 0 -2.0 1e-06 
0.0 -0.9162 0 -2.0 1e-06 
0.0 -0.9161 0 -2.0 1e-06 
0.0 -0.916 0 -2.0 1e-06 
0.0 -0.9159 0 -2.0 1e-06 
0.0 -0.9158 0 -2.0 1e-06 
0.0 -0.9157 0 -2.0 1e-06 
0.0 -0.9156 0 -2.0 1e-06 
0.0 -0.9155 0 -2.0 1e-06 
0.0 -0.9154 0 -2.0 1e-06 
0.0 -0.9153 0 -2.0 1e-06 
0.0 -0.9152 0 -2.0 1e-06 
0.0 -0.9151 0 -2.0 1e-06 
0.0 -0.915 0 -2.0 1e-06 
0.0 -0.9149 0 -2.0 1e-06 
0.0 -0.9148 0 -2.0 1e-06 
0.0 -0.9147 0 -2.0 1e-06 
0.0 -0.9146 0 -2.0 1e-06 
0.0 -0.9145 0 -2.0 1e-06 
0.0 -0.9144 0 -2.0 1e-06 
0.0 -0.9143 0 -2.0 1e-06 
0.0 -0.9142 0 -2.0 1e-06 
0.0 -0.9141 0 -2.0 1e-06 
0.0 -0.914 0 -2.0 1e-06 
0.0 -0.9139 0 -2.0 1e-06 
0.0 -0.9138 0 -2.0 1e-06 
0.0 -0.9137 0 -2.0 1e-06 
0.0 -0.9136 0 -2.0 1e-06 
0.0 -0.9135 0 -2.0 1e-06 
0.0 -0.9134 0 -2.0 1e-06 
0.0 -0.9133 0 -2.0 1e-06 
0.0 -0.9132 0 -2.0 1e-06 
0.0 -0.9131 0 -2.0 1e-06 
0.0 -0.913 0 -2.0 1e-06 
0.0 -0.9129 0 -2.0 1e-06 
0.0 -0.9128 0 -2.0 1e-06 
0.0 -0.9127 0 -2.0 1e-06 
0.0 -0.9126 0 -2.0 1e-06 
0.0 -0.9125 0 -2.0 1e-06 
0.0 -0.9124 0 -2.0 1e-06 
0.0 -0.9123 0 -2.0 1e-06 
0.0 -0.9122 0 -2.0 1e-06 
0.0 -0.9121 0 -2.0 1e-06 
0.0 -0.912 0 -2.0 1e-06 
0.0 -0.9119 0 -2.0 1e-06 
0.0 -0.9118 0 -2.0 1e-06 
0.0 -0.9117 0 -2.0 1e-06 
0.0 -0.9116 0 -2.0 1e-06 
0.0 -0.9115 0 -2.0 1e-06 
0.0 -0.9114 0 -2.0 1e-06 
0.0 -0.9113 0 -2.0 1e-06 
0.0 -0.9112 0 -2.0 1e-06 
0.0 -0.9111 0 -2.0 1e-06 
0.0 -0.911 0 -2.0 1e-06 
0.0 -0.9109 0 -2.0 1e-06 
0.0 -0.9108 0 -2.0 1e-06 
0.0 -0.9107 0 -2.0 1e-06 
0.0 -0.9106 0 -2.0 1e-06 
0.0 -0.9105 0 -2.0 1e-06 
0.0 -0.9104 0 -2.0 1e-06 
0.0 -0.9103 0 -2.0 1e-06 
0.0 -0.9102 0 -2.0 1e-06 
0.0 -0.9101 0 -2.0 1e-06 
0.0 -0.91 0 -2.0 1e-06 
0.0 -0.9099 0 -2.0 1e-06 
0.0 -0.9098 0 -2.0 1e-06 
0.0 -0.9097 0 -2.0 1e-06 
0.0 -0.9096 0 -2.0 1e-06 
0.0 -0.9095 0 -2.0 1e-06 
0.0 -0.9094 0 -2.0 1e-06 
0.0 -0.9093 0 -2.0 1e-06 
0.0 -0.9092 0 -2.0 1e-06 
0.0 -0.9091 0 -2.0 1e-06 
0.0 -0.909 0 -2.0 1e-06 
0.0 -0.9089 0 -2.0 1e-06 
0.0 -0.9088 0 -2.0 1e-06 
0.0 -0.9087 0 -2.0 1e-06 
0.0 -0.9086 0 -2.0 1e-06 
0.0 -0.9085 0 -2.0 1e-06 
0.0 -0.9084 0 -2.0 1e-06 
0.0 -0.9083 0 -2.0 1e-06 
0.0 -0.9082 0 -2.0 1e-06 
0.0 -0.9081 0 -2.0 1e-06 
0.0 -0.908 0 -2.0 1e-06 
0.0 -0.9079 0 -2.0 1e-06 
0.0 -0.9078 0 -2.0 1e-06 
0.0 -0.9077 0 -2.0 1e-06 
0.0 -0.9076 0 -2.0 1e-06 
0.0 -0.9075 0 -2.0 1e-06 
0.0 -0.9074 0 -2.0 1e-06 
0.0 -0.9073 0 -2.0 1e-06 
0.0 -0.9072 0 -2.0 1e-06 
0.0 -0.9071 0 -2.0 1e-06 
0.0 -0.907 0 -2.0 1e-06 
0.0 -0.9069 0 -2.0 1e-06 
0.0 -0.9068 0 -2.0 1e-06 
0.0 -0.9067 0 -2.0 1e-06 
0.0 -0.9066 0 -2.0 1e-06 
0.0 -0.9065 0 -2.0 1e-06 
0.0 -0.9064 0 -2.0 1e-06 
0.0 -0.9063 0 -2.0 1e-06 
0.0 -0.9062 0 -2.0 1e-06 
0.0 -0.9061 0 -2.0 1e-06 
0.0 -0.906 0 -2.0 1e-06 
0.0 -0.9059 0 -2.0 1e-06 
0.0 -0.9058 0 -2.0 1e-06 
0.0 -0.9057 0 -2.0 1e-06 
0.0 -0.9056 0 -2.0 1e-06 
0.0 -0.9055 0 -2.0 1e-06 
0.0 -0.9054 0 -2.0 1e-06 
0.0 -0.9053 0 -2.0 1e-06 
0.0 -0.9052 0 -2.0 1e-06 
0.0 -0.9051 0 -2.0 1e-06 
0.0 -0.905 0 -2.0 1e-06 
0.0 -0.9049 0 -2.0 1e-06 
0.0 -0.9048 0 -2.0 1e-06 
0.0 -0.9047 0 -2.0 1e-06 
0.0 -0.9046 0 -2.0 1e-06 
0.0 -0.9045 0 -2.0 1e-06 
0.0 -0.9044 0 -2.0 1e-06 
0.0 -0.9043 0 -2.0 1e-06 
0.0 -0.9042 0 -2.0 1e-06 
0.0 -0.9041 0 -2.0 1e-06 
0.0 -0.904 0 -2.0 1e-06 
0.0 -0.9039 0 -2.0 1e-06 
0.0 -0.9038 0 -2.0 1e-06 
0.0 -0.9037 0 -2.0 1e-06 
0.0 -0.9036 0 -2.0 1e-06 
0.0 -0.9035 0 -2.0 1e-06 
0.0 -0.9034 0 -2.0 1e-06 
0.0 -0.9033 0 -2.0 1e-06 
0.0 -0.9032 0 -2.0 1e-06 
0.0 -0.9031 0 -2.0 1e-06 
0.0 -0.903 0 -2.0 1e-06 
0.0 -0.9029 0 -2.0 1e-06 
0.0 -0.9028 0 -2.0 1e-06 
0.0 -0.9027 0 -2.0 1e-06 
0.0 -0.9026 0 -2.0 1e-06 
0.0 -0.9025 0 -2.0 1e-06 
0.0 -0.9024 0 -2.0 1e-06 
0.0 -0.9023 0 -2.0 1e-06 
0.0 -0.9022 0 -2.0 1e-06 
0.0 -0.9021 0 -2.0 1e-06 
0.0 -0.902 0 -2.0 1e-06 
0.0 -0.9019 0 -2.0 1e-06 
0.0 -0.9018 0 -2.0 1e-06 
0.0 -0.9017 0 -2.0 1e-06 
0.0 -0.9016 0 -2.0 1e-06 
0.0 -0.9015 0 -2.0 1e-06 
0.0 -0.9014 0 -2.0 1e-06 
0.0 -0.9013 0 -2.0 1e-06 
0.0 -0.9012 0 -2.0 1e-06 
0.0 -0.9011 0 -2.0 1e-06 
0.0 -0.901 0 -2.0 1e-06 
0.0 -0.9009 0 -2.0 1e-06 
0.0 -0.9008 0 -2.0 1e-06 
0.0 -0.9007 0 -2.0 1e-06 
0.0 -0.9006 0 -2.0 1e-06 
0.0 -0.9005 0 -2.0 1e-06 
0.0 -0.9004 0 -2.0 1e-06 
0.0 -0.9003 0 -2.0 1e-06 
0.0 -0.9002 0 -2.0 1e-06 
0.0 -0.9001 0 -2.0 1e-06 
0.0 -0.9 0 -2.0 1e-06 
0.0 -0.8999 0 -2.0 1e-06 
0.0 -0.8998 0 -2.0 1e-06 
0.0 -0.8997 0 -2.0 1e-06 
0.0 -0.8996 0 -2.0 1e-06 
0.0 -0.8995 0 -2.0 1e-06 
0.0 -0.8994 0 -2.0 1e-06 
0.0 -0.8993 0 -2.0 1e-06 
0.0 -0.8992 0 -2.0 1e-06 
0.0 -0.8991 0 -2.0 1e-06 
0.0 -0.899 0 -2.0 1e-06 
0.0 -0.8989 0 -2.0 1e-06 
0.0 -0.8988 0 -2.0 1e-06 
0.0 -0.8987 0 -2.0 1e-06 
0.0 -0.8986 0 -2.0 1e-06 
0.0 -0.8985 0 -2.0 1e-06 
0.0 -0.8984 0 -2.0 1e-06 
0.0 -0.8983 0 -2.0 1e-06 
0.0 -0.8982 0 -2.0 1e-06 
0.0 -0.8981 0 -2.0 1e-06 
0.0 -0.898 0 -2.0 1e-06 
0.0 -0.8979 0 -2.0 1e-06 
0.0 -0.8978 0 -2.0 1e-06 
0.0 -0.8977 0 -2.0 1e-06 
0.0 -0.8976 0 -2.0 1e-06 
0.0 -0.8975 0 -2.0 1e-06 
0.0 -0.8974 0 -2.0 1e-06 
0.0 -0.8973 0 -2.0 1e-06 
0.0 -0.8972 0 -2.0 1e-06 
0.0 -0.8971 0 -2.0 1e-06 
0.0 -0.897 0 -2.0 1e-06 
0.0 -0.8969 0 -2.0 1e-06 
0.0 -0.8968 0 -2.0 1e-06 
0.0 -0.8967 0 -2.0 1e-06 
0.0 -0.8966 0 -2.0 1e-06 
0.0 -0.8965 0 -2.0 1e-06 
0.0 -0.8964 0 -2.0 1e-06 
0.0 -0.8963 0 -2.0 1e-06 
0.0 -0.8962 0 -2.0 1e-06 
0.0 -0.8961 0 -2.0 1e-06 
0.0 -0.896 0 -2.0 1e-06 
0.0 -0.8959 0 -2.0 1e-06 
0.0 -0.8958 0 -2.0 1e-06 
0.0 -0.8957 0 -2.0 1e-06 
0.0 -0.8956 0 -2.0 1e-06 
0.0 -0.8955 0 -2.0 1e-06 
0.0 -0.8954 0 -2.0 1e-06 
0.0 -0.8953 0 -2.0 1e-06 
0.0 -0.8952 0 -2.0 1e-06 
0.0 -0.8951 0 -2.0 1e-06 
0.0 -0.895 0 -2.0 1e-06 
0.0 -0.8949 0 -2.0 1e-06 
0.0 -0.8948 0 -2.0 1e-06 
0.0 -0.8947 0 -2.0 1e-06 
0.0 -0.8946 0 -2.0 1e-06 
0.0 -0.8945 0 -2.0 1e-06 
0.0 -0.8944 0 -2.0 1e-06 
0.0 -0.8943 0 -2.0 1e-06 
0.0 -0.8942 0 -2.0 1e-06 
0.0 -0.8941 0 -2.0 1e-06 
0.0 -0.894 0 -2.0 1e-06 
0.0 -0.8939 0 -2.0 1e-06 
0.0 -0.8938 0 -2.0 1e-06 
0.0 -0.8937 0 -2.0 1e-06 
0.0 -0.8936 0 -2.0 1e-06 
0.0 -0.8935 0 -2.0 1e-06 
0.0 -0.8934 0 -2.0 1e-06 
0.0 -0.8933 0 -2.0 1e-06 
0.0 -0.8932 0 -2.0 1e-06 
0.0 -0.8931 0 -2.0 1e-06 
0.0 -0.893 0 -2.0 1e-06 
0.0 -0.8929 0 -2.0 1e-06 
0.0 -0.8928 0 -2.0 1e-06 
0.0 -0.8927 0 -2.0 1e-06 
0.0 -0.8926 0 -2.0 1e-06 
0.0 -0.8925 0 -2.0 1e-06 
0.0 -0.8924 0 -2.0 1e-06 
0.0 -0.8923 0 -2.0 1e-06 
0.0 -0.8922 0 -2.0 1e-06 
0.0 -0.8921 0 -2.0 1e-06 
0.0 -0.892 0 -2.0 1e-06 
0.0 -0.8919 0 -2.0 1e-06 
0.0 -0.8918 0 -2.0 1e-06 
0.0 -0.8917 0 -2.0 1e-06 
0.0 -0.8916 0 -2.0 1e-06 
0.0 -0.8915 0 -2.0 1e-06 
0.0 -0.8914 0 -2.0 1e-06 
0.0 -0.8913 0 -2.0 1e-06 
0.0 -0.8912 0 -2.0 1e-06 
0.0 -0.8911 0 -2.0 1e-06 
0.0 -0.891 0 -2.0 1e-06 
0.0 -0.8909 0 -2.0 1e-06 
0.0 -0.8908 0 -2.0 1e-06 
0.0 -0.8907 0 -2.0 1e-06 
0.0 -0.8906 0 -2.0 1e-06 
0.0 -0.8905 0 -2.0 1e-06 
0.0 -0.8904 0 -2.0 1e-06 
0.0 -0.8903 0 -2.0 1e-06 
0.0 -0.8902 0 -2.0 1e-06 
0.0 -0.8901 0 -2.0 1e-06 
0.0 -0.89 0 -2.0 1e-06 
0.0 -0.8899 0 -2.0 1e-06 
0.0 -0.8898 0 -2.0 1e-06 
0.0 -0.8897 0 -2.0 1e-06 
0.0 -0.8896 0 -2.0 1e-06 
0.0 -0.8895 0 -2.0 1e-06 
0.0 -0.8894 0 -2.0 1e-06 
0.0 -0.8893 0 -2.0 1e-06 
0.0 -0.8892 0 -2.0 1e-06 
0.0 -0.8891 0 -2.0 1e-06 
0.0 -0.889 0 -2.0 1e-06 
0.0 -0.8889 0 -2.0 1e-06 
0.0 -0.8888 0 -2.0 1e-06 
0.0 -0.8887 0 -2.0 1e-06 
0.0 -0.8886 0 -2.0 1e-06 
0.0 -0.8885 0 -2.0 1e-06 
0.0 -0.8884 0 -2.0 1e-06 
0.0 -0.8883 0 -2.0 1e-06 
0.0 -0.8882 0 -2.0 1e-06 
0.0 -0.8881 0 -2.0 1e-06 
0.0 -0.888 0 -2.0 1e-06 
0.0 -0.8879 0 -2.0 1e-06 
0.0 -0.8878 0 -2.0 1e-06 
0.0 -0.8877 0 -2.0 1e-06 
0.0 -0.8876 0 -2.0 1e-06 
0.0 -0.8875 0 -2.0 1e-06 
0.0 -0.8874 0 -2.0 1e-06 
0.0 -0.8873 0 -2.0 1e-06 
0.0 -0.8872 0 -2.0 1e-06 
0.0 -0.8871 0 -2.0 1e-06 
0.0 -0.887 0 -2.0 1e-06 
0.0 -0.8869 0 -2.0 1e-06 
0.0 -0.8868 0 -2.0 1e-06 
0.0 -0.8867 0 -2.0 1e-06 
0.0 -0.8866 0 -2.0 1e-06 
0.0 -0.8865 0 -2.0 1e-06 
0.0 -0.8864 0 -2.0 1e-06 
0.0 -0.8863 0 -2.0 1e-06 
0.0 -0.8862 0 -2.0 1e-06 
0.0 -0.8861 0 -2.0 1e-06 
0.0 -0.886 0 -2.0 1e-06 
0.0 -0.8859 0 -2.0 1e-06 
0.0 -0.8858 0 -2.0 1e-06 
0.0 -0.8857 0 -2.0 1e-06 
0.0 -0.8856 0 -2.0 1e-06 
0.0 -0.8855 0 -2.0 1e-06 
0.0 -0.8854 0 -2.0 1e-06 
0.0 -0.8853 0 -2.0 1e-06 
0.0 -0.8852 0 -2.0 1e-06 
0.0 -0.8851 0 -2.0 1e-06 
0.0 -0.885 0 -2.0 1e-06 
0.0 -0.8849 0 -2.0 1e-06 
0.0 -0.8848 0 -2.0 1e-06 
0.0 -0.8847 0 -2.0 1e-06 
0.0 -0.8846 0 -2.0 1e-06 
0.0 -0.8845 0 -2.0 1e-06 
0.0 -0.8844 0 -2.0 1e-06 
0.0 -0.8843 0 -2.0 1e-06 
0.0 -0.8842 0 -2.0 1e-06 
0.0 -0.8841 0 -2.0 1e-06 
0.0 -0.884 0 -2.0 1e-06 
0.0 -0.8839 0 -2.0 1e-06 
0.0 -0.8838 0 -2.0 1e-06 
0.0 -0.8837 0 -2.0 1e-06 
0.0 -0.8836 0 -2.0 1e-06 
0.0 -0.8835 0 -2.0 1e-06 
0.0 -0.8834 0 -2.0 1e-06 
0.0 -0.8833 0 -2.0 1e-06 
0.0 -0.8832 0 -2.0 1e-06 
0.0 -0.8831 0 -2.0 1e-06 
0.0 -0.883 0 -2.0 1e-06 
0.0 -0.8829 0 -2.0 1e-06 
0.0 -0.8828 0 -2.0 1e-06 
0.0 -0.8827 0 -2.0 1e-06 
0.0 -0.8826 0 -2.0 1e-06 
0.0 -0.8825 0 -2.0 1e-06 
0.0 -0.8824 0 -2.0 1e-06 
0.0 -0.8823 0 -2.0 1e-06 
0.0 -0.8822 0 -2.0 1e-06 
0.0 -0.8821 0 -2.0 1e-06 
0.0 -0.882 0 -2.0 1e-06 
0.0 -0.8819 0 -2.0 1e-06 
0.0 -0.8818 0 -2.0 1e-06 
0.0 -0.8817 0 -2.0 1e-06 
0.0 -0.8816 0 -2.0 1e-06 
0.0 -0.8815 0 -2.0 1e-06 
0.0 -0.8814 0 -2.0 1e-06 
0.0 -0.8813 0 -2.0 1e-06 
0.0 -0.8812 0 -2.0 1e-06 
0.0 -0.8811 0 -2.0 1e-06 
0.0 -0.881 0 -2.0 1e-06 
0.0 -0.8809 0 -2.0 1e-06 
0.0 -0.8808 0 -2.0 1e-06 
0.0 -0.8807 0 -2.0 1e-06 
0.0 -0.8806 0 -2.0 1e-06 
0.0 -0.8805 0 -2.0 1e-06 
0.0 -0.8804 0 -2.0 1e-06 
0.0 -0.8803 0 -2.0 1e-06 
0.0 -0.8802 0 -2.0 1e-06 
0.0 -0.8801 0 -2.0 1e-06 
0.0 -0.88 0 -2.0 1e-06 
0.0 -0.8799 0 -2.0 1e-06 
0.0 -0.8798 0 -2.0 1e-06 
0.0 -0.8797 0 -2.0 1e-06 
0.0 -0.8796 0 -2.0 1e-06 
0.0 -0.8795 0 -2.0 1e-06 
0.0 -0.8794 0 -2.0 1e-06 
0.0 -0.8793 0 -2.0 1e-06 
0.0 -0.8792 0 -2.0 1e-06 
0.0 -0.8791 0 -2.0 1e-06 
0.0 -0.879 0 -2.0 1e-06 
0.0 -0.8789 0 -2.0 1e-06 
0.0 -0.8788 0 -2.0 1e-06 
0.0 -0.8787 0 -2.0 1e-06 
0.0 -0.8786 0 -2.0 1e-06 
0.0 -0.8785 0 -2.0 1e-06 
0.0 -0.8784 0 -2.0 1e-06 
0.0 -0.8783 0 -2.0 1e-06 
0.0 -0.8782 0 -2.0 1e-06 
0.0 -0.8781 0 -2.0 1e-06 
0.0 -0.878 0 -2.0 1e-06 
0.0 -0.8779 0 -2.0 1e-06 
0.0 -0.8778 0 -2.0 1e-06 
0.0 -0.8777 0 -2.0 1e-06 
0.0 -0.8776 0 -2.0 1e-06 
0.0 -0.8775 0 -2.0 1e-06 
0.0 -0.8774 0 -2.0 1e-06 
0.0 -0.8773 0 -2.0 1e-06 
0.0 -0.8772 0 -2.0 1e-06 
0.0 -0.8771 0 -2.0 1e-06 
0.0 -0.877 0 -2.0 1e-06 
0.0 -0.8769 0 -2.0 1e-06 
0.0 -0.8768 0 -2.0 1e-06 
0.0 -0.8767 0 -2.0 1e-06 
0.0 -0.8766 0 -2.0 1e-06 
0.0 -0.8765 0 -2.0 1e-06 
0.0 -0.8764 0 -2.0 1e-06 
0.0 -0.8763 0 -2.0 1e-06 
0.0 -0.8762 0 -2.0 1e-06 
0.0 -0.8761 0 -2.0 1e-06 
0.0 -0.876 0 -2.0 1e-06 
0.0 -0.8759 0 -2.0 1e-06 
0.0 -0.8758 0 -2.0 1e-06 
0.0 -0.8757 0 -2.0 1e-06 
0.0 -0.8756 0 -2.0 1e-06 
0.0 -0.8755 0 -2.0 1e-06 
0.0 -0.8754 0 -2.0 1e-06 
0.0 -0.8753 0 -2.0 1e-06 
0.0 -0.8752 0 -2.0 1e-06 
0.0 -0.8751 0 -2.0 1e-06 
0.0 -0.875 0 -2.0 1e-06 
0.0 -0.8749 0 -2.0 1e-06 
0.0 -0.8748 0 -2.0 1e-06 
0.0 -0.8747 0 -2.0 1e-06 
0.0 -0.8746 0 -2.0 1e-06 
0.0 -0.8745 0 -2.0 1e-06 
0.0 -0.8744 0 -2.0 1e-06 
0.0 -0.8743 0 -2.0 1e-06 
0.0 -0.8742 0 -2.0 1e-06 
0.0 -0.8741 0 -2.0 1e-06 
0.0 -0.874 0 -2.0 1e-06 
0.0 -0.8739 0 -2.0 1e-06 
0.0 -0.8738 0 -2.0 1e-06 
0.0 -0.8737 0 -2.0 1e-06 
0.0 -0.8736 0 -2.0 1e-06 
0.0 -0.8735 0 -2.0 1e-06 
0.0 -0.8734 0 -2.0 1e-06 
0.0 -0.8733 0 -2.0 1e-06 
0.0 -0.8732 0 -2.0 1e-06 
0.0 -0.8731 0 -2.0 1e-06 
0.0 -0.873 0 -2.0 1e-06 
0.0 -0.8729 0 -2.0 1e-06 
0.0 -0.8728 0 -2.0 1e-06 
0.0 -0.8727 0 -2.0 1e-06 
0.0 -0.8726 0 -2.0 1e-06 
0.0 -0.8725 0 -2.0 1e-06 
0.0 -0.8724 0 -2.0 1e-06 
0.0 -0.8723 0 -2.0 1e-06 
0.0 -0.8722 0 -2.0 1e-06 
0.0 -0.8721 0 -2.0 1e-06 
0.0 -0.872 0 -2.0 1e-06 
0.0 -0.8719 0 -2.0 1e-06 
0.0 -0.8718 0 -2.0 1e-06 
0.0 -0.8717 0 -2.0 1e-06 
0.0 -0.8716 0 -2.0 1e-06 
0.0 -0.8715 0 -2.0 1e-06 
0.0 -0.8714 0 -2.0 1e-06 
0.0 -0.8713 0 -2.0 1e-06 
0.0 -0.8712 0 -2.0 1e-06 
0.0 -0.8711 0 -2.0 1e-06 
0.0 -0.871 0 -2.0 1e-06 
0.0 -0.8709 0 -2.0 1e-06 
0.0 -0.8708 0 -2.0 1e-06 
0.0 -0.8707 0 -2.0 1e-06 
0.0 -0.8706 0 -2.0 1e-06 
0.0 -0.8705 0 -2.0 1e-06 
0.0 -0.8704 0 -2.0 1e-06 
0.0 -0.8703 0 -2.0 1e-06 
0.0 -0.8702 0 -2.0 1e-06 
0.0 -0.8701 0 -2.0 1e-06 
0.0 -0.87 0 -2.0 1e-06 
0.0 -0.8699 0 -2.0 1e-06 
0.0 -0.8698 0 -2.0 1e-06 
0.0 -0.8697 0 -2.0 1e-06 
0.0 -0.8696 0 -2.0 1e-06 
0.0 -0.8695 0 -2.0 1e-06 
0.0 -0.8694 0 -2.0 1e-06 
0.0 -0.8693 0 -2.0 1e-06 
0.0 -0.8692 0 -2.0 1e-06 
0.0 -0.8691 0 -2.0 1e-06 
0.0 -0.869 0 -2.0 1e-06 
0.0 -0.8689 0 -2.0 1e-06 
0.0 -0.8688 0 -2.0 1e-06 
0.0 -0.8687 0 -2.0 1e-06 
0.0 -0.8686 0 -2.0 1e-06 
0.0 -0.8685 0 -2.0 1e-06 
0.0 -0.8684 0 -2.0 1e-06 
0.0 -0.8683 0 -2.0 1e-06 
0.0 -0.8682 0 -2.0 1e-06 
0.0 -0.8681 0 -2.0 1e-06 
0.0 -0.868 0 -2.0 1e-06 
0.0 -0.8679 0 -2.0 1e-06 
0.0 -0.8678 0 -2.0 1e-06 
0.0 -0.8677 0 -2.0 1e-06 
0.0 -0.8676 0 -2.0 1e-06 
0.0 -0.8675 0 -2.0 1e-06 
0.0 -0.8674 0 -2.0 1e-06 
0.0 -0.8673 0 -2.0 1e-06 
0.0 -0.8672 0 -2.0 1e-06 
0.0 -0.8671 0 -2.0 1e-06 
0.0 -0.867 0 -2.0 1e-06 
0.0 -0.8669 0 -2.0 1e-06 
0.0 -0.8668 0 -2.0 1e-06 
0.0 -0.8667 0 -2.0 1e-06 
0.0 -0.8666 0 -2.0 1e-06 
0.0 -0.8665 0 -2.0 1e-06 
0.0 -0.8664 0 -2.0 1e-06 
0.0 -0.8663 0 -2.0 1e-06 
0.0 -0.8662 0 -2.0 1e-06 
0.0 -0.8661 0 -2.0 1e-06 
0.0 -0.866 0 -2.0 1e-06 
0.0 -0.8659 0 -2.0 1e-06 
0.0 -0.8658 0 -2.0 1e-06 
0.0 -0.8657 0 -2.0 1e-06 
0.0 -0.8656 0 -2.0 1e-06 
0.0 -0.8655 0 -2.0 1e-06 
0.0 -0.8654 0 -2.0 1e-06 
0.0 -0.8653 0 -2.0 1e-06 
0.0 -0.8652 0 -2.0 1e-06 
0.0 -0.8651 0 -2.0 1e-06 
0.0 -0.865 0 -2.0 1e-06 
0.0 -0.8649 0 -2.0 1e-06 
0.0 -0.8648 0 -2.0 1e-06 
0.0 -0.8647 0 -2.0 1e-06 
0.0 -0.8646 0 -2.0 1e-06 
0.0 -0.8645 0 -2.0 1e-06 
0.0 -0.8644 0 -2.0 1e-06 
0.0 -0.8643 0 -2.0 1e-06 
0.0 -0.8642 0 -2.0 1e-06 
0.0 -0.8641 0 -2.0 1e-06 
0.0 -0.864 0 -2.0 1e-06 
0.0 -0.8639 0 -2.0 1e-06 
0.0 -0.8638 0 -2.0 1e-06 
0.0 -0.8637 0 -2.0 1e-06 
0.0 -0.8636 0 -2.0 1e-06 
0.0 -0.8635 0 -2.0 1e-06 
0.0 -0.8634 0 -2.0 1e-06 
0.0 -0.8633 0 -2.0 1e-06 
0.0 -0.8632 0 -2.0 1e-06 
0.0 -0.8631 0 -2.0 1e-06 
0.0 -0.863 0 -2.0 1e-06 
0.0 -0.8629 0 -2.0 1e-06 
0.0 -0.8628 0 -2.0 1e-06 
0.0 -0.8627 0 -2.0 1e-06 
0.0 -0.8626 0 -2.0 1e-06 
0.0 -0.8625 0 -2.0 1e-06 
0.0 -0.8624 0 -2.0 1e-06 
0.0 -0.8623 0 -2.0 1e-06 
0.0 -0.8622 0 -2.0 1e-06 
0.0 -0.8621 0 -2.0 1e-06 
0.0 -0.862 0 -2.0 1e-06 
0.0 -0.8619 0 -2.0 1e-06 
0.0 -0.8618 0 -2.0 1e-06 
0.0 -0.8617 0 -2.0 1e-06 
0.0 -0.8616 0 -2.0 1e-06 
0.0 -0.8615 0 -2.0 1e-06 
0.0 -0.8614 0 -2.0 1e-06 
0.0 -0.8613 0 -2.0 1e-06 
0.0 -0.8612 0 -2.0 1e-06 
0.0 -0.8611 0 -2.0 1e-06 
0.0 -0.861 0 -2.0 1e-06 
0.0 -0.8609 0 -2.0 1e-06 
0.0 -0.8608 0 -2.0 1e-06 
0.0 -0.8607 0 -2.0 1e-06 
0.0 -0.8606 0 -2.0 1e-06 
0.0 -0.8605 0 -2.0 1e-06 
0.0 -0.8604 0 -2.0 1e-06 
0.0 -0.8603 0 -2.0 1e-06 
0.0 -0.8602 0 -2.0 1e-06 
0.0 -0.8601 0 -2.0 1e-06 
0.0 -0.86 0 -2.0 1e-06 
0.0 -0.8599 0 -2.0 1e-06 
0.0 -0.8598 0 -2.0 1e-06 
0.0 -0.8597 0 -2.0 1e-06 
0.0 -0.8596 0 -2.0 1e-06 
0.0 -0.8595 0 -2.0 1e-06 
0.0 -0.8594 0 -2.0 1e-06 
0.0 -0.8593 0 -2.0 1e-06 
0.0 -0.8592 0 -2.0 1e-06 
0.0 -0.8591 0 -2.0 1e-06 
0.0 -0.859 0 -2.0 1e-06 
0.0 -0.8589 0 -2.0 1e-06 
0.0 -0.8588 0 -2.0 1e-06 
0.0 -0.8587 0 -2.0 1e-06 
0.0 -0.8586 0 -2.0 1e-06 
0.0 -0.8585 0 -2.0 1e-06 
0.0 -0.8584 0 -2.0 1e-06 
0.0 -0.8583 0 -2.0 1e-06 
0.0 -0.8582 0 -2.0 1e-06 
0.0 -0.8581 0 -2.0 1e-06 
0.0 -0.858 0 -2.0 1e-06 
0.0 -0.8579 0 -2.0 1e-06 
0.0 -0.8578 0 -2.0 1e-06 
0.0 -0.8577 0 -2.0 1e-06 
0.0 -0.8576 0 -2.0 1e-06 
0.0 -0.8575 0 -2.0 1e-06 
0.0 -0.8574 0 -2.0 1e-06 
0.0 -0.8573 0 -2.0 1e-06 
0.0 -0.8572 0 -2.0 1e-06 
0.0 -0.8571 0 -2.0 1e-06 
0.0 -0.857 0 -2.0 1e-06 
0.0 -0.8569 0 -2.0 1e-06 
0.0 -0.8568 0 -2.0 1e-06 
0.0 -0.8567 0 -2.0 1e-06 
0.0 -0.8566 0 -2.0 1e-06 
0.0 -0.8565 0 -2.0 1e-06 
0.0 -0.8564 0 -2.0 1e-06 
0.0 -0.8563 0 -2.0 1e-06 
0.0 -0.8562 0 -2.0 1e-06 
0.0 -0.8561 0 -2.0 1e-06 
0.0 -0.856 0 -2.0 1e-06 
0.0 -0.8559 0 -2.0 1e-06 
0.0 -0.8558 0 -2.0 1e-06 
0.0 -0.8557 0 -2.0 1e-06 
0.0 -0.8556 0 -2.0 1e-06 
0.0 -0.8555 0 -2.0 1e-06 
0.0 -0.8554 0 -2.0 1e-06 
0.0 -0.8553 0 -2.0 1e-06 
0.0 -0.8552 0 -2.0 1e-06 
0.0 -0.8551 0 -2.0 1e-06 
0.0 -0.855 0 -2.0 1e-06 
0.0 -0.8549 0 -2.0 1e-06 
0.0 -0.8548 0 -2.0 1e-06 
0.0 -0.8547 0 -2.0 1e-06 
0.0 -0.8546 0 -2.0 1e-06 
0.0 -0.8545 0 -2.0 1e-06 
0.0 -0.8544 0 -2.0 1e-06 
0.0 -0.8543 0 -2.0 1e-06 
0.0 -0.8542 0 -2.0 1e-06 
0.0 -0.8541 0 -2.0 1e-06 
0.0 -0.854 0 -2.0 1e-06 
0.0 -0.8539 0 -2.0 1e-06 
0.0 -0.8538 0 -2.0 1e-06 
0.0 -0.8537 0 -2.0 1e-06 
0.0 -0.8536 0 -2.0 1e-06 
0.0 -0.8535 0 -2.0 1e-06 
0.0 -0.8534 0 -2.0 1e-06 
0.0 -0.8533 0 -2.0 1e-06 
0.0 -0.8532 0 -2.0 1e-06 
0.0 -0.8531 0 -2.0 1e-06 
0.0 -0.853 0 -2.0 1e-06 
0.0 -0.8529 0 -2.0 1e-06 
0.0 -0.8528 0 -2.0 1e-06 
0.0 -0.8527 0 -2.0 1e-06 
0.0 -0.8526 0 -2.0 1e-06 
0.0 -0.8525 0 -2.0 1e-06 
0.0 -0.8524 0 -2.0 1e-06 
0.0 -0.8523 0 -2.0 1e-06 
0.0 -0.8522 0 -2.0 1e-06 
0.0 -0.8521 0 -2.0 1e-06 
0.0 -0.852 0 -2.0 1e-06 
0.0 -0.8519 0 -2.0 1e-06 
0.0 -0.8518 0 -2.0 1e-06 
0.0 -0.8517 0 -2.0 1e-06 
0.0 -0.8516 0 -2.0 1e-06 
0.0 -0.8515 0 -2.0 1e-06 
0.0 -0.8514 0 -2.0 1e-06 
0.0 -0.8513 0 -2.0 1e-06 
0.0 -0.8512 0 -2.0 1e-06 
0.0 -0.8511 0 -2.0 1e-06 
0.0 -0.851 0 -2.0 1e-06 
0.0 -0.8509 0 -2.0 1e-06 
0.0 -0.8508 0 -2.0 1e-06 
0.0 -0.8507 0 -2.0 1e-06 
0.0 -0.8506 0 -2.0 1e-06 
0.0 -0.8505 0 -2.0 1e-06 
0.0 -0.8504 0 -2.0 1e-06 
0.0 -0.8503 0 -2.0 1e-06 
0.0 -0.8502 0 -2.0 1e-06 
0.0 -0.8501 0 -2.0 1e-06 
0.0 -0.85 0 -2.0 1e-06 
0.0 -0.8499 0 -2.0 1e-06 
0.0 -0.8498 0 -2.0 1e-06 
0.0 -0.8497 0 -2.0 1e-06 
0.0 -0.8496 0 -2.0 1e-06 
0.0 -0.8495 0 -2.0 1e-06 
0.0 -0.8494 0 -2.0 1e-06 
0.0 -0.8493 0 -2.0 1e-06 
0.0 -0.8492 0 -2.0 1e-06 
0.0 -0.8491 0 -2.0 1e-06 
0.0 -0.849 0 -2.0 1e-06 
0.0 -0.8489 0 -2.0 1e-06 
0.0 -0.8488 0 -2.0 1e-06 
0.0 -0.8487 0 -2.0 1e-06 
0.0 -0.8486 0 -2.0 1e-06 
0.0 -0.8485 0 -2.0 1e-06 
0.0 -0.8484 0 -2.0 1e-06 
0.0 -0.8483 0 -2.0 1e-06 
0.0 -0.8482 0 -2.0 1e-06 
0.0 -0.8481 0 -2.0 1e-06 
0.0 -0.848 0 -2.0 1e-06 
0.0 -0.8479 0 -2.0 1e-06 
0.0 -0.8478 0 -2.0 1e-06 
0.0 -0.8477 0 -2.0 1e-06 
0.0 -0.8476 0 -2.0 1e-06 
0.0 -0.8475 0 -2.0 1e-06 
0.0 -0.8474 0 -2.0 1e-06 
0.0 -0.8473 0 -2.0 1e-06 
0.0 -0.8472 0 -2.0 1e-06 
0.0 -0.8471 0 -2.0 1e-06 
0.0 -0.847 0 -2.0 1e-06 
0.0 -0.8469 0 -2.0 1e-06 
0.0 -0.8468 0 -2.0 1e-06 
0.0 -0.8467 0 -2.0 1e-06 
0.0 -0.8466 0 -2.0 1e-06 
0.0 -0.8465 0 -2.0 1e-06 
0.0 -0.8464 0 -2.0 1e-06 
0.0 -0.8463 0 -2.0 1e-06 
0.0 -0.8462 0 -2.0 1e-06 
0.0 -0.8461 0 -2.0 1e-06 
0.0 -0.846 0 -2.0 1e-06 
0.0 -0.8459 0 -2.0 1e-06 
0.0 -0.8458 0 -2.0 1e-06 
0.0 -0.8457 0 -2.0 1e-06 
0.0 -0.8456 0 -2.0 1e-06 
0.0 -0.8455 0 -2.0 1e-06 
0.0 -0.8454 0 -2.0 1e-06 
0.0 -0.8453 0 -2.0 1e-06 
0.0 -0.8452 0 -2.0 1e-06 
0.0 -0.8451 0 -2.0 1e-06 
0.0 -0.845 0 -2.0 1e-06 
0.0 -0.8449 0 -2.0 1e-06 
0.0 -0.8448 0 -2.0 1e-06 
0.0 -0.8447 0 -2.0 1e-06 
0.0 -0.8446 0 -2.0 1e-06 
0.0 -0.8445 0 -2.0 1e-06 
0.0 -0.8444 0 -2.0 1e-06 
0.0 -0.8443 0 -2.0 1e-06 
0.0 -0.8442 0 -2.0 1e-06 
0.0 -0.8441 0 -2.0 1e-06 
0.0 -0.844 0 -2.0 1e-06 
0.0 -0.8439 0 -2.0 1e-06 
0.0 -0.8438 0 -2.0 1e-06 
0.0 -0.8437 0 -2.0 1e-06 
0.0 -0.8436 0 -2.0 1e-06 
0.0 -0.8435 0 -2.0 1e-06 
0.0 -0.8434 0 -2.0 1e-06 
0.0 -0.8433 0 -2.0 1e-06 
0.0 -0.8432 0 -2.0 1e-06 
0.0 -0.8431 0 -2.0 1e-06 
0.0 -0.843 0 -2.0 1e-06 
0.0 -0.8429 0 -2.0 1e-06 
0.0 -0.8428 0 -2.0 1e-06 
0.0 -0.8427 0 -2.0 1e-06 
0.0 -0.8426 0 -2.0 1e-06 
0.0 -0.8425 0 -2.0 1e-06 
0.0 -0.8424 0 -2.0 1e-06 
0.0 -0.8423 0 -2.0 1e-06 
0.0 -0.8422 0 -2.0 1e-06 
0.0 -0.8421 0 -2.0 1e-06 
0.0 -0.842 0 -2.0 1e-06 
0.0 -0.8419 0 -2.0 1e-06 
0.0 -0.8418 0 -2.0 1e-06 
0.0 -0.8417 0 -2.0 1e-06 
0.0 -0.8416 0 -2.0 1e-06 
0.0 -0.8415 0 -2.0 1e-06 
0.0 -0.8414 0 -2.0 1e-06 
0.0 -0.8413 0 -2.0 1e-06 
0.0 -0.8412 0 -2.0 1e-06 
0.0 -0.8411 0 -2.0 1e-06 
0.0 -0.841 0 -2.0 1e-06 
0.0 -0.8409 0 -2.0 1e-06 
0.0 -0.8408 0 -2.0 1e-06 
0.0 -0.8407 0 -2.0 1e-06 
0.0 -0.8406 0 -2.0 1e-06 
0.0 -0.8405 0 -2.0 1e-06 
0.0 -0.8404 0 -2.0 1e-06 
0.0 -0.8403 0 -2.0 1e-06 
0.0 -0.8402 0 -2.0 1e-06 
0.0 -0.8401 0 -2.0 1e-06 
0.0 -0.84 0 -2.0 1e-06 
0.0 -0.8399 0 -2.0 1e-06 
0.0 -0.8398 0 -2.0 1e-06 
0.0 -0.8397 0 -2.0 1e-06 
0.0 -0.8396 0 -2.0 1e-06 
0.0 -0.8395 0 -2.0 1e-06 
0.0 -0.8394 0 -2.0 1e-06 
0.0 -0.8393 0 -2.0 1e-06 
0.0 -0.8392 0 -2.0 1e-06 
0.0 -0.8391 0 -2.0 1e-06 
0.0 -0.839 0 -2.0 1e-06 
0.0 -0.8389 0 -2.0 1e-06 
0.0 -0.8388 0 -2.0 1e-06 
0.0 -0.8387 0 -2.0 1e-06 
0.0 -0.8386 0 -2.0 1e-06 
0.0 -0.8385 0 -2.0 1e-06 
0.0 -0.8384 0 -2.0 1e-06 
0.0 -0.8383 0 -2.0 1e-06 
0.0 -0.8382 0 -2.0 1e-06 
0.0 -0.8381 0 -2.0 1e-06 
0.0 -0.838 0 -2.0 1e-06 
0.0 -0.8379 0 -2.0 1e-06 
0.0 -0.8378 0 -2.0 1e-06 
0.0 -0.8377 0 -2.0 1e-06 
0.0 -0.8376 0 -2.0 1e-06 
0.0 -0.8375 0 -2.0 1e-06 
0.0 -0.8374 0 -2.0 1e-06 
0.0 -0.8373 0 -2.0 1e-06 
0.0 -0.8372 0 -2.0 1e-06 
0.0 -0.8371 0 -2.0 1e-06 
0.0 -0.837 0 -2.0 1e-06 
0.0 -0.8369 0 -2.0 1e-06 
0.0 -0.8368 0 -2.0 1e-06 
0.0 -0.8367 0 -2.0 1e-06 
0.0 -0.8366 0 -2.0 1e-06 
0.0 -0.8365 0 -2.0 1e-06 
0.0 -0.8364 0 -2.0 1e-06 
0.0 -0.8363 0 -2.0 1e-06 
0.0 -0.8362 0 -2.0 1e-06 
0.0 -0.8361 0 -2.0 1e-06 
0.0 -0.836 0 -2.0 1e-06 
0.0 -0.8359 0 -2.0 1e-06 
0.0 -0.8358 0 -2.0 1e-06 
0.0 -0.8357 0 -2.0 1e-06 
0.0 -0.8356 0 -2.0 1e-06 
0.0 -0.8355 0 -2.0 1e-06 
0.0 -0.8354 0 -2.0 1e-06 
0.0 -0.8353 0 -2.0 1e-06 
0.0 -0.8352 0 -2.0 1e-06 
0.0 -0.8351 0 -2.0 1e-06 
0.0 -0.835 0 -2.0 1e-06 
0.0 -0.8349 0 -2.0 1e-06 
0.0 -0.8348 0 -2.0 1e-06 
0.0 -0.8347 0 -2.0 1e-06 
0.0 -0.8346 0 -2.0 1e-06 
0.0 -0.8345 0 -2.0 1e-06 
0.0 -0.8344 0 -2.0 1e-06 
0.0 -0.8343 0 -2.0 1e-06 
0.0 -0.8342 0 -2.0 1e-06 
0.0 -0.8341 0 -2.0 1e-06 
0.0 -0.834 0 -2.0 1e-06 
0.0 -0.8339 0 -2.0 1e-06 
0.0 -0.8338 0 -2.0 1e-06 
0.0 -0.8337 0 -2.0 1e-06 
0.0 -0.8336 0 -2.0 1e-06 
0.0 -0.8335 0 -2.0 1e-06 
0.0 -0.8334 0 -2.0 1e-06 
0.0 -0.8333 0 -2.0 1e-06 
0.0 -0.8332 0 -2.0 1e-06 
0.0 -0.8331 0 -2.0 1e-06 
0.0 -0.833 0 -2.0 1e-06 
0.0 -0.8329 0 -2.0 1e-06 
0.0 -0.8328 0 -2.0 1e-06 
0.0 -0.8327 0 -2.0 1e-06 
0.0 -0.8326 0 -2.0 1e-06 
0.0 -0.8325 0 -2.0 1e-06 
0.0 -0.8324 0 -2.0 1e-06 
0.0 -0.8323 0 -2.0 1e-06 
0.0 -0.8322 0 -2.0 1e-06 
0.0 -0.8321 0 -2.0 1e-06 
0.0 -0.832 0 -2.0 1e-06 
0.0 -0.8319 0 -2.0 1e-06 
0.0 -0.8318 0 -2.0 1e-06 
0.0 -0.8317 0 -2.0 1e-06 
0.0 -0.8316 0 -2.0 1e-06 
0.0 -0.8315 0 -2.0 1e-06 
0.0 -0.8314 0 -2.0 1e-06 
0.0 -0.8313 0 -2.0 1e-06 
0.0 -0.8312 0 -2.0 1e-06 
0.0 -0.8311 0 -2.0 1e-06 
0.0 -0.831 0 -2.0 1e-06 
0.0 -0.8309 0 -2.0 1e-06 
0.0 -0.8308 0 -2.0 1e-06 
0.0 -0.8307 0 -2.0 1e-06 
0.0 -0.8306 0 -2.0 1e-06 
0.0 -0.8305 0 -2.0 1e-06 
0.0 -0.8304 0 -2.0 1e-06 
0.0 -0.8303 0 -2.0 1e-06 
0.0 -0.8302 0 -2.0 1e-06 
0.0 -0.8301 0 -2.0 1e-06 
0.0 -0.83 0 -2.0 1e-06 
0.0 -0.8299 0 -2.0 1e-06 
0.0 -0.8298 0 -2.0 1e-06 
0.0 -0.8297 0 -2.0 1e-06 
0.0 -0.8296 0 -2.0 1e-06 
0.0 -0.8295 0 -2.0 1e-06 
0.0 -0.8294 0 -2.0 1e-06 
0.0 -0.8293 0 -2.0 1e-06 
0.0 -0.8292 0 -2.0 1e-06 
0.0 -0.8291 0 -2.0 1e-06 
0.0 -0.829 0 -2.0 1e-06 
0.0 -0.8289 0 -2.0 1e-06 
0.0 -0.8288 0 -2.0 1e-06 
0.0 -0.8287 0 -2.0 1e-06 
0.0 -0.8286 0 -2.0 1e-06 
0.0 -0.8285 0 -2.0 1e-06 
0.0 -0.8284 0 -2.0 1e-06 
0.0 -0.8283 0 -2.0 1e-06 
0.0 -0.8282 0 -2.0 1e-06 
0.0 -0.8281 0 -2.0 1e-06 
0.0 -0.828 0 -2.0 1e-06 
0.0 -0.8279 0 -2.0 1e-06 
0.0 -0.8278 0 -2.0 1e-06 
0.0 -0.8277 0 -2.0 1e-06 
0.0 -0.8276 0 -2.0 1e-06 
0.0 -0.8275 0 -2.0 1e-06 
0.0 -0.8274 0 -2.0 1e-06 
0.0 -0.8273 0 -2.0 1e-06 
0.0 -0.8272 0 -2.0 1e-06 
0.0 -0.8271 0 -2.0 1e-06 
0.0 -0.827 0 -2.0 1e-06 
0.0 -0.8269 0 -2.0 1e-06 
0.0 -0.8268 0 -2.0 1e-06 
0.0 -0.8267 0 -2.0 1e-06 
0.0 -0.8266 0 -2.0 1e-06 
0.0 -0.8265 0 -2.0 1e-06 
0.0 -0.8264 0 -2.0 1e-06 
0.0 -0.8263 0 -2.0 1e-06 
0.0 -0.8262 0 -2.0 1e-06 
0.0 -0.8261 0 -2.0 1e-06 
0.0 -0.826 0 -2.0 1e-06 
0.0 -0.8259 0 -2.0 1e-06 
0.0 -0.8258 0 -2.0 1e-06 
0.0 -0.8257 0 -2.0 1e-06 
0.0 -0.8256 0 -2.0 1e-06 
0.0 -0.8255 0 -2.0 1e-06 
0.0 -0.8254 0 -2.0 1e-06 
0.0 -0.8253 0 -2.0 1e-06 
0.0 -0.8252 0 -2.0 1e-06 
0.0 -0.8251 0 -2.0 1e-06 
0.0 -0.825 0 -2.0 1e-06 
0.0 -0.8249 0 -2.0 1e-06 
0.0 -0.8248 0 -2.0 1e-06 
0.0 -0.8247 0 -2.0 1e-06 
0.0 -0.8246 0 -2.0 1e-06 
0.0 -0.8245 0 -2.0 1e-06 
0.0 -0.8244 0 -2.0 1e-06 
0.0 -0.8243 0 -2.0 1e-06 
0.0 -0.8242 0 -2.0 1e-06 
0.0 -0.8241 0 -2.0 1e-06 
0.0 -0.824 0 -2.0 1e-06 
0.0 -0.8239 0 -2.0 1e-06 
0.0 -0.8238 0 -2.0 1e-06 
0.0 -0.8237 0 -2.0 1e-06 
0.0 -0.8236 0 -2.0 1e-06 
0.0 -0.8235 0 -2.0 1e-06 
0.0 -0.8234 0 -2.0 1e-06 
0.0 -0.8233 0 -2.0 1e-06 
0.0 -0.8232 0 -2.0 1e-06 
0.0 -0.8231 0 -2.0 1e-06 
0.0 -0.823 0 -2.0 1e-06 
0.0 -0.8229 0 -2.0 1e-06 
0.0 -0.8228 0 -2.0 1e-06 
0.0 -0.8227 0 -2.0 1e-06 
0.0 -0.8226 0 -2.0 1e-06 
0.0 -0.8225 0 -2.0 1e-06 
0.0 -0.8224 0 -2.0 1e-06 
0.0 -0.8223 0 -2.0 1e-06 
0.0 -0.8222 0 -2.0 1e-06 
0.0 -0.8221 0 -2.0 1e-06 
0.0 -0.822 0 -2.0 1e-06 
0.0 -0.8219 0 -2.0 1e-06 
0.0 -0.8218 0 -2.0 1e-06 
0.0 -0.8217 0 -2.0 1e-06 
0.0 -0.8216 0 -2.0 1e-06 
0.0 -0.8215 0 -2.0 1e-06 
0.0 -0.8214 0 -2.0 1e-06 
0.0 -0.8213 0 -2.0 1e-06 
0.0 -0.8212 0 -2.0 1e-06 
0.0 -0.8211 0 -2.0 1e-06 
0.0 -0.821 0 -2.0 1e-06 
0.0 -0.8209 0 -2.0 1e-06 
0.0 -0.8208 0 -2.0 1e-06 
0.0 -0.8207 0 -2.0 1e-06 
0.0 -0.8206 0 -2.0 1e-06 
0.0 -0.8205 0 -2.0 1e-06 
0.0 -0.8204 0 -2.0 1e-06 
0.0 -0.8203 0 -2.0 1e-06 
0.0 -0.8202 0 -2.0 1e-06 
0.0 -0.8201 0 -2.0 1e-06 
0.0 -0.82 0 -2.0 1e-06 
0.0 -0.8199 0 -2.0 1e-06 
0.0 -0.8198 0 -2.0 1e-06 
0.0 -0.8197 0 -2.0 1e-06 
0.0 -0.8196 0 -2.0 1e-06 
0.0 -0.8195 0 -2.0 1e-06 
0.0 -0.8194 0 -2.0 1e-06 
0.0 -0.8193 0 -2.0 1e-06 
0.0 -0.8192 0 -2.0 1e-06 
0.0 -0.8191 0 -2.0 1e-06 
0.0 -0.819 0 -2.0 1e-06 
0.0 -0.8189 0 -2.0 1e-06 
0.0 -0.8188 0 -2.0 1e-06 
0.0 -0.8187 0 -2.0 1e-06 
0.0 -0.8186 0 -2.0 1e-06 
0.0 -0.8185 0 -2.0 1e-06 
0.0 -0.8184 0 -2.0 1e-06 
0.0 -0.8183 0 -2.0 1e-06 
0.0 -0.8182 0 -2.0 1e-06 
0.0 -0.8181 0 -2.0 1e-06 
0.0 -0.818 0 -2.0 1e-06 
0.0 -0.8179 0 -2.0 1e-06 
0.0 -0.8178 0 -2.0 1e-06 
0.0 -0.8177 0 -2.0 1e-06 
0.0 -0.8176 0 -2.0 1e-06 
0.0 -0.8175 0 -2.0 1e-06 
0.0 -0.8174 0 -2.0 1e-06 
0.0 -0.8173 0 -2.0 1e-06 
0.0 -0.8172 0 -2.0 1e-06 
0.0 -0.8171 0 -2.0 1e-06 
0.0 -0.817 0 -2.0 1e-06 
0.0 -0.8169 0 -2.0 1e-06 
0.0 -0.8168 0 -2.0 1e-06 
0.0 -0.8167 0 -2.0 1e-06 
0.0 -0.8166 0 -2.0 1e-06 
0.0 -0.8165 0 -2.0 1e-06 
0.0 -0.8164 0 -2.0 1e-06 
0.0 -0.8163 0 -2.0 1e-06 
0.0 -0.8162 0 -2.0 1e-06 
0.0 -0.8161 0 -2.0 1e-06 
0.0 -0.816 0 -2.0 1e-06 
0.0 -0.8159 0 -2.0 1e-06 
0.0 -0.8158 0 -2.0 1e-06 
0.0 -0.8157 0 -2.0 1e-06 
0.0 -0.8156 0 -2.0 1e-06 
0.0 -0.8155 0 -2.0 1e-06 
0.0 -0.8154 0 -2.0 1e-06 
0.0 -0.8153 0 -2.0 1e-06 
0.0 -0.8152 0 -2.0 1e-06 
0.0 -0.8151 0 -2.0 1e-06 
0.0 -0.815 0 -2.0 1e-06 
0.0 -0.8149 0 -2.0 1e-06 
0.0 -0.8148 0 -2.0 1e-06 
0.0 -0.8147 0 -2.0 1e-06 
0.0 -0.8146 0 -2.0 1e-06 
0.0 -0.8145 0 -2.0 1e-06 
0.0 -0.8144 0 -2.0 1e-06 
0.0 -0.8143 0 -2.0 1e-06 
0.0 -0.8142 0 -2.0 1e-06 
0.0 -0.8141 0 -2.0 1e-06 
0.0 -0.814 0 -2.0 1e-06 
0.0 -0.8139 0 -2.0 1e-06 
0.0 -0.8138 0 -2.0 1e-06 
0.0 -0.8137 0 -2.0 1e-06 
0.0 -0.8136 0 -2.0 1e-06 
0.0 -0.8135 0 -2.0 1e-06 
0.0 -0.8134 0 -2.0 1e-06 
0.0 -0.8133 0 -2.0 1e-06 
0.0 -0.8132 0 -2.0 1e-06 
0.0 -0.8131 0 -2.0 1e-06 
0.0 -0.813 0 -2.0 1e-06 
0.0 -0.8129 0 -2.0 1e-06 
0.0 -0.8128 0 -2.0 1e-06 
0.0 -0.8127 0 -2.0 1e-06 
0.0 -0.8126 0 -2.0 1e-06 
0.0 -0.8125 0 -2.0 1e-06 
0.0 -0.8124 0 -2.0 1e-06 
0.0 -0.8123 0 -2.0 1e-06 
0.0 -0.8122 0 -2.0 1e-06 
0.0 -0.8121 0 -2.0 1e-06 
0.0 -0.812 0 -2.0 1e-06 
0.0 -0.8119 0 -2.0 1e-06 
0.0 -0.8118 0 -2.0 1e-06 
0.0 -0.8117 0 -2.0 1e-06 
0.0 -0.8116 0 -2.0 1e-06 
0.0 -0.8115 0 -2.0 1e-06 
0.0 -0.8114 0 -2.0 1e-06 
0.0 -0.8113 0 -2.0 1e-06 
0.0 -0.8112 0 -2.0 1e-06 
0.0 -0.8111 0 -2.0 1e-06 
0.0 -0.811 0 -2.0 1e-06 
0.0 -0.8109 0 -2.0 1e-06 
0.0 -0.8108 0 -2.0 1e-06 
0.0 -0.8107 0 -2.0 1e-06 
0.0 -0.8106 0 -2.0 1e-06 
0.0 -0.8105 0 -2.0 1e-06 
0.0 -0.8104 0 -2.0 1e-06 
0.0 -0.8103 0 -2.0 1e-06 
0.0 -0.8102 0 -2.0 1e-06 
0.0 -0.8101 0 -2.0 1e-06 
0.0 -0.81 0 -2.0 1e-06 
0.0 -0.8099 0 -2.0 1e-06 
0.0 -0.8098 0 -2.0 1e-06 
0.0 -0.8097 0 -2.0 1e-06 
0.0 -0.8096 0 -2.0 1e-06 
0.0 -0.8095 0 -2.0 1e-06 
0.0 -0.8094 0 -2.0 1e-06 
0.0 -0.8093 0 -2.0 1e-06 
0.0 -0.8092 0 -2.0 1e-06 
0.0 -0.8091 0 -2.0 1e-06 
0.0 -0.809 0 -2.0 1e-06 
0.0 -0.8089 0 -2.0 1e-06 
0.0 -0.8088 0 -2.0 1e-06 
0.0 -0.8087 0 -2.0 1e-06 
0.0 -0.8086 0 -2.0 1e-06 
0.0 -0.8085 0 -2.0 1e-06 
0.0 -0.8084 0 -2.0 1e-06 
0.0 -0.8083 0 -2.0 1e-06 
0.0 -0.8082 0 -2.0 1e-06 
0.0 -0.8081 0 -2.0 1e-06 
0.0 -0.808 0 -2.0 1e-06 
0.0 -0.8079 0 -2.0 1e-06 
0.0 -0.8078 0 -2.0 1e-06 
0.0 -0.8077 0 -2.0 1e-06 
0.0 -0.8076 0 -2.0 1e-06 
0.0 -0.8075 0 -2.0 1e-06 
0.0 -0.8074 0 -2.0 1e-06 
0.0 -0.8073 0 -2.0 1e-06 
0.0 -0.8072 0 -2.0 1e-06 
0.0 -0.8071 0 -2.0 1e-06 
0.0 -0.807 0 -2.0 1e-06 
0.0 -0.8069 0 -2.0 1e-06 
0.0 -0.8068 0 -2.0 1e-06 
0.0 -0.8067 0 -2.0 1e-06 
0.0 -0.8066 0 -2.0 1e-06 
0.0 -0.8065 0 -2.0 1e-06 
0.0 -0.8064 0 -2.0 1e-06 
0.0 -0.8063 0 -2.0 1e-06 
0.0 -0.8062 0 -2.0 1e-06 
0.0 -0.8061 0 -2.0 1e-06 
0.0 -0.806 0 -2.0 1e-06 
0.0 -0.8059 0 -2.0 1e-06 
0.0 -0.8058 0 -2.0 1e-06 
0.0 -0.8057 0 -2.0 1e-06 
0.0 -0.8056 0 -2.0 1e-06 
0.0 -0.8055 0 -2.0 1e-06 
0.0 -0.8054 0 -2.0 1e-06 
0.0 -0.8053 0 -2.0 1e-06 
0.0 -0.8052 0 -2.0 1e-06 
0.0 -0.8051 0 -2.0 1e-06 
0.0 -0.805 0 -2.0 1e-06 
0.0 -0.8049 0 -2.0 1e-06 
0.0 -0.8048 0 -2.0 1e-06 
0.0 -0.8047 0 -2.0 1e-06 
0.0 -0.8046 0 -2.0 1e-06 
0.0 -0.8045 0 -2.0 1e-06 
0.0 -0.8044 0 -2.0 1e-06 
0.0 -0.8043 0 -2.0 1e-06 
0.0 -0.8042 0 -2.0 1e-06 
0.0 -0.8041 0 -2.0 1e-06 
0.0 -0.804 0 -2.0 1e-06 
0.0 -0.8039 0 -2.0 1e-06 
0.0 -0.8038 0 -2.0 1e-06 
0.0 -0.8037 0 -2.0 1e-06 
0.0 -0.8036 0 -2.0 1e-06 
0.0 -0.8035 0 -2.0 1e-06 
0.0 -0.8034 0 -2.0 1e-06 
0.0 -0.8033 0 -2.0 1e-06 
0.0 -0.8032 0 -2.0 1e-06 
0.0 -0.8031 0 -2.0 1e-06 
0.0 -0.803 0 -2.0 1e-06 
0.0 -0.8029 0 -2.0 1e-06 
0.0 -0.8028 0 -2.0 1e-06 
0.0 -0.8027 0 -2.0 1e-06 
0.0 -0.8026 0 -2.0 1e-06 
0.0 -0.8025 0 -2.0 1e-06 
0.0 -0.8024 0 -2.0 1e-06 
0.0 -0.8023 0 -2.0 1e-06 
0.0 -0.8022 0 -2.0 1e-06 
0.0 -0.8021 0 -2.0 1e-06 
0.0 -0.802 0 -2.0 1e-06 
0.0 -0.8019 0 -2.0 1e-06 
0.0 -0.8018 0 -2.0 1e-06 
0.0 -0.8017 0 -2.0 1e-06 
0.0 -0.8016 0 -2.0 1e-06 
0.0 -0.8015 0 -2.0 1e-06 
0.0 -0.8014 0 -2.0 1e-06 
0.0 -0.8013 0 -2.0 1e-06 
0.0 -0.8012 0 -2.0 1e-06 
0.0 -0.8011 0 -2.0 1e-06 
0.0 -0.801 0 -2.0 1e-06 
0.0 -0.8009 0 -2.0 1e-06 
0.0 -0.8008 0 -2.0 1e-06 
0.0 -0.8007 0 -2.0 1e-06 
0.0 -0.8006 0 -2.0 1e-06 
0.0 -0.8005 0 -2.0 1e-06 
0.0 -0.8004 0 -2.0 1e-06 
0.0 -0.8003 0 -2.0 1e-06 
0.0 -0.8002 0 -2.0 1e-06 
0.0 -0.8001 0 -2.0 1e-06 
0.0 -0.8 0 -2.0 1e-06 
0.0 -0.7999 0 -2.0 1e-06 
0.0 -0.7998 0 -2.0 1e-06 
0.0 -0.7997 0 -2.0 1e-06 
0.0 -0.7996 0 -2.0 1e-06 
0.0 -0.7995 0 -2.0 1e-06 
0.0 -0.7994 0 -2.0 1e-06 
0.0 -0.7993 0 -2.0 1e-06 
0.0 -0.7992 0 -2.0 1e-06 
0.0 -0.7991 0 -2.0 1e-06 
0.0 -0.799 0 -2.0 1e-06 
0.0 -0.7989 0 -2.0 1e-06 
0.0 -0.7988 0 -2.0 1e-06 
0.0 -0.7987 0 -2.0 1e-06 
0.0 -0.7986 0 -2.0 1e-06 
0.0 -0.7985 0 -2.0 1e-06 
0.0 -0.7984 0 -2.0 1e-06 
0.0 -0.7983 0 -2.0 1e-06 
0.0 -0.7982 0 -2.0 1e-06 
0.0 -0.7981 0 -2.0 1e-06 
0.0 -0.798 0 -2.0 1e-06 
0.0 -0.7979 0 -2.0 1e-06 
0.0 -0.7978 0 -2.0 1e-06 
0.0 -0.7977 0 -2.0 1e-06 
0.0 -0.7976 0 -2.0 1e-06 
0.0 -0.7975 0 -2.0 1e-06 
0.0 -0.7974 0 -2.0 1e-06 
0.0 -0.7973 0 -2.0 1e-06 
0.0 -0.7972 0 -2.0 1e-06 
0.0 -0.7971 0 -2.0 1e-06 
0.0 -0.797 0 -2.0 1e-06 
0.0 -0.7969 0 -2.0 1e-06 
0.0 -0.7968 0 -2.0 1e-06 
0.0 -0.7967 0 -2.0 1e-06 
0.0 -0.7966 0 -2.0 1e-06 
0.0 -0.7965 0 -2.0 1e-06 
0.0 -0.7964 0 -2.0 1e-06 
0.0 -0.7963 0 -2.0 1e-06 
0.0 -0.7962 0 -2.0 1e-06 
0.0 -0.7961 0 -2.0 1e-06 
0.0 -0.796 0 -2.0 1e-06 
0.0 -0.7959 0 -2.0 1e-06 
0.0 -0.7958 0 -2.0 1e-06 
0.0 -0.7957 0 -2.0 1e-06 
0.0 -0.7956 0 -2.0 1e-06 
0.0 -0.7955 0 -2.0 1e-06 
0.0 -0.7954 0 -2.0 1e-06 
0.0 -0.7953 0 -2.0 1e-06 
0.0 -0.7952 0 -2.0 1e-06 
0.0 -0.7951 0 -2.0 1e-06 
0.0 -0.795 0 -2.0 1e-06 
0.0 -0.7949 0 -2.0 1e-06 
0.0 -0.7948 0 -2.0 1e-06 
0.0 -0.7947 0 -2.0 1e-06 
0.0 -0.7946 0 -2.0 1e-06 
0.0 -0.7945 0 -2.0 1e-06 
0.0 -0.7944 0 -2.0 1e-06 
0.0 -0.7943 0 -2.0 1e-06 
0.0 -0.7942 0 -2.0 1e-06 
0.0 -0.7941 0 -2.0 1e-06 
0.0 -0.794 0 -2.0 1e-06 
0.0 -0.7939 0 -2.0 1e-06 
0.0 -0.7938 0 -2.0 1e-06 
0.0 -0.7937 0 -2.0 1e-06 
0.0 -0.7936 0 -2.0 1e-06 
0.0 -0.7935 0 -2.0 1e-06 
0.0 -0.7934 0 -2.0 1e-06 
0.0 -0.7933 0 -2.0 1e-06 
0.0 -0.7932 0 -2.0 1e-06 
0.0 -0.7931 0 -2.0 1e-06 
0.0 -0.793 0 -2.0 1e-06 
0.0 -0.7929 0 -2.0 1e-06 
0.0 -0.7928 0 -2.0 1e-06 
0.0 -0.7927 0 -2.0 1e-06 
0.0 -0.7926 0 -2.0 1e-06 
0.0 -0.7925 0 -2.0 1e-06 
0.0 -0.7924 0 -2.0 1e-06 
0.0 -0.7923 0 -2.0 1e-06 
0.0 -0.7922 0 -2.0 1e-06 
0.0 -0.7921 0 -2.0 1e-06 
0.0 -0.792 0 -2.0 1e-06 
0.0 -0.7919 0 -2.0 1e-06 
0.0 -0.7918 0 -2.0 1e-06 
0.0 -0.7917 0 -2.0 1e-06 
0.0 -0.7916 0 -2.0 1e-06 
0.0 -0.7915 0 -2.0 1e-06 
0.0 -0.7914 0 -2.0 1e-06 
0.0 -0.7913 0 -2.0 1e-06 
0.0 -0.7912 0 -2.0 1e-06 
0.0 -0.7911 0 -2.0 1e-06 
0.0 -0.791 0 -2.0 1e-06 
0.0 -0.7909 0 -2.0 1e-06 
0.0 -0.7908 0 -2.0 1e-06 
0.0 -0.7907 0 -2.0 1e-06 
0.0 -0.7906 0 -2.0 1e-06 
0.0 -0.7905 0 -2.0 1e-06 
0.0 -0.7904 0 -2.0 1e-06 
0.0 -0.7903 0 -2.0 1e-06 
0.0 -0.7902 0 -2.0 1e-06 
0.0 -0.7901 0 -2.0 1e-06 
0.0 -0.79 0 -2.0 1e-06 
0.0 -0.7899 0 -2.0 1e-06 
0.0 -0.7898 0 -2.0 1e-06 
0.0 -0.7897 0 -2.0 1e-06 
0.0 -0.7896 0 -2.0 1e-06 
0.0 -0.7895 0 -2.0 1e-06 
0.0 -0.7894 0 -2.0 1e-06 
0.0 -0.7893 0 -2.0 1e-06 
0.0 -0.7892 0 -2.0 1e-06 
0.0 -0.7891 0 -2.0 1e-06 
0.0 -0.789 0 -2.0 1e-06 
0.0 -0.7889 0 -2.0 1e-06 
0.0 -0.7888 0 -2.0 1e-06 
0.0 -0.7887 0 -2.0 1e-06 
0.0 -0.7886 0 -2.0 1e-06 
0.0 -0.7885 0 -2.0 1e-06 
0.0 -0.7884 0 -2.0 1e-06 
0.0 -0.7883 0 -2.0 1e-06 
0.0 -0.7882 0 -2.0 1e-06 
0.0 -0.7881 0 -2.0 1e-06 
0.0 -0.788 0 -2.0 1e-06 
0.0 -0.7879 0 -2.0 1e-06 
0.0 -0.7878 0 -2.0 1e-06 
0.0 -0.7877 0 -2.0 1e-06 
0.0 -0.7876 0 -2.0 1e-06 
0.0 -0.7875 0 -2.0 1e-06 
0.0 -0.7874 0 -2.0 1e-06 
0.0 -0.7873 0 -2.0 1e-06 
0.0 -0.7872 0 -2.0 1e-06 
0.0 -0.7871 0 -2.0 1e-06 
0.0 -0.787 0 -2.0 1e-06 
0.0 -0.7869 0 -2.0 1e-06 
0.0 -0.7868 0 -2.0 1e-06 
0.0 -0.7867 0 -2.0 1e-06 
0.0 -0.7866 0 -2.0 1e-06 
0.0 -0.7865 0 -2.0 1e-06 
0.0 -0.7864 0 -2.0 1e-06 
0.0 -0.7863 0 -2.0 1e-06 
0.0 -0.7862 0 -2.0 1e-06 
0.0 -0.7861 0 -2.0 1e-06 
0.0 -0.786 0 -2.0 1e-06 
0.0 -0.7859 0 -2.0 1e-06 
0.0 -0.7858 0 -2.0 1e-06 
0.0 -0.7857 0 -2.0 1e-06 
0.0 -0.7856 0 -2.0 1e-06 
0.0 -0.7855 0 -2.0 1e-06 
0.0 -0.7854 0 -2.0 1e-06 
0.0 -0.7853 0 -2.0 1e-06 
0.0 -0.7852 0 -2.0 1e-06 
0.0 -0.7851 0 -2.0 1e-06 
0.0 -0.785 0 -2.0 1e-06 
0.0 -0.7849 0 -2.0 1e-06 
0.0 -0.7848 0 -2.0 1e-06 
0.0 -0.7847 0 -2.0 1e-06 
0.0 -0.7846 0 -2.0 1e-06 
0.0 -0.7845 0 -2.0 1e-06 
0.0 -0.7844 0 -2.0 1e-06 
0.0 -0.7843 0 -2.0 1e-06 
0.0 -0.7842 0 -2.0 1e-06 
0.0 -0.7841 0 -2.0 1e-06 
0.0 -0.784 0 -2.0 1e-06 
0.0 -0.7839 0 -2.0 1e-06 
0.0 -0.7838 0 -2.0 1e-06 
0.0 -0.7837 0 -2.0 1e-06 
0.0 -0.7836 0 -2.0 1e-06 
0.0 -0.7835 0 -2.0 1e-06 
0.0 -0.7834 0 -2.0 1e-06 
0.0 -0.7833 0 -2.0 1e-06 
0.0 -0.7832 0 -2.0 1e-06 
0.0 -0.7831 0 -2.0 1e-06 
0.0 -0.783 0 -2.0 1e-06 
0.0 -0.7829 0 -2.0 1e-06 
0.0 -0.7828 0 -2.0 1e-06 
0.0 -0.7827 0 -2.0 1e-06 
0.0 -0.7826 0 -2.0 1e-06 
0.0 -0.7825 0 -2.0 1e-06 
0.0 -0.7824 0 -2.0 1e-06 
0.0 -0.7823 0 -2.0 1e-06 
0.0 -0.7822 0 -2.0 1e-06 
0.0 -0.7821 0 -2.0 1e-06 
0.0 -0.782 0 -2.0 1e-06 
0.0 -0.7819 0 -2.0 1e-06 
0.0 -0.7818 0 -2.0 1e-06 
0.0 -0.7817 0 -2.0 1e-06 
0.0 -0.7816 0 -2.0 1e-06 
0.0 -0.7815 0 -2.0 1e-06 
0.0 -0.7814 0 -2.0 1e-06 
0.0 -0.7813 0 -2.0 1e-06 
0.0 -0.7812 0 -2.0 1e-06 
0.0 -0.7811 0 -2.0 1e-06 
0.0 -0.781 0 -2.0 1e-06 
0.0 -0.7809 0 -2.0 1e-06 
0.0 -0.7808 0 -2.0 1e-06 
0.0 -0.7807 0 -2.0 1e-06 
0.0 -0.7806 0 -2.0 1e-06 
0.0 -0.7805 0 -2.0 1e-06 
0.0 -0.7804 0 -2.0 1e-06 
0.0 -0.7803 0 -2.0 1e-06 
0.0 -0.7802 0 -2.0 1e-06 
0.0 -0.7801 0 -2.0 1e-06 
0.0 -0.78 0 -2.0 1e-06 
0.0 -0.7799 0 -2.0 1e-06 
0.0 -0.7798 0 -2.0 1e-06 
0.0 -0.7797 0 -2.0 1e-06 
0.0 -0.7796 0 -2.0 1e-06 
0.0 -0.7795 0 -2.0 1e-06 
0.0 -0.7794 0 -2.0 1e-06 
0.0 -0.7793 0 -2.0 1e-06 
0.0 -0.7792 0 -2.0 1e-06 
0.0 -0.7791 0 -2.0 1e-06 
0.0 -0.779 0 -2.0 1e-06 
0.0 -0.7789 0 -2.0 1e-06 
0.0 -0.7788 0 -2.0 1e-06 
0.0 -0.7787 0 -2.0 1e-06 
0.0 -0.7786 0 -2.0 1e-06 
0.0 -0.7785 0 -2.0 1e-06 
0.0 -0.7784 0 -2.0 1e-06 
0.0 -0.7783 0 -2.0 1e-06 
0.0 -0.7782 0 -2.0 1e-06 
0.0 -0.7781 0 -2.0 1e-06 
0.0 -0.778 0 -2.0 1e-06 
0.0 -0.7779 0 -2.0 1e-06 
0.0 -0.7778 0 -2.0 1e-06 
0.0 -0.7777 0 -2.0 1e-06 
0.0 -0.7776 0 -2.0 1e-06 
0.0 -0.7775 0 -2.0 1e-06 
0.0 -0.7774 0 -2.0 1e-06 
0.0 -0.7773 0 -2.0 1e-06 
0.0 -0.7772 0 -2.0 1e-06 
0.0 -0.7771 0 -2.0 1e-06 
0.0 -0.777 0 -2.0 1e-06 
0.0 -0.7769 0 -2.0 1e-06 
0.0 -0.7768 0 -2.0 1e-06 
0.0 -0.7767 0 -2.0 1e-06 
0.0 -0.7766 0 -2.0 1e-06 
0.0 -0.7765 0 -2.0 1e-06 
0.0 -0.7764 0 -2.0 1e-06 
0.0 -0.7763 0 -2.0 1e-06 
0.0 -0.7762 0 -2.0 1e-06 
0.0 -0.7761 0 -2.0 1e-06 
0.0 -0.776 0 -2.0 1e-06 
0.0 -0.7759 0 -2.0 1e-06 
0.0 -0.7758 0 -2.0 1e-06 
0.0 -0.7757 0 -2.0 1e-06 
0.0 -0.7756 0 -2.0 1e-06 
0.0 -0.7755 0 -2.0 1e-06 
0.0 -0.7754 0 -2.0 1e-06 
0.0 -0.7753 0 -2.0 1e-06 
0.0 -0.7752 0 -2.0 1e-06 
0.0 -0.7751 0 -2.0 1e-06 
0.0 -0.775 0 -2.0 1e-06 
0.0 -0.7749 0 -2.0 1e-06 
0.0 -0.7748 0 -2.0 1e-06 
0.0 -0.7747 0 -2.0 1e-06 
0.0 -0.7746 0 -2.0 1e-06 
0.0 -0.7745 0 -2.0 1e-06 
0.0 -0.7744 0 -2.0 1e-06 
0.0 -0.7743 0 -2.0 1e-06 
0.0 -0.7742 0 -2.0 1e-06 
0.0 -0.7741 0 -2.0 1e-06 
0.0 -0.774 0 -2.0 1e-06 
0.0 -0.7739 0 -2.0 1e-06 
0.0 -0.7738 0 -2.0 1e-06 
0.0 -0.7737 0 -2.0 1e-06 
0.0 -0.7736 0 -2.0 1e-06 
0.0 -0.7735 0 -2.0 1e-06 
0.0 -0.7734 0 -2.0 1e-06 
0.0 -0.7733 0 -2.0 1e-06 
0.0 -0.7732 0 -2.0 1e-06 
0.0 -0.7731 0 -2.0 1e-06 
0.0 -0.773 0 -2.0 1e-06 
0.0 -0.7729 0 -2.0 1e-06 
0.0 -0.7728 0 -2.0 1e-06 
0.0 -0.7727 0 -2.0 1e-06 
0.0 -0.7726 0 -2.0 1e-06 
0.0 -0.7725 0 -2.0 1e-06 
0.0 -0.7724 0 -2.0 1e-06 
0.0 -0.7723 0 -2.0 1e-06 
0.0 -0.7722 0 -2.0 1e-06 
0.0 -0.7721 0 -2.0 1e-06 
0.0 -0.772 0 -2.0 1e-06 
0.0 -0.7719 0 -2.0 1e-06 
0.0 -0.7718 0 -2.0 1e-06 
0.0 -0.7717 0 -2.0 1e-06 
0.0 -0.7716 0 -2.0 1e-06 
0.0 -0.7715 0 -2.0 1e-06 
0.0 -0.7714 0 -2.0 1e-06 
0.0 -0.7713 0 -2.0 1e-06 
0.0 -0.7712 0 -2.0 1e-06 
0.0 -0.7711 0 -2.0 1e-06 
0.0 -0.771 0 -2.0 1e-06 
0.0 -0.7709 0 -2.0 1e-06 
0.0 -0.7708 0 -2.0 1e-06 
0.0 -0.7707 0 -2.0 1e-06 
0.0 -0.7706 0 -2.0 1e-06 
0.0 -0.7705 0 -2.0 1e-06 
0.0 -0.7704 0 -2.0 1e-06 
0.0 -0.7703 0 -2.0 1e-06 
0.0 -0.7702 0 -2.0 1e-06 
0.0 -0.7701 0 -2.0 1e-06 
0.0 -0.77 0 -2.0 1e-06 
0.0 -0.7699 0 -2.0 1e-06 
0.0 -0.7698 0 -2.0 1e-06 
0.0 -0.7697 0 -2.0 1e-06 
0.0 -0.7696 0 -2.0 1e-06 
0.0 -0.7695 0 -2.0 1e-06 
0.0 -0.7694 0 -2.0 1e-06 
0.0 -0.7693 0 -2.0 1e-06 
0.0 -0.7692 0 -2.0 1e-06 
0.0 -0.7691 0 -2.0 1e-06 
0.0 -0.769 0 -2.0 1e-06 
0.0 -0.7689 0 -2.0 1e-06 
0.0 -0.7688 0 -2.0 1e-06 
0.0 -0.7687 0 -2.0 1e-06 
0.0 -0.7686 0 -2.0 1e-06 
0.0 -0.7685 0 -2.0 1e-06 
0.0 -0.7684 0 -2.0 1e-06 
0.0 -0.7683 0 -2.0 1e-06 
0.0 -0.7682 0 -2.0 1e-06 
0.0 -0.7681 0 -2.0 1e-06 
0.0 -0.768 0 -2.0 1e-06 
0.0 -0.7679 0 -2.0 1e-06 
0.0 -0.7678 0 -2.0 1e-06 
0.0 -0.7677 0 -2.0 1e-06 
0.0 -0.7676 0 -2.0 1e-06 
0.0 -0.7675 0 -2.0 1e-06 
0.0 -0.7674 0 -2.0 1e-06 
0.0 -0.7673 0 -2.0 1e-06 
0.0 -0.7672 0 -2.0 1e-06 
0.0 -0.7671 0 -2.0 1e-06 
0.0 -0.767 0 -2.0 1e-06 
0.0 -0.7669 0 -2.0 1e-06 
0.0 -0.7668 0 -2.0 1e-06 
0.0 -0.7667 0 -2.0 1e-06 
0.0 -0.7666 0 -2.0 1e-06 
0.0 -0.7665 0 -2.0 1e-06 
0.0 -0.7664 0 -2.0 1e-06 
0.0 -0.7663 0 -2.0 1e-06 
0.0 -0.7662 0 -2.0 1e-06 
0.0 -0.7661 0 -2.0 1e-06 
0.0 -0.766 0 -2.0 1e-06 
0.0 -0.7659 0 -2.0 1e-06 
0.0 -0.7658 0 -2.0 1e-06 
0.0 -0.7657 0 -2.0 1e-06 
0.0 -0.7656 0 -2.0 1e-06 
0.0 -0.7655 0 -2.0 1e-06 
0.0 -0.7654 0 -2.0 1e-06 
0.0 -0.7653 0 -2.0 1e-06 
0.0 -0.7652 0 -2.0 1e-06 
0.0 -0.7651 0 -2.0 1e-06 
0.0 -0.765 0 -2.0 1e-06 
0.0 -0.7649 0 -2.0 1e-06 
0.0 -0.7648 0 -2.0 1e-06 
0.0 -0.7647 0 -2.0 1e-06 
0.0 -0.7646 0 -2.0 1e-06 
0.0 -0.7645 0 -2.0 1e-06 
0.0 -0.7644 0 -2.0 1e-06 
0.0 -0.7643 0 -2.0 1e-06 
0.0 -0.7642 0 -2.0 1e-06 
0.0 -0.7641 0 -2.0 1e-06 
0.0 -0.764 0 -2.0 1e-06 
0.0 -0.7639 0 -2.0 1e-06 
0.0 -0.7638 0 -2.0 1e-06 
0.0 -0.7637 0 -2.0 1e-06 
0.0 -0.7636 0 -2.0 1e-06 
0.0 -0.7635 0 -2.0 1e-06 
0.0 -0.7634 0 -2.0 1e-06 
0.0 -0.7633 0 -2.0 1e-06 
0.0 -0.7632 0 -2.0 1e-06 
0.0 -0.7631 0 -2.0 1e-06 
0.0 -0.763 0 -2.0 1e-06 
0.0 -0.7629 0 -2.0 1e-06 
0.0 -0.7628 0 -2.0 1e-06 
0.0 -0.7627 0 -2.0 1e-06 
0.0 -0.7626 0 -2.0 1e-06 
0.0 -0.7625 0 -2.0 1e-06 
0.0 -0.7624 0 -2.0 1e-06 
0.0 -0.7623 0 -2.0 1e-06 
0.0 -0.7622 0 -2.0 1e-06 
0.0 -0.7621 0 -2.0 1e-06 
0.0 -0.762 0 -2.0 1e-06 
0.0 -0.7619 0 -2.0 1e-06 
0.0 -0.7618 0 -2.0 1e-06 
0.0 -0.7617 0 -2.0 1e-06 
0.0 -0.7616 0 -2.0 1e-06 
0.0 -0.7615 0 -2.0 1e-06 
0.0 -0.7614 0 -2.0 1e-06 
0.0 -0.7613 0 -2.0 1e-06 
0.0 -0.7612 0 -2.0 1e-06 
0.0 -0.7611 0 -2.0 1e-06 
0.0 -0.761 0 -2.0 1e-06 
0.0 -0.7609 0 -2.0 1e-06 
0.0 -0.7608 0 -2.0 1e-06 
0.0 -0.7607 0 -2.0 1e-06 
0.0 -0.7606 0 -2.0 1e-06 
0.0 -0.7605 0 -2.0 1e-06 
0.0 -0.7604 0 -2.0 1e-06 
0.0 -0.7603 0 -2.0 1e-06 
0.0 -0.7602 0 -2.0 1e-06 
0.0 -0.7601 0 -2.0 1e-06 
0.0 -0.76 0 -2.0 1e-06 
0.0 -0.7599 0 -2.0 1e-06 
0.0 -0.7598 0 -2.0 1e-06 
0.0 -0.7597 0 -2.0 1e-06 
0.0 -0.7596 0 -2.0 1e-06 
0.0 -0.7595 0 -2.0 1e-06 
0.0 -0.7594 0 -2.0 1e-06 
0.0 -0.7593 0 -2.0 1e-06 
0.0 -0.7592 0 -2.0 1e-06 
0.0 -0.7591 0 -2.0 1e-06 
0.0 -0.759 0 -2.0 1e-06 
0.0 -0.7589 0 -2.0 1e-06 
0.0 -0.7588 0 -2.0 1e-06 
0.0 -0.7587 0 -2.0 1e-06 
0.0 -0.7586 0 -2.0 1e-06 
0.0 -0.7585 0 -2.0 1e-06 
0.0 -0.7584 0 -2.0 1e-06 
0.0 -0.7583 0 -2.0 1e-06 
0.0 -0.7582 0 -2.0 1e-06 
0.0 -0.7581 0 -2.0 1e-06 
0.0 -0.758 0 -2.0 1e-06 
0.0 -0.7579 0 -2.0 1e-06 
0.0 -0.7578 0 -2.0 1e-06 
0.0 -0.7577 0 -2.0 1e-06 
0.0 -0.7576 0 -2.0 1e-06 
0.0 -0.7575 0 -2.0 1e-06 
0.0 -0.7574 0 -2.0 1e-06 
0.0 -0.7573 0 -2.0 1e-06 
0.0 -0.7572 0 -2.0 1e-06 
0.0 -0.7571 0 -2.0 1e-06 
0.0 -0.757 0 -2.0 1e-06 
0.0 -0.7569 0 -2.0 1e-06 
0.0 -0.7568 0 -2.0 1e-06 
0.0 -0.7567 0 -2.0 1e-06 
0.0 -0.7566 0 -2.0 1e-06 
0.0 -0.7565 0 -2.0 1e-06 
0.0 -0.7564 0 -2.0 1e-06 
0.0 -0.7563 0 -2.0 1e-06 
0.0 -0.7562 0 -2.0 1e-06 
0.0 -0.7561 0 -2.0 1e-06 
0.0 -0.756 0 -2.0 1e-06 
0.0 -0.7559 0 -2.0 1e-06 
0.0 -0.7558 0 -2.0 1e-06 
0.0 -0.7557 0 -2.0 1e-06 
0.0 -0.7556 0 -2.0 1e-06 
0.0 -0.7555 0 -2.0 1e-06 
0.0 -0.7554 0 -2.0 1e-06 
0.0 -0.7553 0 -2.0 1e-06 
0.0 -0.7552 0 -2.0 1e-06 
0.0 -0.7551 0 -2.0 1e-06 
0.0 -0.755 0 -2.0 1e-06 
0.0 -0.7549 0 -2.0 1e-06 
0.0 -0.7548 0 -2.0 1e-06 
0.0 -0.7547 0 -2.0 1e-06 
0.0 -0.7546 0 -2.0 1e-06 
0.0 -0.7545 0 -2.0 1e-06 
0.0 -0.7544 0 -2.0 1e-06 
0.0 -0.7543 0 -2.0 1e-06 
0.0 -0.7542 0 -2.0 1e-06 
0.0 -0.7541 0 -2.0 1e-06 
0.0 -0.754 0 -2.0 1e-06 
0.0 -0.7539 0 -2.0 1e-06 
0.0 -0.7538 0 -2.0 1e-06 
0.0 -0.7537 0 -2.0 1e-06 
0.0 -0.7536 0 -2.0 1e-06 
0.0 -0.7535 0 -2.0 1e-06 
0.0 -0.7534 0 -2.0 1e-06 
0.0 -0.7533 0 -2.0 1e-06 
0.0 -0.7532 0 -2.0 1e-06 
0.0 -0.7531 0 -2.0 1e-06 
0.0 -0.753 0 -2.0 1e-06 
0.0 -0.7529 0 -2.0 1e-06 
0.0 -0.7528 0 -2.0 1e-06 
0.0 -0.7527 0 -2.0 1e-06 
0.0 -0.7526 0 -2.0 1e-06 
0.0 -0.7525 0 -2.0 1e-06 
0.0 -0.7524 0 -2.0 1e-06 
0.0 -0.7523 0 -2.0 1e-06 
0.0 -0.7522 0 -2.0 1e-06 
0.0 -0.7521 0 -2.0 1e-06 
0.0 -0.752 0 -2.0 1e-06 
0.0 -0.7519 0 -2.0 1e-06 
0.0 -0.7518 0 -2.0 1e-06 
0.0 -0.7517 0 -2.0 1e-06 
0.0 -0.7516 0 -2.0 1e-06 
0.0 -0.7515 0 -2.0 1e-06 
0.0 -0.7514 0 -2.0 1e-06 
0.0 -0.7513 0 -2.0 1e-06 
0.0 -0.7512 0 -2.0 1e-06 
0.0 -0.7511 0 -2.0 1e-06 
0.0 -0.751 0 -2.0 1e-06 
0.0 -0.7509 0 -2.0 1e-06 
0.0 -0.7508 0 -2.0 1e-06 
0.0 -0.7507 0 -2.0 1e-06 
0.0 -0.7506 0 -2.0 1e-06 
0.0 -0.7505 0 -2.0 1e-06 
0.0 -0.7504 0 -2.0 1e-06 
0.0 -0.7503 0 -2.0 1e-06 
0.0 -0.7502 0 -2.0 1e-06 
0.0 -0.7501 0 -2.0 1e-06 
0.0 -0.75 0 -2.0 1e-06 
0.0 -0.7499 0 -2.0 1e-06 
0.0 -0.7498 0 -2.0 1e-06 
0.0 -0.7497 0 -2.0 1e-06 
0.0 -0.7496 0 -2.0 1e-06 
0.0 -0.7495 0 -2.0 1e-06 
0.0 -0.7494 0 -2.0 1e-06 
0.0 -0.7493 0 -2.0 1e-06 
0.0 -0.7492 0 -2.0 1e-06 
0.0 -0.7491 0 -2.0 1e-06 
0.0 -0.749 0 -2.0 1e-06 
0.0 -0.7489 0 -2.0 1e-06 
0.0 -0.7488 0 -2.0 1e-06 
0.0 -0.7487 0 -2.0 1e-06 
0.0 -0.7486 0 -2.0 1e-06 
0.0 -0.7485 0 -2.0 1e-06 
0.0 -0.7484 0 -2.0 1e-06 
0.0 -0.7483 0 -2.0 1e-06 
0.0 -0.7482 0 -2.0 1e-06 
0.0 -0.7481 0 -2.0 1e-06 
0.0 -0.748 0 -2.0 1e-06 
0.0 -0.7479 0 -2.0 1e-06 
0.0 -0.7478 0 -2.0 1e-06 
0.0 -0.7477 0 -2.0 1e-06 
0.0 -0.7476 0 -2.0 1e-06 
0.0 -0.7475 0 -2.0 1e-06 
0.0 -0.7474 0 -2.0 1e-06 
0.0 -0.7473 0 -2.0 1e-06 
0.0 -0.7472 0 -2.0 1e-06 
0.0 -0.7471 0 -2.0 1e-06 
0.0 -0.747 0 -2.0 1e-06 
0.0 -0.7469 0 -2.0 1e-06 
0.0 -0.7468 0 -2.0 1e-06 
0.0 -0.7467 0 -2.0 1e-06 
0.0 -0.7466 0 -2.0 1e-06 
0.0 -0.7465 0 -2.0 1e-06 
0.0 -0.7464 0 -2.0 1e-06 
0.0 -0.7463 0 -2.0 1e-06 
0.0 -0.7462 0 -2.0 1e-06 
0.0 -0.7461 0 -2.0 1e-06 
0.0 -0.746 0 -2.0 1e-06 
0.0 -0.7459 0 -2.0 1e-06 
0.0 -0.7458 0 -2.0 1e-06 
0.0 -0.7457 0 -2.0 1e-06 
0.0 -0.7456 0 -2.0 1e-06 
0.0 -0.7455 0 -2.0 1e-06 
0.0 -0.7454 0 -2.0 1e-06 
0.0 -0.7453 0 -2.0 1e-06 
0.0 -0.7452 0 -2.0 1e-06 
0.0 -0.7451 0 -2.0 1e-06 
0.0 -0.745 0 -2.0 1e-06 
0.0 -0.7449 0 -2.0 1e-06 
0.0 -0.7448 0 -2.0 1e-06 
0.0 -0.7447 0 -2.0 1e-06 
0.0 -0.7446 0 -2.0 1e-06 
0.0 -0.7445 0 -2.0 1e-06 
0.0 -0.7444 0 -2.0 1e-06 
0.0 -0.7443 0 -2.0 1e-06 
0.0 -0.7442 0 -2.0 1e-06 
0.0 -0.7441 0 -2.0 1e-06 
0.0 -0.744 0 -2.0 1e-06 
0.0 -0.7439 0 -2.0 1e-06 
0.0 -0.7438 0 -2.0 1e-06 
0.0 -0.7437 0 -2.0 1e-06 
0.0 -0.7436 0 -2.0 1e-06 
0.0 -0.7435 0 -2.0 1e-06 
0.0 -0.7434 0 -2.0 1e-06 
0.0 -0.7433 0 -2.0 1e-06 
0.0 -0.7432 0 -2.0 1e-06 
0.0 -0.7431 0 -2.0 1e-06 
0.0 -0.743 0 -2.0 1e-06 
0.0 -0.7429 0 -2.0 1e-06 
0.0 -0.7428 0 -2.0 1e-06 
0.0 -0.7427 0 -2.0 1e-06 
0.0 -0.7426 0 -2.0 1e-06 
0.0 -0.7425 0 -2.0 1e-06 
0.0 -0.7424 0 -2.0 1e-06 
0.0 -0.7423 0 -2.0 1e-06 
0.0 -0.7422 0 -2.0 1e-06 
0.0 -0.7421 0 -2.0 1e-06 
0.0 -0.742 0 -2.0 1e-06 
0.0 -0.7419 0 -2.0 1e-06 
0.0 -0.7418 0 -2.0 1e-06 
0.0 -0.7417 0 -2.0 1e-06 
0.0 -0.7416 0 -2.0 1e-06 
0.0 -0.7415 0 -2.0 1e-06 
0.0 -0.7414 0 -2.0 1e-06 
0.0 -0.7413 0 -2.0 1e-06 
0.0 -0.7412 0 -2.0 1e-06 
0.0 -0.7411 0 -2.0 1e-06 
0.0 -0.741 0 -2.0 1e-06 
0.0 -0.7409 0 -2.0 1e-06 
0.0 -0.7408 0 -2.0 1e-06 
0.0 -0.7407 0 -2.0 1e-06 
0.0 -0.7406 0 -2.0 1e-06 
0.0 -0.7405 0 -2.0 1e-06 
0.0 -0.7404 0 -2.0 1e-06 
0.0 -0.7403 0 -2.0 1e-06 
0.0 -0.7402 0 -2.0 1e-06 
0.0 -0.7401 0 -2.0 1e-06 
0.0 -0.74 0 -2.0 1e-06 
0.0 -0.7399 0 -2.0 1e-06 
0.0 -0.7398 0 -2.0 1e-06 
0.0 -0.7397 0 -2.0 1e-06 
0.0 -0.7396 0 -2.0 1e-06 
0.0 -0.7395 0 -2.0 1e-06 
0.0 -0.7394 0 -2.0 1e-06 
0.0 -0.7393 0 -2.0 1e-06 
0.0 -0.7392 0 -2.0 1e-06 
0.0 -0.7391 0 -2.0 1e-06 
0.0 -0.739 0 -2.0 1e-06 
0.0 -0.7389 0 -2.0 1e-06 
0.0 -0.7388 0 -2.0 1e-06 
0.0 -0.7387 0 -2.0 1e-06 
0.0 -0.7386 0 -2.0 1e-06 
0.0 -0.7385 0 -2.0 1e-06 
0.0 -0.7384 0 -2.0 1e-06 
0.0 -0.7383 0 -2.0 1e-06 
0.0 -0.7382 0 -2.0 1e-06 
0.0 -0.7381 0 -2.0 1e-06 
0.0 -0.738 0 -2.0 1e-06 
0.0 -0.7379 0 -2.0 1e-06 
0.0 -0.7378 0 -2.0 1e-06 
0.0 -0.7377 0 -2.0 1e-06 
0.0 -0.7376 0 -2.0 1e-06 
0.0 -0.7375 0 -2.0 1e-06 
0.0 -0.7374 0 -2.0 1e-06 
0.0 -0.7373 0 -2.0 1e-06 
0.0 -0.7372 0 -2.0 1e-06 
0.0 -0.7371 0 -2.0 1e-06 
0.0 -0.737 0 -2.0 1e-06 
0.0 -0.7369 0 -2.0 1e-06 
0.0 -0.7368 0 -2.0 1e-06 
0.0 -0.7367 0 -2.0 1e-06 
0.0 -0.7366 0 -2.0 1e-06 
0.0 -0.7365 0 -2.0 1e-06 
0.0 -0.7364 0 -2.0 1e-06 
0.0 -0.7363 0 -2.0 1e-06 
0.0 -0.7362 0 -2.0 1e-06 
0.0 -0.7361 0 -2.0 1e-06 
0.0 -0.736 0 -2.0 1e-06 
0.0 -0.7359 0 -2.0 1e-06 
0.0 -0.7358 0 -2.0 1e-06 
0.0 -0.7357 0 -2.0 1e-06 
0.0 -0.7356 0 -2.0 1e-06 
0.0 -0.7355 0 -2.0 1e-06 
0.0 -0.7354 0 -2.0 1e-06 
0.0 -0.7353 0 -2.0 1e-06 
0.0 -0.7352 0 -2.0 1e-06 
0.0 -0.7351 0 -2.0 1e-06 
0.0 -0.735 0 -2.0 1e-06 
0.0 -0.7349 0 -2.0 1e-06 
0.0 -0.7348 0 -2.0 1e-06 
0.0 -0.7347 0 -2.0 1e-06 
0.0 -0.7346 0 -2.0 1e-06 
0.0 -0.7345 0 -2.0 1e-06 
0.0 -0.7344 0 -2.0 1e-06 
0.0 -0.7343 0 -2.0 1e-06 
0.0 -0.7342 0 -2.0 1e-06 
0.0 -0.7341 0 -2.0 1e-06 
0.0 -0.734 0 -2.0 1e-06 
0.0 -0.7339 0 -2.0 1e-06 
0.0 -0.7338 0 -2.0 1e-06 
0.0 -0.7337 0 -2.0 1e-06 
0.0 -0.7336 0 -2.0 1e-06 
0.0 -0.7335 0 -2.0 1e-06 
0.0 -0.7334 0 -2.0 1e-06 
0.0 -0.7333 0 -2.0 1e-06 
0.0 -0.7332 0 -2.0 1e-06 
0.0 -0.7331 0 -2.0 1e-06 
0.0 -0.733 0 -2.0 1e-06 
0.0 -0.7329 0 -2.0 1e-06 
0.0 -0.7328 0 -2.0 1e-06 
0.0 -0.7327 0 -2.0 1e-06 
0.0 -0.7326 0 -2.0 1e-06 
0.0 -0.7325 0 -2.0 1e-06 
0.0 -0.7324 0 -2.0 1e-06 
0.0 -0.7323 0 -2.0 1e-06 
0.0 -0.7322 0 -2.0 1e-06 
0.0 -0.7321 0 -2.0 1e-06 
0.0 -0.732 0 -2.0 1e-06 
0.0 -0.7319 0 -2.0 1e-06 
0.0 -0.7318 0 -2.0 1e-06 
0.0 -0.7317 0 -2.0 1e-06 
0.0 -0.7316 0 -2.0 1e-06 
0.0 -0.7315 0 -2.0 1e-06 
0.0 -0.7314 0 -2.0 1e-06 
0.0 -0.7313 0 -2.0 1e-06 
0.0 -0.7312 0 -2.0 1e-06 
0.0 -0.7311 0 -2.0 1e-06 
0.0 -0.731 0 -2.0 1e-06 
0.0 -0.7309 0 -2.0 1e-06 
0.0 -0.7308 0 -2.0 1e-06 
0.0 -0.7307 0 -2.0 1e-06 
0.0 -0.7306 0 -2.0 1e-06 
0.0 -0.7305 0 -2.0 1e-06 
0.0 -0.7304 0 -2.0 1e-06 
0.0 -0.7303 0 -2.0 1e-06 
0.0 -0.7302 0 -2.0 1e-06 
0.0 -0.7301 0 -2.0 1e-06 
0.0 -0.73 0 -2.0 1e-06 
0.0 -0.7299 0 -2.0 1e-06 
0.0 -0.7298 0 -2.0 1e-06 
0.0 -0.7297 0 -2.0 1e-06 
0.0 -0.7296 0 -2.0 1e-06 
0.0 -0.7295 0 -2.0 1e-06 
0.0 -0.7294 0 -2.0 1e-06 
0.0 -0.7293 0 -2.0 1e-06 
0.0 -0.7292 0 -2.0 1e-06 
0.0 -0.7291 0 -2.0 1e-06 
0.0 -0.729 0 -2.0 1e-06 
0.0 -0.7289 0 -2.0 1e-06 
0.0 -0.7288 0 -2.0 1e-06 
0.0 -0.7287 0 -2.0 1e-06 
0.0 -0.7286 0 -2.0 1e-06 
0.0 -0.7285 0 -2.0 1e-06 
0.0 -0.7284 0 -2.0 1e-06 
0.0 -0.7283 0 -2.0 1e-06 
0.0 -0.7282 0 -2.0 1e-06 
0.0 -0.7281 0 -2.0 1e-06 
0.0 -0.728 0 -2.0 1e-06 
0.0 -0.7279 0 -2.0 1e-06 
0.0 -0.7278 0 -2.0 1e-06 
0.0 -0.7277 0 -2.0 1e-06 
0.0 -0.7276 0 -2.0 1e-06 
0.0 -0.7275 0 -2.0 1e-06 
0.0 -0.7274 0 -2.0 1e-06 
0.0 -0.7273 0 -2.0 1e-06 
0.0 -0.7272 0 -2.0 1e-06 
0.0 -0.7271 0 -2.0 1e-06 
0.0 -0.727 0 -2.0 1e-06 
0.0 -0.7269 0 -2.0 1e-06 
0.0 -0.7268 0 -2.0 1e-06 
0.0 -0.7267 0 -2.0 1e-06 
0.0 -0.7266 0 -2.0 1e-06 
0.0 -0.7265 0 -2.0 1e-06 
0.0 -0.7264 0 -2.0 1e-06 
0.0 -0.7263 0 -2.0 1e-06 
0.0 -0.7262 0 -2.0 1e-06 
0.0 -0.7261 0 -2.0 1e-06 
0.0 -0.726 0 -2.0 1e-06 
0.0 -0.7259 0 -2.0 1e-06 
0.0 -0.7258 0 -2.0 1e-06 
0.0 -0.7257 0 -2.0 1e-06 
0.0 -0.7256 0 -2.0 1e-06 
0.0 -0.7255 0 -2.0 1e-06 
0.0 -0.7254 0 -2.0 1e-06 
0.0 -0.7253 0 -2.0 1e-06 
0.0 -0.7252 0 -2.0 1e-06 
0.0 -0.7251 0 -2.0 1e-06 
0.0 -0.725 0 -2.0 1e-06 
0.0 -0.7249 0 -2.0 1e-06 
0.0 -0.7248 0 -2.0 1e-06 
0.0 -0.7247 0 -2.0 1e-06 
0.0 -0.7246 0 -2.0 1e-06 
0.0 -0.7245 0 -2.0 1e-06 
0.0 -0.7244 0 -2.0 1e-06 
0.0 -0.7243 0 -2.0 1e-06 
0.0 -0.7242 0 -2.0 1e-06 
0.0 -0.7241 0 -2.0 1e-06 
0.0 -0.724 0 -2.0 1e-06 
0.0 -0.7239 0 -2.0 1e-06 
0.0 -0.7238 0 -2.0 1e-06 
0.0 -0.7237 0 -2.0 1e-06 
0.0 -0.7236 0 -2.0 1e-06 
0.0 -0.7235 0 -2.0 1e-06 
0.0 -0.7234 0 -2.0 1e-06 
0.0 -0.7233 0 -2.0 1e-06 
0.0 -0.7232 0 -2.0 1e-06 
0.0 -0.7231 0 -2.0 1e-06 
0.0 -0.723 0 -2.0 1e-06 
0.0 -0.7229 0 -2.0 1e-06 
0.0 -0.7228 0 -2.0 1e-06 
0.0 -0.7227 0 -2.0 1e-06 
0.0 -0.7226 0 -2.0 1e-06 
0.0 -0.7225 0 -2.0 1e-06 
0.0 -0.7224 0 -2.0 1e-06 
0.0 -0.7223 0 -2.0 1e-06 
0.0 -0.7222 0 -2.0 1e-06 
0.0 -0.7221 0 -2.0 1e-06 
0.0 -0.722 0 -2.0 1e-06 
0.0 -0.7219 0 -2.0 1e-06 
0.0 -0.7218 0 -2.0 1e-06 
0.0 -0.7217 0 -2.0 1e-06 
0.0 -0.7216 0 -2.0 1e-06 
0.0 -0.7215 0 -2.0 1e-06 
0.0 -0.7214 0 -2.0 1e-06 
0.0 -0.7213 0 -2.0 1e-06 
0.0 -0.7212 0 -2.0 1e-06 
0.0 -0.7211 0 -2.0 1e-06 
0.0 -0.721 0 -2.0 1e-06 
0.0 -0.7209 0 -2.0 1e-06 
0.0 -0.7208 0 -2.0 1e-06 
0.0 -0.7207 0 -2.0 1e-06 
0.0 -0.7206 0 -2.0 1e-06 
0.0 -0.7205 0 -2.0 1e-06 
0.0 -0.7204 0 -2.0 1e-06 
0.0 -0.7203 0 -2.0 1e-06 
0.0 -0.7202 0 -2.0 1e-06 
0.0 -0.7201 0 -2.0 1e-06 
0.0 -0.72 0 -2.0 1e-06 
0.0 -0.7199 0 -2.0 1e-06 
0.0 -0.7198 0 -2.0 1e-06 
0.0 -0.7197 0 -2.0 1e-06 
0.0 -0.7196 0 -2.0 1e-06 
0.0 -0.7195 0 -2.0 1e-06 
0.0 -0.7194 0 -2.0 1e-06 
0.0 -0.7193 0 -2.0 1e-06 
0.0 -0.7192 0 -2.0 1e-06 
0.0 -0.7191 0 -2.0 1e-06 
0.0 -0.719 0 -2.0 1e-06 
0.0 -0.7189 0 -2.0 1e-06 
0.0 -0.7188 0 -2.0 1e-06 
0.0 -0.7187 0 -2.0 1e-06 
0.0 -0.7186 0 -2.0 1e-06 
0.0 -0.7185 0 -2.0 1e-06 
0.0 -0.7184 0 -2.0 1e-06 
0.0 -0.7183 0 -2.0 1e-06 
0.0 -0.7182 0 -2.0 1e-06 
0.0 -0.7181 0 -2.0 1e-06 
0.0 -0.718 0 -2.0 1e-06 
0.0 -0.7179 0 -2.0 1e-06 
0.0 -0.7178 0 -2.0 1e-06 
0.0 -0.7177 0 -2.0 1e-06 
0.0 -0.7176 0 -2.0 1e-06 
0.0 -0.7175 0 -2.0 1e-06 
0.0 -0.7174 0 -2.0 1e-06 
0.0 -0.7173 0 -2.0 1e-06 
0.0 -0.7172 0 -2.0 1e-06 
0.0 -0.7171 0 -2.0 1e-06 
0.0 -0.717 0 -2.0 1e-06 
0.0 -0.7169 0 -2.0 1e-06 
0.0 -0.7168 0 -2.0 1e-06 
0.0 -0.7167 0 -2.0 1e-06 
0.0 -0.7166 0 -2.0 1e-06 
0.0 -0.7165 0 -2.0 1e-06 
0.0 -0.7164 0 -2.0 1e-06 
0.0 -0.7163 0 -2.0 1e-06 
0.0 -0.7162 0 -2.0 1e-06 
0.0 -0.7161 0 -2.0 1e-06 
0.0 -0.716 0 -2.0 1e-06 
0.0 -0.7159 0 -2.0 1e-06 
0.0 -0.7158 0 -2.0 1e-06 
0.0 -0.7157 0 -2.0 1e-06 
0.0 -0.7156 0 -2.0 1e-06 
0.0 -0.7155 0 -2.0 1e-06 
0.0 -0.7154 0 -2.0 1e-06 
0.0 -0.7153 0 -2.0 1e-06 
0.0 -0.7152 0 -2.0 1e-06 
0.0 -0.7151 0 -2.0 1e-06 
0.0 -0.715 0 -2.0 1e-06 
0.0 -0.7149 0 -2.0 1e-06 
0.0 -0.7148 0 -2.0 1e-06 
0.0 -0.7147 0 -2.0 1e-06 
0.0 -0.7146 0 -2.0 1e-06 
0.0 -0.7145 0 -2.0 1e-06 
0.0 -0.7144 0 -2.0 1e-06 
0.0 -0.7143 0 -2.0 1e-06 
0.0 -0.7142 0 -2.0 1e-06 
0.0 -0.7141 0 -2.0 1e-06 
0.0 -0.714 0 -2.0 1e-06 
0.0 -0.7139 0 -2.0 1e-06 
0.0 -0.7138 0 -2.0 1e-06 
0.0 -0.7137 0 -2.0 1e-06 
0.0 -0.7136 0 -2.0 1e-06 
0.0 -0.7135 0 -2.0 1e-06 
0.0 -0.7134 0 -2.0 1e-06 
0.0 -0.7133 0 -2.0 1e-06 
0.0 -0.7132 0 -2.0 1e-06 
0.0 -0.7131 0 -2.0 1e-06 
0.0 -0.713 0 -2.0 1e-06 
0.0 -0.7129 0 -2.0 1e-06 
0.0 -0.7128 0 -2.0 1e-06 
0.0 -0.7127 0 -2.0 1e-06 
0.0 -0.7126 0 -2.0 1e-06 
0.0 -0.7125 0 -2.0 1e-06 
0.0 -0.7124 0 -2.0 1e-06 
0.0 -0.7123 0 -2.0 1e-06 
0.0 -0.7122 0 -2.0 1e-06 
0.0 -0.7121 0 -2.0 1e-06 
0.0 -0.712 0 -2.0 1e-06 
0.0 -0.7119 0 -2.0 1e-06 
0.0 -0.7118 0 -2.0 1e-06 
0.0 -0.7117 0 -2.0 1e-06 
0.0 -0.7116 0 -2.0 1e-06 
0.0 -0.7115 0 -2.0 1e-06 
0.0 -0.7114 0 -2.0 1e-06 
0.0 -0.7113 0 -2.0 1e-06 
0.0 -0.7112 0 -2.0 1e-06 
0.0 -0.7111 0 -2.0 1e-06 
0.0 -0.711 0 -2.0 1e-06 
0.0 -0.7109 0 -2.0 1e-06 
0.0 -0.7108 0 -2.0 1e-06 
0.0 -0.7107 0 -2.0 1e-06 
0.0 -0.7106 0 -2.0 1e-06 
0.0 -0.7105 0 -2.0 1e-06 
0.0 -0.7104 0 -2.0 1e-06 
0.0 -0.7103 0 -2.0 1e-06 
0.0 -0.7102 0 -2.0 1e-06 
0.0 -0.7101 0 -2.0 1e-06 
0.0 -0.71 0 -2.0 1e-06 
0.0 -0.7099 0 -2.0 1e-06 
0.0 -0.7098 0 -2.0 1e-06 
0.0 -0.7097 0 -2.0 1e-06 
0.0 -0.7096 0 -2.0 1e-06 
0.0 -0.7095 0 -2.0 1e-06 
0.0 -0.7094 0 -2.0 1e-06 
0.0 -0.7093 0 -2.0 1e-06 
0.0 -0.7092 0 -2.0 1e-06 
0.0 -0.7091 0 -2.0 1e-06 
0.0 -0.709 0 -2.0 1e-06 
0.0 -0.7089 0 -2.0 1e-06 
0.0 -0.7088 0 -2.0 1e-06 
0.0 -0.7087 0 -2.0 1e-06 
0.0 -0.7086 0 -2.0 1e-06 
0.0 -0.7085 0 -2.0 1e-06 
0.0 -0.7084 0 -2.0 1e-06 
0.0 -0.7083 0 -2.0 1e-06 
0.0 -0.7082 0 -2.0 1e-06 
0.0 -0.7081 0 -2.0 1e-06 
0.0 -0.708 0 -2.0 1e-06 
0.0 -0.7079 0 -2.0 1e-06 
0.0 -0.7078 0 -2.0 1e-06 
0.0 -0.7077 0 -2.0 1e-06 
0.0 -0.7076 0 -2.0 1e-06 
0.0 -0.7075 0 -2.0 1e-06 
0.0 -0.7074 0 -2.0 1e-06 
0.0 -0.7073 0 -2.0 1e-06 
0.0 -0.7072 0 -2.0 1e-06 
0.0 -0.7071 0 -2.0 1e-06 
0.0 -0.707 0 -2.0 1e-06 
0.0 -0.7069 0 -2.0 1e-06 
0.0 -0.7068 0 -2.0 1e-06 
0.0 -0.7067 0 -2.0 1e-06 
0.0 -0.7066 0 -2.0 1e-06 
0.0 -0.7065 0 -2.0 1e-06 
0.0 -0.7064 0 -2.0 1e-06 
0.0 -0.7063 0 -2.0 1e-06 
0.0 -0.7062 0 -2.0 1e-06 
0.0 -0.7061 0 -2.0 1e-06 
0.0 -0.706 0 -2.0 1e-06 
0.0 -0.7059 0 -2.0 1e-06 
0.0 -0.7058 0 -2.0 1e-06 
0.0 -0.7057 0 -2.0 1e-06 
0.0 -0.7056 0 -2.0 1e-06 
0.0 -0.7055 0 -2.0 1e-06 
0.0 -0.7054 0 -2.0 1e-06 
0.0 -0.7053 0 -2.0 1e-06 
0.0 -0.7052 0 -2.0 1e-06 
0.0 -0.7051 0 -2.0 1e-06 
0.0 -0.705 0 -2.0 1e-06 
0.0 -0.7049 0 -2.0 1e-06 
0.0 -0.7048 0 -2.0 1e-06 
0.0 -0.7047 0 -2.0 1e-06 
0.0 -0.7046 0 -2.0 1e-06 
0.0 -0.7045 0 -2.0 1e-06 
0.0 -0.7044 0 -2.0 1e-06 
0.0 -0.7043 0 -2.0 1e-06 
0.0 -0.7042 0 -2.0 1e-06 
0.0 -0.7041 0 -2.0 1e-06 
0.0 -0.704 0 -2.0 1e-06 
0.0 -0.7039 0 -2.0 1e-06 
0.0 -0.7038 0 -2.0 1e-06 
0.0 -0.7037 0 -2.0 1e-06 
0.0 -0.7036 0 -2.0 1e-06 
0.0 -0.7035 0 -2.0 1e-06 
0.0 -0.7034 0 -2.0 1e-06 
0.0 -0.7033 0 -2.0 1e-06 
0.0 -0.7032 0 -2.0 1e-06 
0.0 -0.7031 0 -2.0 1e-06 
0.0 -0.703 0 -2.0 1e-06 
0.0 -0.7029 0 -2.0 1e-06 
0.0 -0.7028 0 -2.0 1e-06 
0.0 -0.7027 0 -2.0 1e-06 
0.0 -0.7026 0 -2.0 1e-06 
0.0 -0.7025 0 -2.0 1e-06 
0.0 -0.7024 0 -2.0 1e-06 
0.0 -0.7023 0 -2.0 1e-06 
0.0 -0.7022 0 -2.0 1e-06 
0.0 -0.7021 0 -2.0 1e-06 
0.0 -0.702 0 -2.0 1e-06 
0.0 -0.7019 0 -2.0 1e-06 
0.0 -0.7018 0 -2.0 1e-06 
0.0 -0.7017 0 -2.0 1e-06 
0.0 -0.7016 0 -2.0 1e-06 
0.0 -0.7015 0 -2.0 1e-06 
0.0 -0.7014 0 -2.0 1e-06 
0.0 -0.7013 0 -2.0 1e-06 
0.0 -0.7012 0 -2.0 1e-06 
0.0 -0.7011 0 -2.0 1e-06 
0.0 -0.701 0 -2.0 1e-06 
0.0 -0.7009 0 -2.0 1e-06 
0.0 -0.7008 0 -2.0 1e-06 
0.0 -0.7007 0 -2.0 1e-06 
0.0 -0.7006 0 -2.0 1e-06 
0.0 -0.7005 0 -2.0 1e-06 
0.0 -0.7004 0 -2.0 1e-06 
0.0 -0.7003 0 -2.0 1e-06 
0.0 -0.7002 0 -2.0 1e-06 
0.0 -0.7001 0 -2.0 1e-06 
0.0 -0.7 0 -2.0 1e-06 
0.0 -0.6999 0 -2.0 1e-06 
0.0 -0.6998 0 -2.0 1e-06 
0.0 -0.6997 0 -2.0 1e-06 
0.0 -0.6996 0 -2.0 1e-06 
0.0 -0.6995 0 -2.0 1e-06 
0.0 -0.6994 0 -2.0 1e-06 
0.0 -0.6993 0 -2.0 1e-06 
0.0 -0.6992 0 -2.0 1e-06 
0.0 -0.6991 0 -2.0 1e-06 
0.0 -0.699 0 -2.0 1e-06 
0.0 -0.6989 0 -2.0 1e-06 
0.0 -0.6988 0 -2.0 1e-06 
0.0 -0.6987 0 -2.0 1e-06 
0.0 -0.6986 0 -2.0 1e-06 
0.0 -0.6985 0 -2.0 1e-06 
0.0 -0.6984 0 -2.0 1e-06 
0.0 -0.6983 0 -2.0 1e-06 
0.0 -0.6982 0 -2.0 1e-06 
0.0 -0.6981 0 -2.0 1e-06 
0.0 -0.698 0 -2.0 1e-06 
0.0 -0.6979 0 -2.0 1e-06 
0.0 -0.6978 0 -2.0 1e-06 
0.0 -0.6977 0 -2.0 1e-06 
0.0 -0.6976 0 -2.0 1e-06 
0.0 -0.6975 0 -2.0 1e-06 
0.0 -0.6974 0 -2.0 1e-06 
0.0 -0.6973 0 -2.0 1e-06 
0.0 -0.6972 0 -2.0 1e-06 
0.0 -0.6971 0 -2.0 1e-06 
0.0 -0.697 0 -2.0 1e-06 
0.0 -0.6969 0 -2.0 1e-06 
0.0 -0.6968 0 -2.0 1e-06 
0.0 -0.6967 0 -2.0 1e-06 
0.0 -0.6966 0 -2.0 1e-06 
0.0 -0.6965 0 -2.0 1e-06 
0.0 -0.6964 0 -2.0 1e-06 
0.0 -0.6963 0 -2.0 1e-06 
0.0 -0.6962 0 -2.0 1e-06 
0.0 -0.6961 0 -2.0 1e-06 
0.0 -0.696 0 -2.0 1e-06 
0.0 -0.6959 0 -2.0 1e-06 
0.0 -0.6958 0 -2.0 1e-06 
0.0 -0.6957 0 -2.0 1e-06 
0.0 -0.6956 0 -2.0 1e-06 
0.0 -0.6955 0 -2.0 1e-06 
0.0 -0.6954 0 -2.0 1e-06 
0.0 -0.6953 0 -2.0 1e-06 
0.0 -0.6952 0 -2.0 1e-06 
0.0 -0.6951 0 -2.0 1e-06 
0.0 -0.695 0 -2.0 1e-06 
0.0 -0.6949 0 -2.0 1e-06 
0.0 -0.6948 0 -2.0 1e-06 
0.0 -0.6947 0 -2.0 1e-06 
0.0 -0.6946 0 -2.0 1e-06 
0.0 -0.6945 0 -2.0 1e-06 
0.0 -0.6944 0 -2.0 1e-06 
0.0 -0.6943 0 -2.0 1e-06 
0.0 -0.6942 0 -2.0 1e-06 
0.0 -0.6941 0 -2.0 1e-06 
0.0 -0.694 0 -2.0 1e-06 
0.0 -0.6939 0 -2.0 1e-06 
0.0 -0.6938 0 -2.0 1e-06 
0.0 -0.6937 0 -2.0 1e-06 
0.0 -0.6936 0 -2.0 1e-06 
0.0 -0.6935 0 -2.0 1e-06 
0.0 -0.6934 0 -2.0 1e-06 
0.0 -0.6933 0 -2.0 1e-06 
0.0 -0.6932 0 -2.0 1e-06 
0.0 -0.6931 0 -2.0 1e-06 
0.0 -0.693 0 -2.0 1e-06 
0.0 -0.6929 0 -2.0 1e-06 
0.0 -0.6928 0 -2.0 1e-06 
0.0 -0.6927 0 -2.0 1e-06 
0.0 -0.6926 0 -2.0 1e-06 
0.0 -0.6925 0 -2.0 1e-06 
0.0 -0.6924 0 -2.0 1e-06 
0.0 -0.6923 0 -2.0 1e-06 
0.0 -0.6922 0 -2.0 1e-06 
0.0 -0.6921 0 -2.0 1e-06 
0.0 -0.692 0 -2.0 1e-06 
0.0 -0.6919 0 -2.0 1e-06 
0.0 -0.6918 0 -2.0 1e-06 
0.0 -0.6917 0 -2.0 1e-06 
0.0 -0.6916 0 -2.0 1e-06 
0.0 -0.6915 0 -2.0 1e-06 
0.0 -0.6914 0 -2.0 1e-06 
0.0 -0.6913 0 -2.0 1e-06 
0.0 -0.6912 0 -2.0 1e-06 
0.0 -0.6911 0 -2.0 1e-06 
0.0 -0.691 0 -2.0 1e-06 
0.0 -0.6909 0 -2.0 1e-06 
0.0 -0.6908 0 -2.0 1e-06 
0.0 -0.6907 0 -2.0 1e-06 
0.0 -0.6906 0 -2.0 1e-06 
0.0 -0.6905 0 -2.0 1e-06 
0.0 -0.6904 0 -2.0 1e-06 
0.0 -0.6903 0 -2.0 1e-06 
0.0 -0.6902 0 -2.0 1e-06 
0.0 -0.6901 0 -2.0 1e-06 
0.0 -0.69 0 -2.0 1e-06 
0.0 -0.6899 0 -2.0 1e-06 
0.0 -0.6898 0 -2.0 1e-06 
0.0 -0.6897 0 -2.0 1e-06 
0.0 -0.6896 0 -2.0 1e-06 
0.0 -0.6895 0 -2.0 1e-06 
0.0 -0.6894 0 -2.0 1e-06 
0.0 -0.6893 0 -2.0 1e-06 
0.0 -0.6892 0 -2.0 1e-06 
0.0 -0.6891 0 -2.0 1e-06 
0.0 -0.689 0 -2.0 1e-06 
0.0 -0.6889 0 -2.0 1e-06 
0.0 -0.6888 0 -2.0 1e-06 
0.0 -0.6887 0 -2.0 1e-06 
0.0 -0.6886 0 -2.0 1e-06 
0.0 -0.6885 0 -2.0 1e-06 
0.0 -0.6884 0 -2.0 1e-06 
0.0 -0.6883 0 -2.0 1e-06 
0.0 -0.6882 0 -2.0 1e-06 
0.0 -0.6881 0 -2.0 1e-06 
0.0 -0.688 0 -2.0 1e-06 
0.0 -0.6879 0 -2.0 1e-06 
0.0 -0.6878 0 -2.0 1e-06 
0.0 -0.6877 0 -2.0 1e-06 
0.0 -0.6876 0 -2.0 1e-06 
0.0 -0.6875 0 -2.0 1e-06 
0.0 -0.6874 0 -2.0 1e-06 
0.0 -0.6873 0 -2.0 1e-06 
0.0 -0.6872 0 -2.0 1e-06 
0.0 -0.6871 0 -2.0 1e-06 
0.0 -0.687 0 -2.0 1e-06 
0.0 -0.6869 0 -2.0 1e-06 
0.0 -0.6868 0 -2.0 1e-06 
0.0 -0.6867 0 -2.0 1e-06 
0.0 -0.6866 0 -2.0 1e-06 
0.0 -0.6865 0 -2.0 1e-06 
0.0 -0.6864 0 -2.0 1e-06 
0.0 -0.6863 0 -2.0 1e-06 
0.0 -0.6862 0 -2.0 1e-06 
0.0 -0.6861 0 -2.0 1e-06 
0.0 -0.686 0 -2.0 1e-06 
0.0 -0.6859 0 -2.0 1e-06 
0.0 -0.6858 0 -2.0 1e-06 
0.0 -0.6857 0 -2.0 1e-06 
0.0 -0.6856 0 -2.0 1e-06 
0.0 -0.6855 0 -2.0 1e-06 
0.0 -0.6854 0 -2.0 1e-06 
0.0 -0.6853 0 -2.0 1e-06 
0.0 -0.6852 0 -2.0 1e-06 
0.0 -0.6851 0 -2.0 1e-06 
0.0 -0.685 0 -2.0 1e-06 
0.0 -0.6849 0 -2.0 1e-06 
0.0 -0.6848 0 -2.0 1e-06 
0.0 -0.6847 0 -2.0 1e-06 
0.0 -0.6846 0 -2.0 1e-06 
0.0 -0.6845 0 -2.0 1e-06 
0.0 -0.6844 0 -2.0 1e-06 
0.0 -0.6843 0 -2.0 1e-06 
0.0 -0.6842 0 -2.0 1e-06 
0.0 -0.6841 0 -2.0 1e-06 
0.0 -0.684 0 -2.0 1e-06 
0.0 -0.6839 0 -2.0 1e-06 
0.0 -0.6838 0 -2.0 1e-06 
0.0 -0.6837 0 -2.0 1e-06 
0.0 -0.6836 0 -2.0 1e-06 
0.0 -0.6835 0 -2.0 1e-06 
0.0 -0.6834 0 -2.0 1e-06 
0.0 -0.6833 0 -2.0 1e-06 
0.0 -0.6832 0 -2.0 1e-06 
0.0 -0.6831 0 -2.0 1e-06 
0.0 -0.683 0 -2.0 1e-06 
0.0 -0.6829 0 -2.0 1e-06 
0.0 -0.6828 0 -2.0 1e-06 
0.0 -0.6827 0 -2.0 1e-06 
0.0 -0.6826 0 -2.0 1e-06 
0.0 -0.6825 0 -2.0 1e-06 
0.0 -0.6824 0 -2.0 1e-06 
0.0 -0.6823 0 -2.0 1e-06 
0.0 -0.6822 0 -2.0 1e-06 
0.0 -0.6821 0 -2.0 1e-06 
0.0 -0.682 0 -2.0 1e-06 
0.0 -0.6819 0 -2.0 1e-06 
0.0 -0.6818 0 -2.0 1e-06 
0.0 -0.6817 0 -2.0 1e-06 
0.0 -0.6816 0 -2.0 1e-06 
0.0 -0.6815 0 -2.0 1e-06 
0.0 -0.6814 0 -2.0 1e-06 
0.0 -0.6813 0 -2.0 1e-06 
0.0 -0.6812 0 -2.0 1e-06 
0.0 -0.6811 0 -2.0 1e-06 
0.0 -0.681 0 -2.0 1e-06 
0.0 -0.6809 0 -2.0 1e-06 
0.0 -0.6808 0 -2.0 1e-06 
0.0 -0.6807 0 -2.0 1e-06 
0.0 -0.6806 0 -2.0 1e-06 
0.0 -0.6805 0 -2.0 1e-06 
0.0 -0.6804 0 -2.0 1e-06 
0.0 -0.6803 0 -2.0 1e-06 
0.0 -0.6802 0 -2.0 1e-06 
0.0 -0.6801 0 -2.0 1e-06 
0.0 -0.68 0 -2.0 1e-06 
0.0 -0.6799 0 -2.0 1e-06 
0.0 -0.6798 0 -2.0 1e-06 
0.0 -0.6797 0 -2.0 1e-06 
0.0 -0.6796 0 -2.0 1e-06 
0.0 -0.6795 0 -2.0 1e-06 
0.0 -0.6794 0 -2.0 1e-06 
0.0 -0.6793 0 -2.0 1e-06 
0.0 -0.6792 0 -2.0 1e-06 
0.0 -0.6791 0 -2.0 1e-06 
0.0 -0.679 0 -2.0 1e-06 
0.0 -0.6789 0 -2.0 1e-06 
0.0 -0.6788 0 -2.0 1e-06 
0.0 -0.6787 0 -2.0 1e-06 
0.0 -0.6786 0 -2.0 1e-06 
0.0 -0.6785 0 -2.0 1e-06 
0.0 -0.6784 0 -2.0 1e-06 
0.0 -0.6783 0 -2.0 1e-06 
0.0 -0.6782 0 -2.0 1e-06 
0.0 -0.6781 0 -2.0 1e-06 
0.0 -0.678 0 -2.0 1e-06 
0.0 -0.6779 0 -2.0 1e-06 
0.0 -0.6778 0 -2.0 1e-06 
0.0 -0.6777 0 -2.0 1e-06 
0.0 -0.6776 0 -2.0 1e-06 
0.0 -0.6775 0 -2.0 1e-06 
0.0 -0.6774 0 -2.0 1e-06 
0.0 -0.6773 0 -2.0 1e-06 
0.0 -0.6772 0 -2.0 1e-06 
0.0 -0.6771 0 -2.0 1e-06 
0.0 -0.677 0 -2.0 1e-06 
0.0 -0.6769 0 -2.0 1e-06 
0.0 -0.6768 0 -2.0 1e-06 
0.0 -0.6767 0 -2.0 1e-06 
0.0 -0.6766 0 -2.0 1e-06 
0.0 -0.6765 0 -2.0 1e-06 
0.0 -0.6764 0 -2.0 1e-06 
0.0 -0.6763 0 -2.0 1e-06 
0.0 -0.6762 0 -2.0 1e-06 
0.0 -0.6761 0 -2.0 1e-06 
0.0 -0.676 0 -2.0 1e-06 
0.0 -0.6759 0 -2.0 1e-06 
0.0 -0.6758 0 -2.0 1e-06 
0.0 -0.6757 0 -2.0 1e-06 
0.0 -0.6756 0 -2.0 1e-06 
0.0 -0.6755 0 -2.0 1e-06 
0.0 -0.6754 0 -2.0 1e-06 
0.0 -0.6753 0 -2.0 1e-06 
0.0 -0.6752 0 -2.0 1e-06 
0.0 -0.6751 0 -2.0 1e-06 
0.0 -0.675 0 -2.0 1e-06 
0.0 -0.6749 0 -2.0 1e-06 
0.0 -0.6748 0 -2.0 1e-06 
0.0 -0.6747 0 -2.0 1e-06 
0.0 -0.6746 0 -2.0 1e-06 
0.0 -0.6745 0 -2.0 1e-06 
0.0 -0.6744 0 -2.0 1e-06 
0.0 -0.6743 0 -2.0 1e-06 
0.0 -0.6742 0 -2.0 1e-06 
0.0 -0.6741 0 -2.0 1e-06 
0.0 -0.674 0 -2.0 1e-06 
0.0 -0.6739 0 -2.0 1e-06 
0.0 -0.6738 0 -2.0 1e-06 
0.0 -0.6737 0 -2.0 1e-06 
0.0 -0.6736 0 -2.0 1e-06 
0.0 -0.6735 0 -2.0 1e-06 
0.0 -0.6734 0 -2.0 1e-06 
0.0 -0.6733 0 -2.0 1e-06 
0.0 -0.6732 0 -2.0 1e-06 
0.0 -0.6731 0 -2.0 1e-06 
0.0 -0.673 0 -2.0 1e-06 
0.0 -0.6729 0 -2.0 1e-06 
0.0 -0.6728 0 -2.0 1e-06 
0.0 -0.6727 0 -2.0 1e-06 
0.0 -0.6726 0 -2.0 1e-06 
0.0 -0.6725 0 -2.0 1e-06 
0.0 -0.6724 0 -2.0 1e-06 
0.0 -0.6723 0 -2.0 1e-06 
0.0 -0.6722 0 -2.0 1e-06 
0.0 -0.6721 0 -2.0 1e-06 
0.0 -0.672 0 -2.0 1e-06 
0.0 -0.6719 0 -2.0 1e-06 
0.0 -0.6718 0 -2.0 1e-06 
0.0 -0.6717 0 -2.0 1e-06 
0.0 -0.6716 0 -2.0 1e-06 
0.0 -0.6715 0 -2.0 1e-06 
0.0 -0.6714 0 -2.0 1e-06 
0.0 -0.6713 0 -2.0 1e-06 
0.0 -0.6712 0 -2.0 1e-06 
0.0 -0.6711 0 -2.0 1e-06 
0.0 -0.671 0 -2.0 1e-06 
0.0 -0.6709 0 -2.0 1e-06 
0.0 -0.6708 0 -2.0 1e-06 
0.0 -0.6707 0 -2.0 1e-06 
0.0 -0.6706 0 -2.0 1e-06 
0.0 -0.6705 0 -2.0 1e-06 
0.0 -0.6704 0 -2.0 1e-06 
0.0 -0.6703 0 -2.0 1e-06 
0.0 -0.6702 0 -2.0 1e-06 
0.0 -0.6701 0 -2.0 1e-06 
0.0 -0.67 0 -2.0 1e-06 
0.0 -0.6699 0 -2.0 1e-06 
0.0 -0.6698 0 -2.0 1e-06 
0.0 -0.6697 0 -2.0 1e-06 
0.0 -0.6696 0 -2.0 1e-06 
0.0 -0.6695 0 -2.0 1e-06 
0.0 -0.6694 0 -2.0 1e-06 
0.0 -0.6693 0 -2.0 1e-06 
0.0 -0.6692 0 -2.0 1e-06 
0.0 -0.6691 0 -2.0 1e-06 
0.0 -0.669 0 -2.0 1e-06 
0.0 -0.6689 0 -2.0 1e-06 
0.0 -0.6688 0 -2.0 1e-06 
0.0 -0.6687 0 -2.0 1e-06 
0.0 -0.6686 0 -2.0 1e-06 
0.0 -0.6685 0 -2.0 1e-06 
0.0 -0.6684 0 -2.0 1e-06 
0.0 -0.6683 0 -2.0 1e-06 
0.0 -0.6682 0 -2.0 1e-06 
0.0 -0.6681 0 -2.0 1e-06 
0.0 -0.668 0 -2.0 1e-06 
0.0 -0.6679 0 -2.0 1e-06 
0.0 -0.6678 0 -2.0 1e-06 
0.0 -0.6677 0 -2.0 1e-06 
0.0 -0.6676 0 -2.0 1e-06 
0.0 -0.6675 0 -2.0 1e-06 
0.0 -0.6674 0 -2.0 1e-06 
0.0 -0.6673 0 -2.0 1e-06 
0.0 -0.6672 0 -2.0 1e-06 
0.0 -0.6671 0 -2.0 1e-06 
0.0 -0.667 0 -2.0 1e-06 
0.0 -0.6669 0 -2.0 1e-06 
0.0 -0.6668 0 -2.0 1e-06 
0.0 -0.6667 0 -2.0 1e-06 
0.0 -0.6666 0 -2.0 1e-06 
0.0 -0.6665 0 -2.0 1e-06 
0.0 -0.6664 0 -2.0 1e-06 
0.0 -0.6663 0 -2.0 1e-06 
0.0 -0.6662 0 -2.0 1e-06 
0.0 -0.6661 0 -2.0 1e-06 
0.0 -0.666 0 -2.0 1e-06 
0.0 -0.6659 0 -2.0 1e-06 
0.0 -0.6658 0 -2.0 1e-06 
0.0 -0.6657 0 -2.0 1e-06 
0.0 -0.6656 0 -2.0 1e-06 
0.0 -0.6655 0 -2.0 1e-06 
0.0 -0.6654 0 -2.0 1e-06 
0.0 -0.6653 0 -2.0 1e-06 
0.0 -0.6652 0 -2.0 1e-06 
0.0 -0.6651 0 -2.0 1e-06 
0.0 -0.665 0 -2.0 1e-06 
0.0 -0.6649 0 -2.0 1e-06 
0.0 -0.6648 0 -2.0 1e-06 
0.0 -0.6647 0 -2.0 1e-06 
0.0 -0.6646 0 -2.0 1e-06 
0.0 -0.6645 0 -2.0 1e-06 
0.0 -0.6644 0 -2.0 1e-06 
0.0 -0.6643 0 -2.0 1e-06 
0.0 -0.6642 0 -2.0 1e-06 
0.0 -0.6641 0 -2.0 1e-06 
0.0 -0.664 0 -2.0 1e-06 
0.0 -0.6639 0 -2.0 1e-06 
0.0 -0.6638 0 -2.0 1e-06 
0.0 -0.6637 0 -2.0 1e-06 
0.0 -0.6636 0 -2.0 1e-06 
0.0 -0.6635 0 -2.0 1e-06 
0.0 -0.6634 0 -2.0 1e-06 
0.0 -0.6633 0 -2.0 1e-06 
0.0 -0.6632 0 -2.0 1e-06 
0.0 -0.6631 0 -2.0 1e-06 
0.0 -0.663 0 -2.0 1e-06 
0.0 -0.6629 0 -2.0 1e-06 
0.0 -0.6628 0 -2.0 1e-06 
0.0 -0.6627 0 -2.0 1e-06 
0.0 -0.6626 0 -2.0 1e-06 
0.0 -0.6625 0 -2.0 1e-06 
0.0 -0.6624 0 -2.0 1e-06 
0.0 -0.6623 0 -2.0 1e-06 
0.0 -0.6622 0 -2.0 1e-06 
0.0 -0.6621 0 -2.0 1e-06 
0.0 -0.662 0 -2.0 1e-06 
0.0 -0.6619 0 -2.0 1e-06 
0.0 -0.6618 0 -2.0 1e-06 
0.0 -0.6617 0 -2.0 1e-06 
0.0 -0.6616 0 -2.0 1e-06 
0.0 -0.6615 0 -2.0 1e-06 
0.0 -0.6614 0 -2.0 1e-06 
0.0 -0.6613 0 -2.0 1e-06 
0.0 -0.6612 0 -2.0 1e-06 
0.0 -0.6611 0 -2.0 1e-06 
0.0 -0.661 0 -2.0 1e-06 
0.0 -0.6609 0 -2.0 1e-06 
0.0 -0.6608 0 -2.0 1e-06 
0.0 -0.6607 0 -2.0 1e-06 
0.0 -0.6606 0 -2.0 1e-06 
0.0 -0.6605 0 -2.0 1e-06 
0.0 -0.6604 0 -2.0 1e-06 
0.0 -0.6603 0 -2.0 1e-06 
0.0 -0.6602 0 -2.0 1e-06 
0.0 -0.6601 0 -2.0 1e-06 
0.0 -0.66 0 -2.0 1e-06 
0.0 -0.6599 0 -2.0 1e-06 
0.0 -0.6598 0 -2.0 1e-06 
0.0 -0.6597 0 -2.0 1e-06 
0.0 -0.6596 0 -2.0 1e-06 
0.0 -0.6595 0 -2.0 1e-06 
0.0 -0.6594 0 -2.0 1e-06 
0.0 -0.6593 0 -2.0 1e-06 
0.0 -0.6592 0 -2.0 1e-06 
0.0 -0.6591 0 -2.0 1e-06 
0.0 -0.659 0 -2.0 1e-06 
0.0 -0.6589 0 -2.0 1e-06 
0.0 -0.6588 0 -2.0 1e-06 
0.0 -0.6587 0 -2.0 1e-06 
0.0 -0.6586 0 -2.0 1e-06 
0.0 -0.6585 0 -2.0 1e-06 
0.0 -0.6584 0 -2.0 1e-06 
0.0 -0.6583 0 -2.0 1e-06 
0.0 -0.6582 0 -2.0 1e-06 
0.0 -0.6581 0 -2.0 1e-06 
0.0 -0.658 0 -2.0 1e-06 
0.0 -0.6579 0 -2.0 1e-06 
0.0 -0.6578 0 -2.0 1e-06 
0.0 -0.6577 0 -2.0 1e-06 
0.0 -0.6576 0 -2.0 1e-06 
0.0 -0.6575 0 -2.0 1e-06 
0.0 -0.6574 0 -2.0 1e-06 
0.0 -0.6573 0 -2.0 1e-06 
0.0 -0.6572 0 -2.0 1e-06 
0.0 -0.6571 0 -2.0 1e-06 
0.0 -0.657 0 -2.0 1e-06 
0.0 -0.6569 0 -2.0 1e-06 
0.0 -0.6568 0 -2.0 1e-06 
0.0 -0.6567 0 -2.0 1e-06 
0.0 -0.6566 0 -2.0 1e-06 
0.0 -0.6565 0 -2.0 1e-06 
0.0 -0.6564 0 -2.0 1e-06 
0.0 -0.6563 0 -2.0 1e-06 
0.0 -0.6562 0 -2.0 1e-06 
0.0 -0.6561 0 -2.0 1e-06 
0.0 -0.656 0 -2.0 1e-06 
0.0 -0.6559 0 -2.0 1e-06 
0.0 -0.6558 0 -2.0 1e-06 
0.0 -0.6557 0 -2.0 1e-06 
0.0 -0.6556 0 -2.0 1e-06 
0.0 -0.6555 0 -2.0 1e-06 
0.0 -0.6554 0 -2.0 1e-06 
0.0 -0.6553 0 -2.0 1e-06 
0.0 -0.6552 0 -2.0 1e-06 
0.0 -0.6551 0 -2.0 1e-06 
0.0 -0.655 0 -2.0 1e-06 
0.0 -0.6549 0 -2.0 1e-06 
0.0 -0.6548 0 -2.0 1e-06 
0.0 -0.6547 0 -2.0 1e-06 
0.0 -0.6546 0 -2.0 1e-06 
0.0 -0.6545 0 -2.0 1e-06 
0.0 -0.6544 0 -2.0 1e-06 
0.0 -0.6543 0 -2.0 1e-06 
0.0 -0.6542 0 -2.0 1e-06 
0.0 -0.6541 0 -2.0 1e-06 
0.0 -0.654 0 -2.0 1e-06 
0.0 -0.6539 0 -2.0 1e-06 
0.0 -0.6538 0 -2.0 1e-06 
0.0 -0.6537 0 -2.0 1e-06 
0.0 -0.6536 0 -2.0 1e-06 
0.0 -0.6535 0 -2.0 1e-06 
0.0 -0.6534 0 -2.0 1e-06 
0.0 -0.6533 0 -2.0 1e-06 
0.0 -0.6532 0 -2.0 1e-06 
0.0 -0.6531 0 -2.0 1e-06 
0.0 -0.653 0 -2.0 1e-06 
0.0 -0.6529 0 -2.0 1e-06 
0.0 -0.6528 0 -2.0 1e-06 
0.0 -0.6527 0 -2.0 1e-06 
0.0 -0.6526 0 -2.0 1e-06 
0.0 -0.6525 0 -2.0 1e-06 
0.0 -0.6524 0 -2.0 1e-06 
0.0 -0.6523 0 -2.0 1e-06 
0.0 -0.6522 0 -2.0 1e-06 
0.0 -0.6521 0 -2.0 1e-06 
0.0 -0.652 0 -2.0 1e-06 
0.0 -0.6519 0 -2.0 1e-06 
0.0 -0.6518 0 -2.0 1e-06 
0.0 -0.6517 0 -2.0 1e-06 
0.0 -0.6516 0 -2.0 1e-06 
0.0 -0.6515 0 -2.0 1e-06 
0.0 -0.6514 0 -2.0 1e-06 
0.0 -0.6513 0 -2.0 1e-06 
0.0 -0.6512 0 -2.0 1e-06 
0.0 -0.6511 0 -2.0 1e-06 
0.0 -0.651 0 -2.0 1e-06 
0.0 -0.6509 0 -2.0 1e-06 
0.0 -0.6508 0 -2.0 1e-06 
0.0 -0.6507 0 -2.0 1e-06 
0.0 -0.6506 0 -2.0 1e-06 
0.0 -0.6505 0 -2.0 1e-06 
0.0 -0.6504 0 -2.0 1e-06 
0.0 -0.6503 0 -2.0 1e-06 
0.0 -0.6502 0 -2.0 1e-06 
0.0 -0.6501 0 -2.0 1e-06 
0.0 -0.65 0 -2.0 1e-06 
0.0 -0.6499 0 -2.0 1e-06 
0.0 -0.6498 0 -2.0 1e-06 
0.0 -0.6497 0 -2.0 1e-06 
0.0 -0.6496 0 -2.0 1e-06 
0.0 -0.6495 0 -2.0 1e-06 
0.0 -0.6494 0 -2.0 1e-06 
0.0 -0.6493 0 -2.0 1e-06 
0.0 -0.6492 0 -2.0 1e-06 
0.0 -0.6491 0 -2.0 1e-06 
0.0 -0.649 0 -2.0 1e-06 
0.0 -0.6489 0 -2.0 1e-06 
0.0 -0.6488 0 -2.0 1e-06 
0.0 -0.6487 0 -2.0 1e-06 
0.0 -0.6486 0 -2.0 1e-06 
0.0 -0.6485 0 -2.0 1e-06 
0.0 -0.6484 0 -2.0 1e-06 
0.0 -0.6483 0 -2.0 1e-06 
0.0 -0.6482 0 -2.0 1e-06 
0.0 -0.6481 0 -2.0 1e-06 
0.0 -0.648 0 -2.0 1e-06 
0.0 -0.6479 0 -2.0 1e-06 
0.0 -0.6478 0 -2.0 1e-06 
0.0 -0.6477 0 -2.0 1e-06 
0.0 -0.6476 0 -2.0 1e-06 
0.0 -0.6475 0 -2.0 1e-06 
0.0 -0.6474 0 -2.0 1e-06 
0.0 -0.6473 0 -2.0 1e-06 
0.0 -0.6472 0 -2.0 1e-06 
0.0 -0.6471 0 -2.0 1e-06 
0.0 -0.647 0 -2.0 1e-06 
0.0 -0.6469 0 -2.0 1e-06 
0.0 -0.6468 0 -2.0 1e-06 
0.0 -0.6467 0 -2.0 1e-06 
0.0 -0.6466 0 -2.0 1e-06 
0.0 -0.6465 0 -2.0 1e-06 
0.0 -0.6464 0 -2.0 1e-06 
0.0 -0.6463 0 -2.0 1e-06 
0.0 -0.6462 0 -2.0 1e-06 
0.0 -0.6461 0 -2.0 1e-06 
0.0 -0.646 0 -2.0 1e-06 
0.0 -0.6459 0 -2.0 1e-06 
0.0 -0.6458 0 -2.0 1e-06 
0.0 -0.6457 0 -2.0 1e-06 
0.0 -0.6456 0 -2.0 1e-06 
0.0 -0.6455 0 -2.0 1e-06 
0.0 -0.6454 0 -2.0 1e-06 
0.0 -0.6453 0 -2.0 1e-06 
0.0 -0.6452 0 -2.0 1e-06 
0.0 -0.6451 0 -2.0 1e-06 
0.0 -0.645 0 -2.0 1e-06 
0.0 -0.6449 0 -2.0 1e-06 
0.0 -0.6448 0 -2.0 1e-06 
0.0 -0.6447 0 -2.0 1e-06 
0.0 -0.6446 0 -2.0 1e-06 
0.0 -0.6445 0 -2.0 1e-06 
0.0 -0.6444 0 -2.0 1e-06 
0.0 -0.6443 0 -2.0 1e-06 
0.0 -0.6442 0 -2.0 1e-06 
0.0 -0.6441 0 -2.0 1e-06 
0.0 -0.644 0 -2.0 1e-06 
0.0 -0.6439 0 -2.0 1e-06 
0.0 -0.6438 0 -2.0 1e-06 
0.0 -0.6437 0 -2.0 1e-06 
0.0 -0.6436 0 -2.0 1e-06 
0.0 -0.6435 0 -2.0 1e-06 
0.0 -0.6434 0 -2.0 1e-06 
0.0 -0.6433 0 -2.0 1e-06 
0.0 -0.6432 0 -2.0 1e-06 
0.0 -0.6431 0 -2.0 1e-06 
0.0 -0.643 0 -2.0 1e-06 
0.0 -0.6429 0 -2.0 1e-06 
0.0 -0.6428 0 -2.0 1e-06 
0.0 -0.6427 0 -2.0 1e-06 
0.0 -0.6426 0 -2.0 1e-06 
0.0 -0.6425 0 -2.0 1e-06 
0.0 -0.6424 0 -2.0 1e-06 
0.0 -0.6423 0 -2.0 1e-06 
0.0 -0.6422 0 -2.0 1e-06 
0.0 -0.6421 0 -2.0 1e-06 
0.0 -0.642 0 -2.0 1e-06 
0.0 -0.6419 0 -2.0 1e-06 
0.0 -0.6418 0 -2.0 1e-06 
0.0 -0.6417 0 -2.0 1e-06 
0.0 -0.6416 0 -2.0 1e-06 
0.0 -0.6415 0 -2.0 1e-06 
0.0 -0.6414 0 -2.0 1e-06 
0.0 -0.6413 0 -2.0 1e-06 
0.0 -0.6412 0 -2.0 1e-06 
0.0 -0.6411 0 -2.0 1e-06 
0.0 -0.641 0 -2.0 1e-06 
0.0 -0.6409 0 -2.0 1e-06 
0.0 -0.6408 0 -2.0 1e-06 
0.0 -0.6407 0 -2.0 1e-06 
0.0 -0.6406 0 -2.0 1e-06 
0.0 -0.6405 0 -2.0 1e-06 
0.0 -0.6404 0 -2.0 1e-06 
0.0 -0.6403 0 -2.0 1e-06 
0.0 -0.6402 0 -2.0 1e-06 
0.0 -0.6401 0 -2.0 1e-06 
0.0 -0.64 0 -2.0 1e-06 
0.0 -0.6399 0 -2.0 1e-06 
0.0 -0.6398 0 -2.0 1e-06 
0.0 -0.6397 0 -2.0 1e-06 
0.0 -0.6396 0 -2.0 1e-06 
0.0 -0.6395 0 -2.0 1e-06 
0.0 -0.6394 0 -2.0 1e-06 
0.0 -0.6393 0 -2.0 1e-06 
0.0 -0.6392 0 -2.0 1e-06 
0.0 -0.6391 0 -2.0 1e-06 
0.0 -0.639 0 -2.0 1e-06 
0.0 -0.6389 0 -2.0 1e-06 
0.0 -0.6388 0 -2.0 1e-06 
0.0 -0.6387 0 -2.0 1e-06 
0.0 -0.6386 0 -2.0 1e-06 
0.0 -0.6385 0 -2.0 1e-06 
0.0 -0.6384 0 -2.0 1e-06 
0.0 -0.6383 0 -2.0 1e-06 
0.0 -0.6382 0 -2.0 1e-06 
0.0 -0.6381 0 -2.0 1e-06 
0.0 -0.638 0 -2.0 1e-06 
0.0 -0.6379 0 -2.0 1e-06 
0.0 -0.6378 0 -2.0 1e-06 
0.0 -0.6377 0 -2.0 1e-06 
0.0 -0.6376 0 -2.0 1e-06 
0.0 -0.6375 0 -2.0 1e-06 
0.0 -0.6374 0 -2.0 1e-06 
0.0 -0.6373 0 -2.0 1e-06 
0.0 -0.6372 0 -2.0 1e-06 
0.0 -0.6371 0 -2.0 1e-06 
0.0 -0.637 0 -2.0 1e-06 
0.0 -0.6369 0 -2.0 1e-06 
0.0 -0.6368 0 -2.0 1e-06 
0.0 -0.6367 0 -2.0 1e-06 
0.0 -0.6366 0 -2.0 1e-06 
0.0 -0.6365 0 -2.0 1e-06 
0.0 -0.6364 0 -2.0 1e-06 
0.0 -0.6363 0 -2.0 1e-06 
0.0 -0.6362 0 -2.0 1e-06 
0.0 -0.6361 0 -2.0 1e-06 
0.0 -0.636 0 -2.0 1e-06 
0.0 -0.6359 0 -2.0 1e-06 
0.0 -0.6358 0 -2.0 1e-06 
0.0 -0.6357 0 -2.0 1e-06 
0.0 -0.6356 0 -2.0 1e-06 
0.0 -0.6355 0 -2.0 1e-06 
0.0 -0.6354 0 -2.0 1e-06 
0.0 -0.6353 0 -2.0 1e-06 
0.0 -0.6352 0 -2.0 1e-06 
0.0 -0.6351 0 -2.0 1e-06 
0.0 -0.635 0 -2.0 1e-06 
0.0 -0.6349 0 -2.0 1e-06 
0.0 -0.6348 0 -2.0 1e-06 
0.0 -0.6347 0 -2.0 1e-06 
0.0 -0.6346 0 -2.0 1e-06 
0.0 -0.6345 0 -2.0 1e-06 
0.0 -0.6344 0 -2.0 1e-06 
0.0 -0.6343 0 -2.0 1e-06 
0.0 -0.6342 0 -2.0 1e-06 
0.0 -0.6341 0 -2.0 1e-06 
0.0 -0.634 0 -2.0 1e-06 
0.0 -0.6339 0 -2.0 1e-06 
0.0 -0.6338 0 -2.0 1e-06 
0.0 -0.6337 0 -2.0 1e-06 
0.0 -0.6336 0 -2.0 1e-06 
0.0 -0.6335 0 -2.0 1e-06 
0.0 -0.6334 0 -2.0 1e-06 
0.0 -0.6333 0 -2.0 1e-06 
0.0 -0.6332 0 -2.0 1e-06 
0.0 -0.6331 0 -2.0 1e-06 
0.0 -0.633 0 -2.0 1e-06 
0.0 -0.6329 0 -2.0 1e-06 
0.0 -0.6328 0 -2.0 1e-06 
0.0 -0.6327 0 -2.0 1e-06 
0.0 -0.6326 0 -2.0 1e-06 
0.0 -0.6325 0 -2.0 1e-06 
0.0 -0.6324 0 -2.0 1e-06 
0.0 -0.6323 0 -2.0 1e-06 
0.0 -0.6322 0 -2.0 1e-06 
0.0 -0.6321 0 -2.0 1e-06 
0.0 -0.632 0 -2.0 1e-06 
0.0 -0.6319 0 -2.0 1e-06 
0.0 -0.6318 0 -2.0 1e-06 
0.0 -0.6317 0 -2.0 1e-06 
0.0 -0.6316 0 -2.0 1e-06 
0.0 -0.6315 0 -2.0 1e-06 
0.0 -0.6314 0 -2.0 1e-06 
0.0 -0.6313 0 -2.0 1e-06 
0.0 -0.6312 0 -2.0 1e-06 
0.0 -0.6311 0 -2.0 1e-06 
0.0 -0.631 0 -2.0 1e-06 
0.0 -0.6309 0 -2.0 1e-06 
0.0 -0.6308 0 -2.0 1e-06 
0.0 -0.6307 0 -2.0 1e-06 
0.0 -0.6306 0 -2.0 1e-06 
0.0 -0.6305 0 -2.0 1e-06 
0.0 -0.6304 0 -2.0 1e-06 
0.0 -0.6303 0 -2.0 1e-06 
0.0 -0.6302 0 -2.0 1e-06 
0.0 -0.6301 0 -2.0 1e-06 
0.0 -0.63 0 -2.0 1e-06 
0.0 -0.6299 0 -2.0 1e-06 
0.0 -0.6298 0 -2.0 1e-06 
0.0 -0.6297 0 -2.0 1e-06 
0.0 -0.6296 0 -2.0 1e-06 
0.0 -0.6295 0 -2.0 1e-06 
0.0 -0.6294 0 -2.0 1e-06 
0.0 -0.6293 0 -2.0 1e-06 
0.0 -0.6292 0 -2.0 1e-06 
0.0 -0.6291 0 -2.0 1e-06 
0.0 -0.629 0 -2.0 1e-06 
0.0 -0.6289 0 -2.0 1e-06 
0.0 -0.6288 0 -2.0 1e-06 
0.0 -0.6287 0 -2.0 1e-06 
0.0 -0.6286 0 -2.0 1e-06 
0.0 -0.6285 0 -2.0 1e-06 
0.0 -0.6284 0 -2.0 1e-06 
0.0 -0.6283 0 -2.0 1e-06 
0.0 -0.6282 0 -2.0 1e-06 
0.0 -0.6281 0 -2.0 1e-06 
0.0 -0.628 0 -2.0 1e-06 
0.0 -0.6279 0 -2.0 1e-06 
0.0 -0.6278 0 -2.0 1e-06 
0.0 -0.6277 0 -2.0 1e-06 
0.0 -0.6276 0 -2.0 1e-06 
0.0 -0.6275 0 -2.0 1e-06 
0.0 -0.6274 0 -2.0 1e-06 
0.0 -0.6273 0 -2.0 1e-06 
0.0 -0.6272 0 -2.0 1e-06 
0.0 -0.6271 0 -2.0 1e-06 
0.0 -0.627 0 -2.0 1e-06 
0.0 -0.6269 0 -2.0 1e-06 
0.0 -0.6268 0 -2.0 1e-06 
0.0 -0.6267 0 -2.0 1e-06 
0.0 -0.6266 0 -2.0 1e-06 
0.0 -0.6265 0 -2.0 1e-06 
0.0 -0.6264 0 -2.0 1e-06 
0.0 -0.6263 0 -2.0 1e-06 
0.0 -0.6262 0 -2.0 1e-06 
0.0 -0.6261 0 -2.0 1e-06 
0.0 -0.626 0 -2.0 1e-06 
0.0 -0.6259 0 -2.0 1e-06 
0.0 -0.6258 0 -2.0 1e-06 
0.0 -0.6257 0 -2.0 1e-06 
0.0 -0.6256 0 -2.0 1e-06 
0.0 -0.6255 0 -2.0 1e-06 
0.0 -0.6254 0 -2.0 1e-06 
0.0 -0.6253 0 -2.0 1e-06 
0.0 -0.6252 0 -2.0 1e-06 
0.0 -0.6251 0 -2.0 1e-06 
0.0 -0.625 0 -2.0 1e-06 
0.0 -0.6249 0 -2.0 1e-06 
0.0 -0.6248 0 -2.0 1e-06 
0.0 -0.6247 0 -2.0 1e-06 
0.0 -0.6246 0 -2.0 1e-06 
0.0 -0.6245 0 -2.0 1e-06 
0.0 -0.6244 0 -2.0 1e-06 
0.0 -0.6243 0 -2.0 1e-06 
0.0 -0.6242 0 -2.0 1e-06 
0.0 -0.6241 0 -2.0 1e-06 
0.0 -0.624 0 -2.0 1e-06 
0.0 -0.6239 0 -2.0 1e-06 
0.0 -0.6238 0 -2.0 1e-06 
0.0 -0.6237 0 -2.0 1e-06 
0.0 -0.6236 0 -2.0 1e-06 
0.0 -0.6235 0 -2.0 1e-06 
0.0 -0.6234 0 -2.0 1e-06 
0.0 -0.6233 0 -2.0 1e-06 
0.0 -0.6232 0 -2.0 1e-06 
0.0 -0.6231 0 -2.0 1e-06 
0.0 -0.623 0 -2.0 1e-06 
0.0 -0.6229 0 -2.0 1e-06 
0.0 -0.6228 0 -2.0 1e-06 
0.0 -0.6227 0 -2.0 1e-06 
0.0 -0.6226 0 -2.0 1e-06 
0.0 -0.6225 0 -2.0 1e-06 
0.0 -0.6224 0 -2.0 1e-06 
0.0 -0.6223 0 -2.0 1e-06 
0.0 -0.6222 0 -2.0 1e-06 
0.0 -0.6221 0 -2.0 1e-06 
0.0 -0.622 0 -2.0 1e-06 
0.0 -0.6219 0 -2.0 1e-06 
0.0 -0.6218 0 -2.0 1e-06 
0.0 -0.6217 0 -2.0 1e-06 
0.0 -0.6216 0 -2.0 1e-06 
0.0 -0.6215 0 -2.0 1e-06 
0.0 -0.6214 0 -2.0 1e-06 
0.0 -0.6213 0 -2.0 1e-06 
0.0 -0.6212 0 -2.0 1e-06 
0.0 -0.6211 0 -2.0 1e-06 
0.0 -0.621 0 -2.0 1e-06 
0.0 -0.6209 0 -2.0 1e-06 
0.0 -0.6208 0 -2.0 1e-06 
0.0 -0.6207 0 -2.0 1e-06 
0.0 -0.6206 0 -2.0 1e-06 
0.0 -0.6205 0 -2.0 1e-06 
0.0 -0.6204 0 -2.0 1e-06 
0.0 -0.6203 0 -2.0 1e-06 
0.0 -0.6202 0 -2.0 1e-06 
0.0 -0.6201 0 -2.0 1e-06 
0.0 -0.62 0 -2.0 1e-06 
0.0 -0.6199 0 -2.0 1e-06 
0.0 -0.6198 0 -2.0 1e-06 
0.0 -0.6197 0 -2.0 1e-06 
0.0 -0.6196 0 -2.0 1e-06 
0.0 -0.6195 0 -2.0 1e-06 
0.0 -0.6194 0 -2.0 1e-06 
0.0 -0.6193 0 -2.0 1e-06 
0.0 -0.6192 0 -2.0 1e-06 
0.0 -0.6191 0 -2.0 1e-06 
0.0 -0.619 0 -2.0 1e-06 
0.0 -0.6189 0 -2.0 1e-06 
0.0 -0.6188 0 -2.0 1e-06 
0.0 -0.6187 0 -2.0 1e-06 
0.0 -0.6186 0 -2.0 1e-06 
0.0 -0.6185 0 -2.0 1e-06 
0.0 -0.6184 0 -2.0 1e-06 
0.0 -0.6183 0 -2.0 1e-06 
0.0 -0.6182 0 -2.0 1e-06 
0.0 -0.6181 0 -2.0 1e-06 
0.0 -0.618 0 -2.0 1e-06 
0.0 -0.6179 0 -2.0 1e-06 
0.0 -0.6178 0 -2.0 1e-06 
0.0 -0.6177 0 -2.0 1e-06 
0.0 -0.6176 0 -2.0 1e-06 
0.0 -0.6175 0 -2.0 1e-06 
0.0 -0.6174 0 -2.0 1e-06 
0.0 -0.6173 0 -2.0 1e-06 
0.0 -0.6172 0 -2.0 1e-06 
0.0 -0.6171 0 -2.0 1e-06 
0.0 -0.617 0 -2.0 1e-06 
0.0 -0.6169 0 -2.0 1e-06 
0.0 -0.6168 0 -2.0 1e-06 
0.0 -0.6167 0 -2.0 1e-06 
0.0 -0.6166 0 -2.0 1e-06 
0.0 -0.6165 0 -2.0 1e-06 
0.0 -0.6164 0 -2.0 1e-06 
0.0 -0.6163 0 -2.0 1e-06 
0.0 -0.6162 0 -2.0 1e-06 
0.0 -0.6161 0 -2.0 1e-06 
0.0 -0.616 0 -2.0 1e-06 
0.0 -0.6159 0 -2.0 1e-06 
0.0 -0.6158 0 -2.0 1e-06 
0.0 -0.6157 0 -2.0 1e-06 
0.0 -0.6156 0 -2.0 1e-06 
0.0 -0.6155 0 -2.0 1e-06 
0.0 -0.6154 0 -2.0 1e-06 
0.0 -0.6153 0 -2.0 1e-06 
0.0 -0.6152 0 -2.0 1e-06 
0.0 -0.6151 0 -2.0 1e-06 
0.0 -0.615 0 -2.0 1e-06 
0.0 -0.6149 0 -2.0 1e-06 
0.0 -0.6148 0 -2.0 1e-06 
0.0 -0.6147 0 -2.0 1e-06 
0.0 -0.6146 0 -2.0 1e-06 
0.0 -0.6145 0 -2.0 1e-06 
0.0 -0.6144 0 -2.0 1e-06 
0.0 -0.6143 0 -2.0 1e-06 
0.0 -0.6142 0 -2.0 1e-06 
0.0 -0.6141 0 -2.0 1e-06 
0.0 -0.614 0 -2.0 1e-06 
0.0 -0.6139 0 -2.0 1e-06 
0.0 -0.6138 0 -2.0 1e-06 
0.0 -0.6137 0 -2.0 1e-06 
0.0 -0.6136 0 -2.0 1e-06 
0.0 -0.6135 0 -2.0 1e-06 
0.0 -0.6134 0 -2.0 1e-06 
0.0 -0.6133 0 -2.0 1e-06 
0.0 -0.6132 0 -2.0 1e-06 
0.0 -0.6131 0 -2.0 1e-06 
0.0 -0.613 0 -2.0 1e-06 
0.0 -0.6129 0 -2.0 1e-06 
0.0 -0.6128 0 -2.0 1e-06 
0.0 -0.6127 0 -2.0 1e-06 
0.0 -0.6126 0 -2.0 1e-06 
0.0 -0.6125 0 -2.0 1e-06 
0.0 -0.6124 0 -2.0 1e-06 
0.0 -0.6123 0 -2.0 1e-06 
0.0 -0.6122 0 -2.0 1e-06 
0.0 -0.6121 0 -2.0 1e-06 
0.0 -0.612 0 -2.0 1e-06 
0.0 -0.6119 0 -2.0 1e-06 
0.0 -0.6118 0 -2.0 1e-06 
0.0 -0.6117 0 -2.0 1e-06 
0.0 -0.6116 0 -2.0 1e-06 
0.0 -0.6115 0 -2.0 1e-06 
0.0 -0.6114 0 -2.0 1e-06 
0.0 -0.6113 0 -2.0 1e-06 
0.0 -0.6112 0 -2.0 1e-06 
0.0 -0.6111 0 -2.0 1e-06 
0.0 -0.611 0 -2.0 1e-06 
0.0 -0.6109 0 -2.0 1e-06 
0.0 -0.6108 0 -2.0 1e-06 
0.0 -0.6107 0 -2.0 1e-06 
0.0 -0.6106 0 -2.0 1e-06 
0.0 -0.6105 0 -2.0 1e-06 
0.0 -0.6104 0 -2.0 1e-06 
0.0 -0.6103 0 -2.0 1e-06 
0.0 -0.6102 0 -2.0 1e-06 
0.0 -0.6101 0 -2.0 1e-06 
0.0 -0.61 0 -2.0 1e-06 
0.0 -0.6099 0 -2.0 1e-06 
0.0 -0.6098 0 -2.0 1e-06 
0.0 -0.6097 0 -2.0 1e-06 
0.0 -0.6096 0 -2.0 1e-06 
0.0 -0.6095 0 -2.0 1e-06 
0.0 -0.6094 0 -2.0 1e-06 
0.0 -0.6093 0 -2.0 1e-06 
0.0 -0.6092 0 -2.0 1e-06 
0.0 -0.6091 0 -2.0 1e-06 
0.0 -0.609 0 -2.0 1e-06 
0.0 -0.6089 0 -2.0 1e-06 
0.0 -0.6088 0 -2.0 1e-06 
0.0 -0.6087 0 -2.0 1e-06 
0.0 -0.6086 0 -2.0 1e-06 
0.0 -0.6085 0 -2.0 1e-06 
0.0 -0.6084 0 -2.0 1e-06 
0.0 -0.6083 0 -2.0 1e-06 
0.0 -0.6082 0 -2.0 1e-06 
0.0 -0.6081 0 -2.0 1e-06 
0.0 -0.608 0 -2.0 1e-06 
0.0 -0.6079 0 -2.0 1e-06 
0.0 -0.6078 0 -2.0 1e-06 
0.0 -0.6077 0 -2.0 1e-06 
0.0 -0.6076 0 -2.0 1e-06 
0.0 -0.6075 0 -2.0 1e-06 
0.0 -0.6074 0 -2.0 1e-06 
0.0 -0.6073 0 -2.0 1e-06 
0.0 -0.6072 0 -2.0 1e-06 
0.0 -0.6071 0 -2.0 1e-06 
0.0 -0.607 0 -2.0 1e-06 
0.0 -0.6069 0 -2.0 1e-06 
0.0 -0.6068 0 -2.0 1e-06 
0.0 -0.6067 0 -2.0 1e-06 
0.0 -0.6066 0 -2.0 1e-06 
0.0 -0.6065 0 -2.0 1e-06 
0.0 -0.6064 0 -2.0 1e-06 
0.0 -0.6063 0 -2.0 1e-06 
0.0 -0.6062 0 -2.0 1e-06 
0.0 -0.6061 0 -2.0 1e-06 
0.0 -0.606 0 -2.0 1e-06 
0.0 -0.6059 0 -2.0 1e-06 
0.0 -0.6058 0 -2.0 1e-06 
0.0 -0.6057 0 -2.0 1e-06 
0.0 -0.6056 0 -2.0 1e-06 
0.0 -0.6055 0 -2.0 1e-06 
0.0 -0.6054 0 -2.0 1e-06 
0.0 -0.6053 0 -2.0 1e-06 
0.0 -0.6052 0 -2.0 1e-06 
0.0 -0.6051 0 -2.0 1e-06 
0.0 -0.605 0 -2.0 1e-06 
0.0 -0.6049 0 -2.0 1e-06 
0.0 -0.6048 0 -2.0 1e-06 
0.0 -0.6047 0 -2.0 1e-06 
0.0 -0.6046 0 -2.0 1e-06 
0.0 -0.6045 0 -2.0 1e-06 
0.0 -0.6044 0 -2.0 1e-06 
0.0 -0.6043 0 -2.0 1e-06 
0.0 -0.6042 0 -2.0 1e-06 
0.0 -0.6041 0 -2.0 1e-06 
0.0 -0.604 0 -2.0 1e-06 
0.0 -0.6039 0 -2.0 1e-06 
0.0 -0.6038 0 -2.0 1e-06 
0.0 -0.6037 0 -2.0 1e-06 
0.0 -0.6036 0 -2.0 1e-06 
0.0 -0.6035 0 -2.0 1e-06 
0.0 -0.6034 0 -2.0 1e-06 
0.0 -0.6033 0 -2.0 1e-06 
0.0 -0.6032 0 -2.0 1e-06 
0.0 -0.6031 0 -2.0 1e-06 
0.0 -0.603 0 -2.0 1e-06 
0.0 -0.6029 0 -2.0 1e-06 
0.0 -0.6028 0 -2.0 1e-06 
0.0 -0.6027 0 -2.0 1e-06 
0.0 -0.6026 0 -2.0 1e-06 
0.0 -0.6025 0 -2.0 1e-06 
0.0 -0.6024 0 -2.0 1e-06 
0.0 -0.6023 0 -2.0 1e-06 
0.0 -0.6022 0 -2.0 1e-06 
0.0 -0.6021 0 -2.0 1e-06 
0.0 -0.602 0 -2.0 1e-06 
0.0 -0.6019 0 -2.0 1e-06 
0.0 -0.6018 0 -2.0 1e-06 
0.0 -0.6017 0 -2.0 1e-06 
0.0 -0.6016 0 -2.0 1e-06 
0.0 -0.6015 0 -2.0 1e-06 
0.0 -0.6014 0 -2.0 1e-06 
0.0 -0.6013 0 -2.0 1e-06 
0.0 -0.6012 0 -2.0 1e-06 
0.0 -0.6011 0 -2.0 1e-06 
0.0 -0.601 0 -2.0 1e-06 
0.0 -0.6009 0 -2.0 1e-06 
0.0 -0.6008 0 -2.0 1e-06 
0.0 -0.6007 0 -2.0 1e-06 
0.0 -0.6006 0 -2.0 1e-06 
0.0 -0.6005 0 -2.0 1e-06 
0.0 -0.6004 0 -2.0 1e-06 
0.0 -0.6003 0 -2.0 1e-06 
0.0 -0.6002 0 -2.0 1e-06 
0.0 -0.6001 0 -2.0 1e-06 
0.0 -0.6 0 -2.0 1e-06 
0.0 -0.5999 0 -2.0 1e-06 
0.0 -0.5998 0 -2.0 1e-06 
0.0 -0.5997 0 -2.0 1e-06 
0.0 -0.5996 0 -2.0 1e-06 
0.0 -0.5995 0 -2.0 1e-06 
0.0 -0.5994 0 -2.0 1e-06 
0.0 -0.5993 0 -2.0 1e-06 
0.0 -0.5992 0 -2.0 1e-06 
0.0 -0.5991 0 -2.0 1e-06 
0.0 -0.599 0 -2.0 1e-06 
0.0 -0.5989 0 -2.0 1e-06 
0.0 -0.5988 0 -2.0 1e-06 
0.0 -0.5987 0 -2.0 1e-06 
0.0 -0.5986 0 -2.0 1e-06 
0.0 -0.5985 0 -2.0 1e-06 
0.0 -0.5984 0 -2.0 1e-06 
0.0 -0.5983 0 -2.0 1e-06 
0.0 -0.5982 0 -2.0 1e-06 
0.0 -0.5981 0 -2.0 1e-06 
0.0 -0.598 0 -2.0 1e-06 
0.0 -0.5979 0 -2.0 1e-06 
0.0 -0.5978 0 -2.0 1e-06 
0.0 -0.5977 0 -2.0 1e-06 
0.0 -0.5976 0 -2.0 1e-06 
0.0 -0.5975 0 -2.0 1e-06 
0.0 -0.5974 0 -2.0 1e-06 
0.0 -0.5973 0 -2.0 1e-06 
0.0 -0.5972 0 -2.0 1e-06 
0.0 -0.5971 0 -2.0 1e-06 
0.0 -0.597 0 -2.0 1e-06 
0.0 -0.5969 0 -2.0 1e-06 
0.0 -0.5968 0 -2.0 1e-06 
0.0 -0.5967 0 -2.0 1e-06 
0.0 -0.5966 0 -2.0 1e-06 
0.0 -0.5965 0 -2.0 1e-06 
0.0 -0.5964 0 -2.0 1e-06 
0.0 -0.5963 0 -2.0 1e-06 
0.0 -0.5962 0 -2.0 1e-06 
0.0 -0.5961 0 -2.0 1e-06 
0.0 -0.596 0 -2.0 1e-06 
0.0 -0.5959 0 -2.0 1e-06 
0.0 -0.5958 0 -2.0 1e-06 
0.0 -0.5957 0 -2.0 1e-06 
0.0 -0.5956 0 -2.0 1e-06 
0.0 -0.5955 0 -2.0 1e-06 
0.0 -0.5954 0 -2.0 1e-06 
0.0 -0.5953 0 -2.0 1e-06 
0.0 -0.5952 0 -2.0 1e-06 
0.0 -0.5951 0 -2.0 1e-06 
0.0 -0.595 0 -2.0 1e-06 
0.0 -0.5949 0 -2.0 1e-06 
0.0 -0.5948 0 -2.0 1e-06 
0.0 -0.5947 0 -2.0 1e-06 
0.0 -0.5946 0 -2.0 1e-06 
0.0 -0.5945 0 -2.0 1e-06 
0.0 -0.5944 0 -2.0 1e-06 
0.0 -0.5943 0 -2.0 1e-06 
0.0 -0.5942 0 -2.0 1e-06 
0.0 -0.5941 0 -2.0 1e-06 
0.0 -0.594 0 -2.0 1e-06 
0.0 -0.5939 0 -2.0 1e-06 
0.0 -0.5938 0 -2.0 1e-06 
0.0 -0.5937 0 -2.0 1e-06 
0.0 -0.5936 0 -2.0 1e-06 
0.0 -0.5935 0 -2.0 1e-06 
0.0 -0.5934 0 -2.0 1e-06 
0.0 -0.5933 0 -2.0 1e-06 
0.0 -0.5932 0 -2.0 1e-06 
0.0 -0.5931 0 -2.0 1e-06 
0.0 -0.593 0 -2.0 1e-06 
0.0 -0.5929 0 -2.0 1e-06 
0.0 -0.5928 0 -2.0 1e-06 
0.0 -0.5927 0 -2.0 1e-06 
0.0 -0.5926 0 -2.0 1e-06 
0.0 -0.5925 0 -2.0 1e-06 
0.0 -0.5924 0 -2.0 1e-06 
0.0 -0.5923 0 -2.0 1e-06 
0.0 -0.5922 0 -2.0 1e-06 
0.0 -0.5921 0 -2.0 1e-06 
0.0 -0.592 0 -2.0 1e-06 
0.0 -0.5919 0 -2.0 1e-06 
0.0 -0.5918 0 -2.0 1e-06 
0.0 -0.5917 0 -2.0 1e-06 
0.0 -0.5916 0 -2.0 1e-06 
0.0 -0.5915 0 -2.0 1e-06 
0.0 -0.5914 0 -2.0 1e-06 
0.0 -0.5913 0 -2.0 1e-06 
0.0 -0.5912 0 -2.0 1e-06 
0.0 -0.5911 0 -2.0 1e-06 
0.0 -0.591 0 -2.0 1e-06 
0.0 -0.5909 0 -2.0 1e-06 
0.0 -0.5908 0 -2.0 1e-06 
0.0 -0.5907 0 -2.0 1e-06 
0.0 -0.5906 0 -2.0 1e-06 
0.0 -0.5905 0 -2.0 1e-06 
0.0 -0.5904 0 -2.0 1e-06 
0.0 -0.5903 0 -2.0 1e-06 
0.0 -0.5902 0 -2.0 1e-06 
0.0 -0.5901 0 -2.0 1e-06 
0.0 -0.59 0 -2.0 1e-06 
0.0 -0.5899 0 -2.0 1e-06 
0.0 -0.5898 0 -2.0 1e-06 
0.0 -0.5897 0 -2.0 1e-06 
0.0 -0.5896 0 -2.0 1e-06 
0.0 -0.5895 0 -2.0 1e-06 
0.0 -0.5894 0 -2.0 1e-06 
0.0 -0.5893 0 -2.0 1e-06 
0.0 -0.5892 0 -2.0 1e-06 
0.0 -0.5891 0 -2.0 1e-06 
0.0 -0.589 0 -2.0 1e-06 
0.0 -0.5889 0 -2.0 1e-06 
0.0 -0.5888 0 -2.0 1e-06 
0.0 -0.5887 0 -2.0 1e-06 
0.0 -0.5886 0 -2.0 1e-06 
0.0 -0.5885 0 -2.0 1e-06 
0.0 -0.5884 0 -2.0 1e-06 
0.0 -0.5883 0 -2.0 1e-06 
0.0 -0.5882 0 -2.0 1e-06 
0.0 -0.5881 0 -2.0 1e-06 
0.0 -0.588 0 -2.0 1e-06 
0.0 -0.5879 0 -2.0 1e-06 
0.0 -0.5878 0 -2.0 1e-06 
0.0 -0.5877 0 -2.0 1e-06 
0.0 -0.5876 0 -2.0 1e-06 
0.0 -0.5875 0 -2.0 1e-06 
0.0 -0.5874 0 -2.0 1e-06 
0.0 -0.5873 0 -2.0 1e-06 
0.0 -0.5872 0 -2.0 1e-06 
0.0 -0.5871 0 -2.0 1e-06 
0.0 -0.587 0 -2.0 1e-06 
0.0 -0.5869 0 -2.0 1e-06 
0.0 -0.5868 0 -2.0 1e-06 
0.0 -0.5867 0 -2.0 1e-06 
0.0 -0.5866 0 -2.0 1e-06 
0.0 -0.5865 0 -2.0 1e-06 
0.0 -0.5864 0 -2.0 1e-06 
0.0 -0.5863 0 -2.0 1e-06 
0.0 -0.5862 0 -2.0 1e-06 
0.0 -0.5861 0 -2.0 1e-06 
0.0 -0.586 0 -2.0 1e-06 
0.0 -0.5859 0 -2.0 1e-06 
0.0 -0.5858 0 -2.0 1e-06 
0.0 -0.5857 0 -2.0 1e-06 
0.0 -0.5856 0 -2.0 1e-06 
0.0 -0.5855 0 -2.0 1e-06 
0.0 -0.5854 0 -2.0 1e-06 
0.0 -0.5853 0 -2.0 1e-06 
0.0 -0.5852 0 -2.0 1e-06 
0.0 -0.5851 0 -2.0 1e-06 
0.0 -0.585 0 -2.0 1e-06 
0.0 -0.5849 0 -2.0 1e-06 
0.0 -0.5848 0 -2.0 1e-06 
0.0 -0.5847 0 -2.0 1e-06 
0.0 -0.5846 0 -2.0 1e-06 
0.0 -0.5845 0 -2.0 1e-06 
0.0 -0.5844 0 -2.0 1e-06 
0.0 -0.5843 0 -2.0 1e-06 
0.0 -0.5842 0 -2.0 1e-06 
0.0 -0.5841 0 -2.0 1e-06 
0.0 -0.584 0 -2.0 1e-06 
0.0 -0.5839 0 -2.0 1e-06 
0.0 -0.5838 0 -2.0 1e-06 
0.0 -0.5837 0 -2.0 1e-06 
0.0 -0.5836 0 -2.0 1e-06 
0.0 -0.5835 0 -2.0 1e-06 
0.0 -0.5834 0 -2.0 1e-06 
0.0 -0.5833 0 -2.0 1e-06 
0.0 -0.5832 0 -2.0 1e-06 
0.0 -0.5831 0 -2.0 1e-06 
0.0 -0.583 0 -2.0 1e-06 
0.0 -0.5829 0 -2.0 1e-06 
0.0 -0.5828 0 -2.0 1e-06 
0.0 -0.5827 0 -2.0 1e-06 
0.0 -0.5826 0 -2.0 1e-06 
0.0 -0.5825 0 -2.0 1e-06 
0.0 -0.5824 0 -2.0 1e-06 
0.0 -0.5823 0 -2.0 1e-06 
0.0 -0.5822 0 -2.0 1e-06 
0.0 -0.5821 0 -2.0 1e-06 
0.0 -0.582 0 -2.0 1e-06 
0.0 -0.5819 0 -2.0 1e-06 
0.0 -0.5818 0 -2.0 1e-06 
0.0 -0.5817 0 -2.0 1e-06 
0.0 -0.5816 0 -2.0 1e-06 
0.0 -0.5815 0 -2.0 1e-06 
0.0 -0.5814 0 -2.0 1e-06 
0.0 -0.5813 0 -2.0 1e-06 
0.0 -0.5812 0 -2.0 1e-06 
0.0 -0.5811 0 -2.0 1e-06 
0.0 -0.581 0 -2.0 1e-06 
0.0 -0.5809 0 -2.0 1e-06 
0.0 -0.5808 0 -2.0 1e-06 
0.0 -0.5807 0 -2.0 1e-06 
0.0 -0.5806 0 -2.0 1e-06 
0.0 -0.5805 0 -2.0 1e-06 
0.0 -0.5804 0 -2.0 1e-06 
0.0 -0.5803 0 -2.0 1e-06 
0.0 -0.5802 0 -2.0 1e-06 
0.0 -0.5801 0 -2.0 1e-06 
0.0 -0.58 0 -2.0 1e-06 
0.0 -0.5799 0 -2.0 1e-06 
0.0 -0.5798 0 -2.0 1e-06 
0.0 -0.5797 0 -2.0 1e-06 
0.0 -0.5796 0 -2.0 1e-06 
0.0 -0.5795 0 -2.0 1e-06 
0.0 -0.5794 0 -2.0 1e-06 
0.0 -0.5793 0 -2.0 1e-06 
0.0 -0.5792 0 -2.0 1e-06 
0.0 -0.5791 0 -2.0 1e-06 
0.0 -0.579 0 -2.0 1e-06 
0.0 -0.5789 0 -2.0 1e-06 
0.0 -0.5788 0 -2.0 1e-06 
0.0 -0.5787 0 -2.0 1e-06 
0.0 -0.5786 0 -2.0 1e-06 
0.0 -0.5785 0 -2.0 1e-06 
0.0 -0.5784 0 -2.0 1e-06 
0.0 -0.5783 0 -2.0 1e-06 
0.0 -0.5782 0 -2.0 1e-06 
0.0 -0.5781 0 -2.0 1e-06 
0.0 -0.578 0 -2.0 1e-06 
0.0 -0.5779 0 -2.0 1e-06 
0.0 -0.5778 0 -2.0 1e-06 
0.0 -0.5777 0 -2.0 1e-06 
0.0 -0.5776 0 -2.0 1e-06 
0.0 -0.5775 0 -2.0 1e-06 
0.0 -0.5774 0 -2.0 1e-06 
0.0 -0.5773 0 -2.0 1e-06 
0.0 -0.5772 0 -2.0 1e-06 
0.0 -0.5771 0 -2.0 1e-06 
0.0 -0.577 0 -2.0 1e-06 
0.0 -0.5769 0 -2.0 1e-06 
0.0 -0.5768 0 -2.0 1e-06 
0.0 -0.5767 0 -2.0 1e-06 
0.0 -0.5766 0 -2.0 1e-06 
0.0 -0.5765 0 -2.0 1e-06 
0.0 -0.5764 0 -2.0 1e-06 
0.0 -0.5763 0 -2.0 1e-06 
0.0 -0.5762 0 -2.0 1e-06 
0.0 -0.5761 0 -2.0 1e-06 
0.0 -0.576 0 -2.0 1e-06 
0.0 -0.5759 0 -2.0 1e-06 
0.0 -0.5758 0 -2.0 1e-06 
0.0 -0.5757 0 -2.0 1e-06 
0.0 -0.5756 0 -2.0 1e-06 
0.0 -0.5755 0 -2.0 1e-06 
0.0 -0.5754 0 -2.0 1e-06 
0.0 -0.5753 0 -2.0 1e-06 
0.0 -0.5752 0 -2.0 1e-06 
0.0 -0.5751 0 -2.0 1e-06 
0.0 -0.575 0 -2.0 1e-06 
0.0 -0.5749 0 -2.0 1e-06 
0.0 -0.5748 0 -2.0 1e-06 
0.0 -0.5747 0 -2.0 1e-06 
0.0 -0.5746 0 -2.0 1e-06 
0.0 -0.5745 0 -2.0 1e-06 
0.0 -0.5744 0 -2.0 1e-06 
0.0 -0.5743 0 -2.0 1e-06 
0.0 -0.5742 0 -2.0 1e-06 
0.0 -0.5741 0 -2.0 1e-06 
0.0 -0.574 0 -2.0 1e-06 
0.0 -0.5739 0 -2.0 1e-06 
0.0 -0.5738 0 -2.0 1e-06 
0.0 -0.5737 0 -2.0 1e-06 
0.0 -0.5736 0 -2.0 1e-06 
0.0 -0.5735 0 -2.0 1e-06 
0.0 -0.5734 0 -2.0 1e-06 
0.0 -0.5733 0 -2.0 1e-06 
0.0 -0.5732 0 -2.0 1e-06 
0.0 -0.5731 0 -2.0 1e-06 
0.0 -0.573 0 -2.0 1e-06 
0.0 -0.5729 0 -2.0 1e-06 
0.0 -0.5728 0 -2.0 1e-06 
0.0 -0.5727 0 -2.0 1e-06 
0.0 -0.5726 0 -2.0 1e-06 
0.0 -0.5725 0 -2.0 1e-06 
0.0 -0.5724 0 -2.0 1e-06 
0.0 -0.5723 0 -2.0 1e-06 
0.0 -0.5722 0 -2.0 1e-06 
0.0 -0.5721 0 -2.0 1e-06 
0.0 -0.572 0 -2.0 1e-06 
0.0 -0.5719 0 -2.0 1e-06 
0.0 -0.5718 0 -2.0 1e-06 
0.0 -0.5717 0 -2.0 1e-06 
0.0 -0.5716 0 -2.0 1e-06 
0.0 -0.5715 0 -2.0 1e-06 
0.0 -0.5714 0 -2.0 1e-06 
0.0 -0.5713 0 -2.0 1e-06 
0.0 -0.5712 0 -2.0 1e-06 
0.0 -0.5711 0 -2.0 1e-06 
0.0 -0.571 0 -2.0 1e-06 
0.0 -0.5709 0 -2.0 1e-06 
0.0 -0.5708 0 -2.0 1e-06 
0.0 -0.5707 0 -2.0 1e-06 
0.0 -0.5706 0 -2.0 1e-06 
0.0 -0.5705 0 -2.0 1e-06 
0.0 -0.5704 0 -2.0 1e-06 
0.0 -0.5703 0 -2.0 1e-06 
0.0 -0.5702 0 -2.0 1e-06 
0.0 -0.5701 0 -2.0 1e-06 
0.0 -0.57 0 -2.0 1e-06 
0.0 -0.5699 0 -2.0 1e-06 
0.0 -0.5698 0 -2.0 1e-06 
0.0 -0.5697 0 -2.0 1e-06 
0.0 -0.5696 0 -2.0 1e-06 
0.0 -0.5695 0 -2.0 1e-06 
0.0 -0.5694 0 -2.0 1e-06 
0.0 -0.5693 0 -2.0 1e-06 
0.0 -0.5692 0 -2.0 1e-06 
0.0 -0.5691 0 -2.0 1e-06 
0.0 -0.569 0 -2.0 1e-06 
0.0 -0.5689 0 -2.0 1e-06 
0.0 -0.5688 0 -2.0 1e-06 
0.0 -0.5687 0 -2.0 1e-06 
0.0 -0.5686 0 -2.0 1e-06 
0.0 -0.5685 0 -2.0 1e-06 
0.0 -0.5684 0 -2.0 1e-06 
0.0 -0.5683 0 -2.0 1e-06 
0.0 -0.5682 0 -2.0 1e-06 
0.0 -0.5681 0 -2.0 1e-06 
0.0 -0.568 0 -2.0 1e-06 
0.0 -0.5679 0 -2.0 1e-06 
0.0 -0.5678 0 -2.0 1e-06 
0.0 -0.5677 0 -2.0 1e-06 
0.0 -0.5676 0 -2.0 1e-06 
0.0 -0.5675 0 -2.0 1e-06 
0.0 -0.5674 0 -2.0 1e-06 
0.0 -0.5673 0 -2.0 1e-06 
0.0 -0.5672 0 -2.0 1e-06 
0.0 -0.5671 0 -2.0 1e-06 
0.0 -0.567 0 -2.0 1e-06 
0.0 -0.5669 0 -2.0 1e-06 
0.0 -0.5668 0 -2.0 1e-06 
0.0 -0.5667 0 -2.0 1e-06 
0.0 -0.5666 0 -2.0 1e-06 
0.0 -0.5665 0 -2.0 1e-06 
0.0 -0.5664 0 -2.0 1e-06 
0.0 -0.5663 0 -2.0 1e-06 
0.0 -0.5662 0 -2.0 1e-06 
0.0 -0.5661 0 -2.0 1e-06 
0.0 -0.566 0 -2.0 1e-06 
0.0 -0.5659 0 -2.0 1e-06 
0.0 -0.5658 0 -2.0 1e-06 
0.0 -0.5657 0 -2.0 1e-06 
0.0 -0.5656 0 -2.0 1e-06 
0.0 -0.5655 0 -2.0 1e-06 
0.0 -0.5654 0 -2.0 1e-06 
0.0 -0.5653 0 -2.0 1e-06 
0.0 -0.5652 0 -2.0 1e-06 
0.0 -0.5651 0 -2.0 1e-06 
0.0 -0.565 0 -2.0 1e-06 
0.0 -0.5649 0 -2.0 1e-06 
0.0 -0.5648 0 -2.0 1e-06 
0.0 -0.5647 0 -2.0 1e-06 
0.0 -0.5646 0 -2.0 1e-06 
0.0 -0.5645 0 -2.0 1e-06 
0.0 -0.5644 0 -2.0 1e-06 
0.0 -0.5643 0 -2.0 1e-06 
0.0 -0.5642 0 -2.0 1e-06 
0.0 -0.5641 0 -2.0 1e-06 
0.0 -0.564 0 -2.0 1e-06 
0.0 -0.5639 0 -2.0 1e-06 
0.0 -0.5638 0 -2.0 1e-06 
0.0 -0.5637 0 -2.0 1e-06 
0.0 -0.5636 0 -2.0 1e-06 
0.0 -0.5635 0 -2.0 1e-06 
0.0 -0.5634 0 -2.0 1e-06 
0.0 -0.5633 0 -2.0 1e-06 
0.0 -0.5632 0 -2.0 1e-06 
0.0 -0.5631 0 -2.0 1e-06 
0.0 -0.563 0 -2.0 1e-06 
0.0 -0.5629 0 -2.0 1e-06 
0.0 -0.5628 0 -2.0 1e-06 
0.0 -0.5627 0 -2.0 1e-06 
0.0 -0.5626 0 -2.0 1e-06 
0.0 -0.5625 0 -2.0 1e-06 
0.0 -0.5624 0 -2.0 1e-06 
0.0 -0.5623 0 -2.0 1e-06 
0.0 -0.5622 0 -2.0 1e-06 
0.0 -0.5621 0 -2.0 1e-06 
0.0 -0.562 0 -2.0 1e-06 
0.0 -0.5619 0 -2.0 1e-06 
0.0 -0.5618 0 -2.0 1e-06 
0.0 -0.5617 0 -2.0 1e-06 
0.0 -0.5616 0 -2.0 1e-06 
0.0 -0.5615 0 -2.0 1e-06 
0.0 -0.5614 0 -2.0 1e-06 
0.0 -0.5613 0 -2.0 1e-06 
0.0 -0.5612 0 -2.0 1e-06 
0.0 -0.5611 0 -2.0 1e-06 
0.0 -0.561 0 -2.0 1e-06 
0.0 -0.5609 0 -2.0 1e-06 
0.0 -0.5608 0 -2.0 1e-06 
0.0 -0.5607 0 -2.0 1e-06 
0.0 -0.5606 0 -2.0 1e-06 
0.0 -0.5605 0 -2.0 1e-06 
0.0 -0.5604 0 -2.0 1e-06 
0.0 -0.5603 0 -2.0 1e-06 
0.0 -0.5602 0 -2.0 1e-06 
0.0 -0.5601 0 -2.0 1e-06 
0.0 -0.56 0 -2.0 1e-06 
0.0 -0.5599 0 -2.0 1e-06 
0.0 -0.5598 0 -2.0 1e-06 
0.0 -0.5597 0 -2.0 1e-06 
0.0 -0.5596 0 -2.0 1e-06 
0.0 -0.5595 0 -2.0 1e-06 
0.0 -0.5594 0 -2.0 1e-06 
0.0 -0.5593 0 -2.0 1e-06 
0.0 -0.5592 0 -2.0 1e-06 
0.0 -0.5591 0 -2.0 1e-06 
0.0 -0.559 0 -2.0 1e-06 
0.0 -0.5589 0 -2.0 1e-06 
0.0 -0.5588 0 -2.0 1e-06 
0.0 -0.5587 0 -2.0 1e-06 
0.0 -0.5586 0 -2.0 1e-06 
0.0 -0.5585 0 -2.0 1e-06 
0.0 -0.5584 0 -2.0 1e-06 
0.0 -0.5583 0 -2.0 1e-06 
0.0 -0.5582 0 -2.0 1e-06 
0.0 -0.5581 0 -2.0 1e-06 
0.0 -0.558 0 -2.0 1e-06 
0.0 -0.5579 0 -2.0 1e-06 
0.0 -0.5578 0 -2.0 1e-06 
0.0 -0.5577 0 -2.0 1e-06 
0.0 -0.5576 0 -2.0 1e-06 
0.0 -0.5575 0 -2.0 1e-06 
0.0 -0.5574 0 -2.0 1e-06 
0.0 -0.5573 0 -2.0 1e-06 
0.0 -0.5572 0 -2.0 1e-06 
0.0 -0.5571 0 -2.0 1e-06 
0.0 -0.557 0 -2.0 1e-06 
0.0 -0.5569 0 -2.0 1e-06 
0.0 -0.5568 0 -2.0 1e-06 
0.0 -0.5567 0 -2.0 1e-06 
0.0 -0.5566 0 -2.0 1e-06 
0.0 -0.5565 0 -2.0 1e-06 
0.0 -0.5564 0 -2.0 1e-06 
0.0 -0.5563 0 -2.0 1e-06 
0.0 -0.5562 0 -2.0 1e-06 
0.0 -0.5561 0 -2.0 1e-06 
0.0 -0.556 0 -2.0 1e-06 
0.0 -0.5559 0 -2.0 1e-06 
0.0 -0.5558 0 -2.0 1e-06 
0.0 -0.5557 0 -2.0 1e-06 
0.0 -0.5556 0 -2.0 1e-06 
0.0 -0.5555 0 -2.0 1e-06 
0.0 -0.5554 0 -2.0 1e-06 
0.0 -0.5553 0 -2.0 1e-06 
0.0 -0.5552 0 -2.0 1e-06 
0.0 -0.5551 0 -2.0 1e-06 
0.0 -0.555 0 -2.0 1e-06 
0.0 -0.5549 0 -2.0 1e-06 
0.0 -0.5548 0 -2.0 1e-06 
0.0 -0.5547 0 -2.0 1e-06 
0.0 -0.5546 0 -2.0 1e-06 
0.0 -0.5545 0 -2.0 1e-06 
0.0 -0.5544 0 -2.0 1e-06 
0.0 -0.5543 0 -2.0 1e-06 
0.0 -0.5542 0 -2.0 1e-06 
0.0 -0.5541 0 -2.0 1e-06 
0.0 -0.554 0 -2.0 1e-06 
0.0 -0.5539 0 -2.0 1e-06 
0.0 -0.5538 0 -2.0 1e-06 
0.0 -0.5537 0 -2.0 1e-06 
0.0 -0.5536 0 -2.0 1e-06 
0.0 -0.5535 0 -2.0 1e-06 
0.0 -0.5534 0 -2.0 1e-06 
0.0 -0.5533 0 -2.0 1e-06 
0.0 -0.5532 0 -2.0 1e-06 
0.0 -0.5531 0 -2.0 1e-06 
0.0 -0.553 0 -2.0 1e-06 
0.0 -0.5529 0 -2.0 1e-06 
0.0 -0.5528 0 -2.0 1e-06 
0.0 -0.5527 0 -2.0 1e-06 
0.0 -0.5526 0 -2.0 1e-06 
0.0 -0.5525 0 -2.0 1e-06 
0.0 -0.5524 0 -2.0 1e-06 
0.0 -0.5523 0 -2.0 1e-06 
0.0 -0.5522 0 -2.0 1e-06 
0.0 -0.5521 0 -2.0 1e-06 
0.0 -0.552 0 -2.0 1e-06 
0.0 -0.5519 0 -2.0 1e-06 
0.0 -0.5518 0 -2.0 1e-06 
0.0 -0.5517 0 -2.0 1e-06 
0.0 -0.5516 0 -2.0 1e-06 
0.0 -0.5515 0 -2.0 1e-06 
0.0 -0.5514 0 -2.0 1e-06 
0.0 -0.5513 0 -2.0 1e-06 
0.0 -0.5512 0 -2.0 1e-06 
0.0 -0.5511 0 -2.0 1e-06 
0.0 -0.551 0 -2.0 1e-06 
0.0 -0.5509 0 -2.0 1e-06 
0.0 -0.5508 0 -2.0 1e-06 
0.0 -0.5507 0 -2.0 1e-06 
0.0 -0.5506 0 -2.0 1e-06 
0.0 -0.5505 0 -2.0 1e-06 
0.0 -0.5504 0 -2.0 1e-06 
0.0 -0.5503 0 -2.0 1e-06 
0.0 -0.5502 0 -2.0 1e-06 
0.0 -0.5501 0 -2.0 1e-06 
0.0 -0.55 0 -2.0 1e-06 
0.0 -0.5499 0 -2.0 1e-06 
0.0 -0.5498 0 -2.0 1e-06 
0.0 -0.5497 0 -2.0 1e-06 
0.0 -0.5496 0 -2.0 1e-06 
0.0 -0.5495 0 -2.0 1e-06 
0.0 -0.5494 0 -2.0 1e-06 
0.0 -0.5493 0 -2.0 1e-06 
0.0 -0.5492 0 -2.0 1e-06 
0.0 -0.5491 0 -2.0 1e-06 
0.0 -0.549 0 -2.0 1e-06 
0.0 -0.5489 0 -2.0 1e-06 
0.0 -0.5488 0 -2.0 1e-06 
0.0 -0.5487 0 -2.0 1e-06 
0.0 -0.5486 0 -2.0 1e-06 
0.0 -0.5485 0 -2.0 1e-06 
0.0 -0.5484 0 -2.0 1e-06 
0.0 -0.5483 0 -2.0 1e-06 
0.0 -0.5482 0 -2.0 1e-06 
0.0 -0.5481 0 -2.0 1e-06 
0.0 -0.548 0 -2.0 1e-06 
0.0 -0.5479 0 -2.0 1e-06 
0.0 -0.5478 0 -2.0 1e-06 
0.0 -0.5477 0 -2.0 1e-06 
0.0 -0.5476 0 -2.0 1e-06 
0.0 -0.5475 0 -2.0 1e-06 
0.0 -0.5474 0 -2.0 1e-06 
0.0 -0.5473 0 -2.0 1e-06 
0.0 -0.5472 0 -2.0 1e-06 
0.0 -0.5471 0 -2.0 1e-06 
0.0 -0.547 0 -2.0 1e-06 
0.0 -0.5469 0 -2.0 1e-06 
0.0 -0.5468 0 -2.0 1e-06 
0.0 -0.5467 0 -2.0 1e-06 
0.0 -0.5466 0 -2.0 1e-06 
0.0 -0.5465 0 -2.0 1e-06 
0.0 -0.5464 0 -2.0 1e-06 
0.0 -0.5463 0 -2.0 1e-06 
0.0 -0.5462 0 -2.0 1e-06 
0.0 -0.5461 0 -2.0 1e-06 
0.0 -0.546 0 -2.0 1e-06 
0.0 -0.5459 0 -2.0 1e-06 
0.0 -0.5458 0 -2.0 1e-06 
0.0 -0.5457 0 -2.0 1e-06 
0.0 -0.5456 0 -2.0 1e-06 
0.0 -0.5455 0 -2.0 1e-06 
0.0 -0.5454 0 -2.0 1e-06 
0.0 -0.5453 0 -2.0 1e-06 
0.0 -0.5452 0 -2.0 1e-06 
0.0 -0.5451 0 -2.0 1e-06 
0.0 -0.545 0 -2.0 1e-06 
0.0 -0.5449 0 -2.0 1e-06 
0.0 -0.5448 0 -2.0 1e-06 
0.0 -0.5447 0 -2.0 1e-06 
0.0 -0.5446 0 -2.0 1e-06 
0.0 -0.5445 0 -2.0 1e-06 
0.0 -0.5444 0 -2.0 1e-06 
0.0 -0.5443 0 -2.0 1e-06 
0.0 -0.5442 0 -2.0 1e-06 
0.0 -0.5441 0 -2.0 1e-06 
0.0 -0.544 0 -2.0 1e-06 
0.0 -0.5439 0 -2.0 1e-06 
0.0 -0.5438 0 -2.0 1e-06 
0.0 -0.5437 0 -2.0 1e-06 
0.0 -0.5436 0 -2.0 1e-06 
0.0 -0.5435 0 -2.0 1e-06 
0.0 -0.5434 0 -2.0 1e-06 
0.0 -0.5433 0 -2.0 1e-06 
0.0 -0.5432 0 -2.0 1e-06 
0.0 -0.5431 0 -2.0 1e-06 
0.0 -0.543 0 -2.0 1e-06 
0.0 -0.5429 0 -2.0 1e-06 
0.0 -0.5428 0 -2.0 1e-06 
0.0 -0.5427 0 -2.0 1e-06 
0.0 -0.5426 0 -2.0 1e-06 
0.0 -0.5425 0 -2.0 1e-06 
0.0 -0.5424 0 -2.0 1e-06 
0.0 -0.5423 0 -2.0 1e-06 
0.0 -0.5422 0 -2.0 1e-06 
0.0 -0.5421 0 -2.0 1e-06 
0.0 -0.542 0 -2.0 1e-06 
0.0 -0.5419 0 -2.0 1e-06 
0.0 -0.5418 0 -2.0 1e-06 
0.0 -0.5417 0 -2.0 1e-06 
0.0 -0.5416 0 -2.0 1e-06 
0.0 -0.5415 0 -2.0 1e-06 
0.0 -0.5414 0 -2.0 1e-06 
0.0 -0.5413 0 -2.0 1e-06 
0.0 -0.5412 0 -2.0 1e-06 
0.0 -0.5411 0 -2.0 1e-06 
0.0 -0.541 0 -2.0 1e-06 
0.0 -0.5409 0 -2.0 1e-06 
0.0 -0.5408 0 -2.0 1e-06 
0.0 -0.5407 0 -2.0 1e-06 
0.0 -0.5406 0 -2.0 1e-06 
0.0 -0.5405 0 -2.0 1e-06 
0.0 -0.5404 0 -2.0 1e-06 
0.0 -0.5403 0 -2.0 1e-06 
0.0 -0.5402 0 -2.0 1e-06 
0.0 -0.5401 0 -2.0 1e-06 
0.0 -0.54 0 -2.0 1e-06 
0.0 -0.5399 0 -2.0 1e-06 
0.0 -0.5398 0 -2.0 1e-06 
0.0 -0.5397 0 -2.0 1e-06 
0.0 -0.5396 0 -2.0 1e-06 
0.0 -0.5395 0 -2.0 1e-06 
0.0 -0.5394 0 -2.0 1e-06 
0.0 -0.5393 0 -2.0 1e-06 
0.0 -0.5392 0 -2.0 1e-06 
0.0 -0.5391 0 -2.0 1e-06 
0.0 -0.539 0 -2.0 1e-06 
0.0 -0.5389 0 -2.0 1e-06 
0.0 -0.5388 0 -2.0 1e-06 
0.0 -0.5387 0 -2.0 1e-06 
0.0 -0.5386 0 -2.0 1e-06 
0.0 -0.5385 0 -2.0 1e-06 
0.0 -0.5384 0 -2.0 1e-06 
0.0 -0.5383 0 -2.0 1e-06 
0.0 -0.5382 0 -2.0 1e-06 
0.0 -0.5381 0 -2.0 1e-06 
0.0 -0.538 0 -2.0 1e-06 
0.0 -0.5379 0 -2.0 1e-06 
0.0 -0.5378 0 -2.0 1e-06 
0.0 -0.5377 0 -2.0 1e-06 
0.0 -0.5376 0 -2.0 1e-06 
0.0 -0.5375 0 -2.0 1e-06 
0.0 -0.5374 0 -2.0 1e-06 
0.0 -0.5373 0 -2.0 1e-06 
0.0 -0.5372 0 -2.0 1e-06 
0.0 -0.5371 0 -2.0 1e-06 
0.0 -0.537 0 -2.0 1e-06 
0.0 -0.5369 0 -2.0 1e-06 
0.0 -0.5368 0 -2.0 1e-06 
0.0 -0.5367 0 -2.0 1e-06 
0.0 -0.5366 0 -2.0 1e-06 
0.0 -0.5365 0 -2.0 1e-06 
0.0 -0.5364 0 -2.0 1e-06 
0.0 -0.5363 0 -2.0 1e-06 
0.0 -0.5362 0 -2.0 1e-06 
0.0 -0.5361 0 -2.0 1e-06 
0.0 -0.536 0 -2.0 1e-06 
0.0 -0.5359 0 -2.0 1e-06 
0.0 -0.5358 0 -2.0 1e-06 
0.0 -0.5357 0 -2.0 1e-06 
0.0 -0.5356 0 -2.0 1e-06 
0.0 -0.5355 0 -2.0 1e-06 
0.0 -0.5354 0 -2.0 1e-06 
0.0 -0.5353 0 -2.0 1e-06 
0.0 -0.5352 0 -2.0 1e-06 
0.0 -0.5351 0 -2.0 1e-06 
0.0 -0.535 0 -2.0 1e-06 
0.0 -0.5349 0 -2.0 1e-06 
0.0 -0.5348 0 -2.0 1e-06 
0.0 -0.5347 0 -2.0 1e-06 
0.0 -0.5346 0 -2.0 1e-06 
0.0 -0.5345 0 -2.0 1e-06 
0.0 -0.5344 0 -2.0 1e-06 
0.0 -0.5343 0 -2.0 1e-06 
0.0 -0.5342 0 -2.0 1e-06 
0.0 -0.5341 0 -2.0 1e-06 
0.0 -0.534 0 -2.0 1e-06 
0.0 -0.5339 0 -2.0 1e-06 
0.0 -0.5338 0 -2.0 1e-06 
0.0 -0.5337 0 -2.0 1e-06 
0.0 -0.5336 0 -2.0 1e-06 
0.0 -0.5335 0 -2.0 1e-06 
0.0 -0.5334 0 -2.0 1e-06 
0.0 -0.5333 0 -2.0 1e-06 
0.0 -0.5332 0 -2.0 1e-06 
0.0 -0.5331 0 -2.0 1e-06 
0.0 -0.533 0 -2.0 1e-06 
0.0 -0.5329 0 -2.0 1e-06 
0.0 -0.5328 0 -2.0 1e-06 
0.0 -0.5327 0 -2.0 1e-06 
0.0 -0.5326 0 -2.0 1e-06 
0.0 -0.5325 0 -2.0 1e-06 
0.0 -0.5324 0 -2.0 1e-06 
0.0 -0.5323 0 -2.0 1e-06 
0.0 -0.5322 0 -2.0 1e-06 
0.0 -0.5321 0 -2.0 1e-06 
0.0 -0.532 0 -2.0 1e-06 
0.0 -0.5319 0 -2.0 1e-06 
0.0 -0.5318 0 -2.0 1e-06 
0.0 -0.5317 0 -2.0 1e-06 
0.0 -0.5316 0 -2.0 1e-06 
0.0 -0.5315 0 -2.0 1e-06 
0.0 -0.5314 0 -2.0 1e-06 
0.0 -0.5313 0 -2.0 1e-06 
0.0 -0.5312 0 -2.0 1e-06 
0.0 -0.5311 0 -2.0 1e-06 
0.0 -0.531 0 -2.0 1e-06 
0.0 -0.5309 0 -2.0 1e-06 
0.0 -0.5308 0 -2.0 1e-06 
0.0 -0.5307 0 -2.0 1e-06 
0.0 -0.5306 0 -2.0 1e-06 
0.0 -0.5305 0 -2.0 1e-06 
0.0 -0.5304 0 -2.0 1e-06 
0.0 -0.5303 0 -2.0 1e-06 
0.0 -0.5302 0 -2.0 1e-06 
0.0 -0.5301 0 -2.0 1e-06 
0.0 -0.53 0 -2.0 1e-06 
0.0 -0.5299 0 -2.0 1e-06 
0.0 -0.5298 0 -2.0 1e-06 
0.0 -0.5297 0 -2.0 1e-06 
0.0 -0.5296 0 -2.0 1e-06 
0.0 -0.5295 0 -2.0 1e-06 
0.0 -0.5294 0 -2.0 1e-06 
0.0 -0.5293 0 -2.0 1e-06 
0.0 -0.5292 0 -2.0 1e-06 
0.0 -0.5291 0 -2.0 1e-06 
0.0 -0.529 0 -2.0 1e-06 
0.0 -0.5289 0 -2.0 1e-06 
0.0 -0.5288 0 -2.0 1e-06 
0.0 -0.5287 0 -2.0 1e-06 
0.0 -0.5286 0 -2.0 1e-06 
0.0 -0.5285 0 -2.0 1e-06 
0.0 -0.5284 0 -2.0 1e-06 
0.0 -0.5283 0 -2.0 1e-06 
0.0 -0.5282 0 -2.0 1e-06 
0.0 -0.5281 0 -2.0 1e-06 
0.0 -0.528 0 -2.0 1e-06 
0.0 -0.5279 0 -2.0 1e-06 
0.0 -0.5278 0 -2.0 1e-06 
0.0 -0.5277 0 -2.0 1e-06 
0.0 -0.5276 0 -2.0 1e-06 
0.0 -0.5275 0 -2.0 1e-06 
0.0 -0.5274 0 -2.0 1e-06 
0.0 -0.5273 0 -2.0 1e-06 
0.0 -0.5272 0 -2.0 1e-06 
0.0 -0.5271 0 -2.0 1e-06 
0.0 -0.527 0 -2.0 1e-06 
0.0 -0.5269 0 -2.0 1e-06 
0.0 -0.5268 0 -2.0 1e-06 
0.0 -0.5267 0 -2.0 1e-06 
0.0 -0.5266 0 -2.0 1e-06 
0.0 -0.5265 0 -2.0 1e-06 
0.0 -0.5264 0 -2.0 1e-06 
0.0 -0.5263 0 -2.0 1e-06 
0.0 -0.5262 0 -2.0 1e-06 
0.0 -0.5261 0 -2.0 1e-06 
0.0 -0.526 0 -2.0 1e-06 
0.0 -0.5259 0 -2.0 1e-06 
0.0 -0.5258 0 -2.0 1e-06 
0.0 -0.5257 0 -2.0 1e-06 
0.0 -0.5256 0 -2.0 1e-06 
0.0 -0.5255 0 -2.0 1e-06 
0.0 -0.5254 0 -2.0 1e-06 
0.0 -0.5253 0 -2.0 1e-06 
0.0 -0.5252 0 -2.0 1e-06 
0.0 -0.5251 0 -2.0 1e-06 
0.0 -0.525 0 -2.0 1e-06 
0.0 -0.5249 0 -2.0 1e-06 
0.0 -0.5248 0 -2.0 1e-06 
0.0 -0.5247 0 -2.0 1e-06 
0.0 -0.5246 0 -2.0 1e-06 
0.0 -0.5245 0 -2.0 1e-06 
0.0 -0.5244 0 -2.0 1e-06 
0.0 -0.5243 0 -2.0 1e-06 
0.0 -0.5242 0 -2.0 1e-06 
0.0 -0.5241 0 -2.0 1e-06 
0.0 -0.524 0 -2.0 1e-06 
0.0 -0.5239 0 -2.0 1e-06 
0.0 -0.5238 0 -2.0 1e-06 
0.0 -0.5237 0 -2.0 1e-06 
0.0 -0.5236 0 -2.0 1e-06 
0.0 -0.5235 0 -2.0 1e-06 
0.0 -0.5234 0 -2.0 1e-06 
0.0 -0.5233 0 -2.0 1e-06 
0.0 -0.5232 0 -2.0 1e-06 
0.0 -0.5231 0 -2.0 1e-06 
0.0 -0.523 0 -2.0 1e-06 
0.0 -0.5229 0 -2.0 1e-06 
0.0 -0.5228 0 -2.0 1e-06 
0.0 -0.5227 0 -2.0 1e-06 
0.0 -0.5226 0 -2.0 1e-06 
0.0 -0.5225 0 -2.0 1e-06 
0.0 -0.5224 0 -2.0 1e-06 
0.0 -0.5223 0 -2.0 1e-06 
0.0 -0.5222 0 -2.0 1e-06 
0.0 -0.5221 0 -2.0 1e-06 
0.0 -0.522 0 -2.0 1e-06 
0.0 -0.5219 0 -2.0 1e-06 
0.0 -0.5218 0 -2.0 1e-06 
0.0 -0.5217 0 -2.0 1e-06 
0.0 -0.5216 0 -2.0 1e-06 
0.0 -0.5215 0 -2.0 1e-06 
0.0 -0.5214 0 -2.0 1e-06 
0.0 -0.5213 0 -2.0 1e-06 
0.0 -0.5212 0 -2.0 1e-06 
0.0 -0.5211 0 -2.0 1e-06 
0.0 -0.521 0 -2.0 1e-06 
0.0 -0.5209 0 -2.0 1e-06 
0.0 -0.5208 0 -2.0 1e-06 
0.0 -0.5207 0 -2.0 1e-06 
0.0 -0.5206 0 -2.0 1e-06 
0.0 -0.5205 0 -2.0 1e-06 
0.0 -0.5204 0 -2.0 1e-06 
0.0 -0.5203 0 -2.0 1e-06 
0.0 -0.5202 0 -2.0 1e-06 
0.0 -0.5201 0 -2.0 1e-06 
0.0 -0.52 0 -2.0 1e-06 
0.0 -0.5199 0 -2.0 1e-06 
0.0 -0.5198 0 -2.0 1e-06 
0.0 -0.5197 0 -2.0 1e-06 
0.0 -0.5196 0 -2.0 1e-06 
0.0 -0.5195 0 -2.0 1e-06 
0.0 -0.5194 0 -2.0 1e-06 
0.0 -0.5193 0 -2.0 1e-06 
0.0 -0.5192 0 -2.0 1e-06 
0.0 -0.5191 0 -2.0 1e-06 
0.0 -0.519 0 -2.0 1e-06 
0.0 -0.5189 0 -2.0 1e-06 
0.0 -0.5188 0 -2.0 1e-06 
0.0 -0.5187 0 -2.0 1e-06 
0.0 -0.5186 0 -2.0 1e-06 
0.0 -0.5185 0 -2.0 1e-06 
0.0 -0.5184 0 -2.0 1e-06 
0.0 -0.5183 0 -2.0 1e-06 
0.0 -0.5182 0 -2.0 1e-06 
0.0 -0.5181 0 -2.0 1e-06 
0.0 -0.518 0 -2.0 1e-06 
0.0 -0.5179 0 -2.0 1e-06 
0.0 -0.5178 0 -2.0 1e-06 
0.0 -0.5177 0 -2.0 1e-06 
0.0 -0.5176 0 -2.0 1e-06 
0.0 -0.5175 0 -2.0 1e-06 
0.0 -0.5174 0 -2.0 1e-06 
0.0 -0.5173 0 -2.0 1e-06 
0.0 -0.5172 0 -2.0 1e-06 
0.0 -0.5171 0 -2.0 1e-06 
0.0 -0.517 0 -2.0 1e-06 
0.0 -0.5169 0 -2.0 1e-06 
0.0 -0.5168 0 -2.0 1e-06 
0.0 -0.5167 0 -2.0 1e-06 
0.0 -0.5166 0 -2.0 1e-06 
0.0 -0.5165 0 -2.0 1e-06 
0.0 -0.5164 0 -2.0 1e-06 
0.0 -0.5163 0 -2.0 1e-06 
0.0 -0.5162 0 -2.0 1e-06 
0.0 -0.5161 0 -2.0 1e-06 
0.0 -0.516 0 -2.0 1e-06 
0.0 -0.5159 0 -2.0 1e-06 
0.0 -0.5158 0 -2.0 1e-06 
0.0 -0.5157 0 -2.0 1e-06 
0.0 -0.5156 0 -2.0 1e-06 
0.0 -0.5155 0 -2.0 1e-06 
0.0 -0.5154 0 -2.0 1e-06 
0.0 -0.5153 0 -2.0 1e-06 
0.0 -0.5152 0 -2.0 1e-06 
0.0 -0.5151 0 -2.0 1e-06 
0.0 -0.515 0 -2.0 1e-06 
0.0 -0.5149 0 -2.0 1e-06 
0.0 -0.5148 0 -2.0 1e-06 
0.0 -0.5147 0 -2.0 1e-06 
0.0 -0.5146 0 -2.0 1e-06 
0.0 -0.5145 0 -2.0 1e-06 
0.0 -0.5144 0 -2.0 1e-06 
0.0 -0.5143 0 -2.0 1e-06 
0.0 -0.5142 0 -2.0 1e-06 
0.0 -0.5141 0 -2.0 1e-06 
0.0 -0.514 0 -2.0 1e-06 
0.0 -0.5139 0 -2.0 1e-06 
0.0 -0.5138 0 -2.0 1e-06 
0.0 -0.5137 0 -2.0 1e-06 
0.0 -0.5136 0 -2.0 1e-06 
0.0 -0.5135 0 -2.0 1e-06 
0.0 -0.5134 0 -2.0 1e-06 
0.0 -0.5133 0 -2.0 1e-06 
0.0 -0.5132 0 -2.0 1e-06 
0.0 -0.5131 0 -2.0 1e-06 
0.0 -0.513 0 -2.0 1e-06 
0.0 -0.5129 0 -2.0 1e-06 
0.0 -0.5128 0 -2.0 1e-06 
0.0 -0.5127 0 -2.0 1e-06 
0.0 -0.5126 0 -2.0 1e-06 
0.0 -0.5125 0 -2.0 1e-06 
0.0 -0.5124 0 -2.0 1e-06 
0.0 -0.5123 0 -2.0 1e-06 
0.0 -0.5122 0 -2.0 1e-06 
0.0 -0.5121 0 -2.0 1e-06 
0.0 -0.512 0 -2.0 1e-06 
0.0 -0.5119 0 -2.0 1e-06 
0.0 -0.5118 0 -2.0 1e-06 
0.0 -0.5117 0 -2.0 1e-06 
0.0 -0.5116 0 -2.0 1e-06 
0.0 -0.5115 0 -2.0 1e-06 
0.0 -0.5114 0 -2.0 1e-06 
0.0 -0.5113 0 -2.0 1e-06 
0.0 -0.5112 0 -2.0 1e-06 
0.0 -0.5111 0 -2.0 1e-06 
0.0 -0.511 0 -2.0 1e-06 
0.0 -0.5109 0 -2.0 1e-06 
0.0 -0.5108 0 -2.0 1e-06 
0.0 -0.5107 0 -2.0 1e-06 
0.0 -0.5106 0 -2.0 1e-06 
0.0 -0.5105 0 -2.0 1e-06 
0.0 -0.5104 0 -2.0 1e-06 
0.0 -0.5103 0 -2.0 1e-06 
0.0 -0.5102 0 -2.0 1e-06 
0.0 -0.5101 0 -2.0 1e-06 
0.0 -0.51 0 -2.0 1e-06 
0.0 -0.5099 0 -2.0 1e-06 
0.0 -0.5098 0 -2.0 1e-06 
0.0 -0.5097 0 -2.0 1e-06 
0.0 -0.5096 0 -2.0 1e-06 
0.0 -0.5095 0 -2.0 1e-06 
0.0 -0.5094 0 -2.0 1e-06 
0.0 -0.5093 0 -2.0 1e-06 
0.0 -0.5092 0 -2.0 1e-06 
0.0 -0.5091 0 -2.0 1e-06 
0.0 -0.509 0 -2.0 1e-06 
0.0 -0.5089 0 -2.0 1e-06 
0.0 -0.5088 0 -2.0 1e-06 
0.0 -0.5087 0 -2.0 1e-06 
0.0 -0.5086 0 -2.0 1e-06 
0.0 -0.5085 0 -2.0 1e-06 
0.0 -0.5084 0 -2.0 1e-06 
0.0 -0.5083 0 -2.0 1e-06 
0.0 -0.5082 0 -2.0 1e-06 
0.0 -0.5081 0 -2.0 1e-06 
0.0 -0.508 0 -2.0 1e-06 
0.0 -0.5079 0 -2.0 1e-06 
0.0 -0.5078 0 -2.0 1e-06 
0.0 -0.5077 0 -2.0 1e-06 
0.0 -0.5076 0 -2.0 1e-06 
0.0 -0.5075 0 -2.0 1e-06 
0.0 -0.5074 0 -2.0 1e-06 
0.0 -0.5073 0 -2.0 1e-06 
0.0 -0.5072 0 -2.0 1e-06 
0.0 -0.5071 0 -2.0 1e-06 
0.0 -0.507 0 -2.0 1e-06 
0.0 -0.5069 0 -2.0 1e-06 
0.0 -0.5068 0 -2.0 1e-06 
0.0 -0.5067 0 -2.0 1e-06 
0.0 -0.5066 0 -2.0 1e-06 
0.0 -0.5065 0 -2.0 1e-06 
0.0 -0.5064 0 -2.0 1e-06 
0.0 -0.5063 0 -2.0 1e-06 
0.0 -0.5062 0 -2.0 1e-06 
0.0 -0.5061 0 -2.0 1e-06 
0.0 -0.506 0 -2.0 1e-06 
0.0 -0.5059 0 -2.0 1e-06 
0.0 -0.5058 0 -2.0 1e-06 
0.0 -0.5057 0 -2.0 1e-06 
0.0 -0.5056 0 -2.0 1e-06 
0.0 -0.5055 0 -2.0 1e-06 
0.0 -0.5054 0 -2.0 1e-06 
0.0 -0.5053 0 -2.0 1e-06 
0.0 -0.5052 0 -2.0 1e-06 
0.0 -0.5051 0 -2.0 1e-06 
0.0 -0.505 0 -2.0 1e-06 
0.0 -0.5049 0 -2.0 1e-06 
0.0 -0.5048 0 -2.0 1e-06 
0.0 -0.5047 0 -2.0 1e-06 
0.0 -0.5046 0 -2.0 1e-06 
0.0 -0.5045 0 -2.0 1e-06 
0.0 -0.5044 0 -2.0 1e-06 
0.0 -0.5043 0 -2.0 1e-06 
0.0 -0.5042 0 -2.0 1e-06 
0.0 -0.5041 0 -2.0 1e-06 
0.0 -0.504 0 -2.0 1e-06 
0.0 -0.5039 0 -2.0 1e-06 
0.0 -0.5038 0 -2.0 1e-06 
0.0 -0.5037 0 -2.0 1e-06 
0.0 -0.5036 0 -2.0 1e-06 
0.0 -0.5035 0 -2.0 1e-06 
0.0 -0.5034 0 -2.0 1e-06 
0.0 -0.5033 0 -2.0 1e-06 
0.0 -0.5032 0 -2.0 1e-06 
0.0 -0.5031 0 -2.0 1e-06 
0.0 -0.503 0 -2.0 1e-06 
0.0 -0.5029 0 -2.0 1e-06 
0.0 -0.5028 0 -2.0 1e-06 
0.0 -0.5027 0 -2.0 1e-06 
0.0 -0.5026 0 -2.0 1e-06 
0.0 -0.5025 0 -2.0 1e-06 
0.0 -0.5024 0 -2.0 1e-06 
0.0 -0.5023 0 -2.0 1e-06 
0.0 -0.5022 0 -2.0 1e-06 
0.0 -0.5021 0 -2.0 1e-06 
0.0 -0.502 0 -2.0 1e-06 
0.0 -0.5019 0 -2.0 1e-06 
0.0 -0.5018 0 -2.0 1e-06 
0.0 -0.5017 0 -2.0 1e-06 
0.0 -0.5016 0 -2.0 1e-06 
0.0 -0.5015 0 -2.0 1e-06 
0.0 -0.5014 0 -2.0 1e-06 
0.0 -0.5013 0 -2.0 1e-06 
0.0 -0.5012 0 -2.0 1e-06 
0.0 -0.5011 0 -2.0 1e-06 
0.0 -0.501 0 -2.0 1e-06 
0.0 -0.5009 0 -2.0 1e-06 
0.0 -0.5008 0 -2.0 1e-06 
0.0 -0.5007 0 -2.0 1e-06 
0.0 -0.5006 0 -2.0 1e-06 
0.0 -0.5005 0 -2.0 1e-06 
0.0 -0.5004 0 -2.0 1e-06 
0.0 -0.5003 0 -2.0 1e-06 
0.0 -0.5002 0 -2.0 1e-06 
0.0 -0.5001 0 -2.0 1e-06 
0.0 -0.5 0 -2.0 1e-06 
0.0 -0.4999 0 -2.0 1e-06 
0.0 -0.4998 0 -2.0 1e-06 
0.0 -0.4997 0 -2.0 1e-06 
0.0 -0.4996 0 -2.0 1e-06 
0.0 -0.4995 0 -2.0 1e-06 
0.0 -0.4994 0 -2.0 1e-06 
0.0 -0.4993 0 -2.0 1e-06 
0.0 -0.4992 0 -2.0 1e-06 
0.0 -0.4991 0 -2.0 1e-06 
0.0 -0.499 0 -2.0 1e-06 
0.0 -0.4989 0 -2.0 1e-06 
0.0 -0.4988 0 -2.0 1e-06 
0.0 -0.4987 0 -2.0 1e-06 
0.0 -0.4986 0 -2.0 1e-06 
0.0 -0.4985 0 -2.0 1e-06 
0.0 -0.4984 0 -2.0 1e-06 
0.0 -0.4983 0 -2.0 1e-06 
0.0 -0.4982 0 -2.0 1e-06 
0.0 -0.4981 0 -2.0 1e-06 
0.0 -0.498 0 -2.0 1e-06 
0.0 -0.4979 0 -2.0 1e-06 
0.0 -0.4978 0 -2.0 1e-06 
0.0 -0.4977 0 -2.0 1e-06 
0.0 -0.4976 0 -2.0 1e-06 
0.0 -0.4975 0 -2.0 1e-06 
0.0 -0.4974 0 -2.0 1e-06 
0.0 -0.4973 0 -2.0 1e-06 
0.0 -0.4972 0 -2.0 1e-06 
0.0 -0.4971 0 -2.0 1e-06 
0.0 -0.497 0 -2.0 1e-06 
0.0 -0.4969 0 -2.0 1e-06 
0.0 -0.4968 0 -2.0 1e-06 
0.0 -0.4967 0 -2.0 1e-06 
0.0 -0.4966 0 -2.0 1e-06 
0.0 -0.4965 0 -2.0 1e-06 
0.0 -0.4964 0 -2.0 1e-06 
0.0 -0.4963 0 -2.0 1e-06 
0.0 -0.4962 0 -2.0 1e-06 
0.0 -0.4961 0 -2.0 1e-06 
0.0 -0.496 0 -2.0 1e-06 
0.0 -0.4959 0 -2.0 1e-06 
0.0 -0.4958 0 -2.0 1e-06 
0.0 -0.4957 0 -2.0 1e-06 
0.0 -0.4956 0 -2.0 1e-06 
0.0 -0.4955 0 -2.0 1e-06 
0.0 -0.4954 0 -2.0 1e-06 
0.0 -0.4953 0 -2.0 1e-06 
0.0 -0.4952 0 -2.0 1e-06 
0.0 -0.4951 0 -2.0 1e-06 
0.0 -0.495 0 -2.0 1e-06 
0.0 -0.4949 0 -2.0 1e-06 
0.0 -0.4948 0 -2.0 1e-06 
0.0 -0.4947 0 -2.0 1e-06 
0.0 -0.4946 0 -2.0 1e-06 
0.0 -0.4945 0 -2.0 1e-06 
0.0 -0.4944 0 -2.0 1e-06 
0.0 -0.4943 0 -2.0 1e-06 
0.0 -0.4942 0 -2.0 1e-06 
0.0 -0.4941 0 -2.0 1e-06 
0.0 -0.494 0 -2.0 1e-06 
0.0 -0.4939 0 -2.0 1e-06 
0.0 -0.4938 0 -2.0 1e-06 
0.0 -0.4937 0 -2.0 1e-06 
0.0 -0.4936 0 -2.0 1e-06 
0.0 -0.4935 0 -2.0 1e-06 
0.0 -0.4934 0 -2.0 1e-06 
0.0 -0.4933 0 -2.0 1e-06 
0.0 -0.4932 0 -2.0 1e-06 
0.0 -0.4931 0 -2.0 1e-06 
0.0 -0.493 0 -2.0 1e-06 
0.0 -0.4929 0 -2.0 1e-06 
0.0 -0.4928 0 -2.0 1e-06 
0.0 -0.4927 0 -2.0 1e-06 
0.0 -0.4926 0 -2.0 1e-06 
0.0 -0.4925 0 -2.0 1e-06 
0.0 -0.4924 0 -2.0 1e-06 
0.0 -0.4923 0 -2.0 1e-06 
0.0 -0.4922 0 -2.0 1e-06 
0.0 -0.4921 0 -2.0 1e-06 
0.0 -0.492 0 -2.0 1e-06 
0.0 -0.4919 0 -2.0 1e-06 
0.0 -0.4918 0 -2.0 1e-06 
0.0 -0.4917 0 -2.0 1e-06 
0.0 -0.4916 0 -2.0 1e-06 
0.0 -0.4915 0 -2.0 1e-06 
0.0 -0.4914 0 -2.0 1e-06 
0.0 -0.4913 0 -2.0 1e-06 
0.0 -0.4912 0 -2.0 1e-06 
0.0 -0.4911 0 -2.0 1e-06 
0.0 -0.491 0 -2.0 1e-06 
0.0 -0.4909 0 -2.0 1e-06 
0.0 -0.4908 0 -2.0 1e-06 
0.0 -0.4907 0 -2.0 1e-06 
0.0 -0.4906 0 -2.0 1e-06 
0.0 -0.4905 0 -2.0 1e-06 
0.0 -0.4904 0 -2.0 1e-06 
0.0 -0.4903 0 -2.0 1e-06 
0.0 -0.4902 0 -2.0 1e-06 
0.0 -0.4901 0 -2.0 1e-06 
0.0 -0.49 0 -2.0 1e-06 
0.0 -0.4899 0 -2.0 1e-06 
0.0 -0.4898 0 -2.0 1e-06 
0.0 -0.4897 0 -2.0 1e-06 
0.0 -0.4896 0 -2.0 1e-06 
0.0 -0.4895 0 -2.0 1e-06 
0.0 -0.4894 0 -2.0 1e-06 
0.0 -0.4893 0 -2.0 1e-06 
0.0 -0.4892 0 -2.0 1e-06 
0.0 -0.4891 0 -2.0 1e-06 
0.0 -0.489 0 -2.0 1e-06 
0.0 -0.4889 0 -2.0 1e-06 
0.0 -0.4888 0 -2.0 1e-06 
0.0 -0.4887 0 -2.0 1e-06 
0.0 -0.4886 0 -2.0 1e-06 
0.0 -0.4885 0 -2.0 1e-06 
0.0 -0.4884 0 -2.0 1e-06 
0.0 -0.4883 0 -2.0 1e-06 
0.0 -0.4882 0 -2.0 1e-06 
0.0 -0.4881 0 -2.0 1e-06 
0.0 -0.488 0 -2.0 1e-06 
0.0 -0.4879 0 -2.0 1e-06 
0.0 -0.4878 0 -2.0 1e-06 
0.0 -0.4877 0 -2.0 1e-06 
0.0 -0.4876 0 -2.0 1e-06 
0.0 -0.4875 0 -2.0 1e-06 
0.0 -0.4874 0 -2.0 1e-06 
0.0 -0.4873 0 -2.0 1e-06 
0.0 -0.4872 0 -2.0 1e-06 
0.0 -0.4871 0 -2.0 1e-06 
0.0 -0.487 0 -2.0 1e-06 
0.0 -0.4869 0 -2.0 1e-06 
0.0 -0.4868 0 -2.0 1e-06 
0.0 -0.4867 0 -2.0 1e-06 
0.0 -0.4866 0 -2.0 1e-06 
0.0 -0.4865 0 -2.0 1e-06 
0.0 -0.4864 0 -2.0 1e-06 
0.0 -0.4863 0 -2.0 1e-06 
0.0 -0.4862 0 -2.0 1e-06 
0.0 -0.4861 0 -2.0 1e-06 
0.0 -0.486 0 -2.0 1e-06 
0.0 -0.4859 0 -2.0 1e-06 
0.0 -0.4858 0 -2.0 1e-06 
0.0 -0.4857 0 -2.0 1e-06 
0.0 -0.4856 0 -2.0 1e-06 
0.0 -0.4855 0 -2.0 1e-06 
0.0 -0.4854 0 -2.0 1e-06 
0.0 -0.4853 0 -2.0 1e-06 
0.0 -0.4852 0 -2.0 1e-06 
0.0 -0.4851 0 -2.0 1e-06 
0.0 -0.485 0 -2.0 1e-06 
0.0 -0.4849 0 -2.0 1e-06 
0.0 -0.4848 0 -2.0 1e-06 
0.0 -0.4847 0 -2.0 1e-06 
0.0 -0.4846 0 -2.0 1e-06 
0.0 -0.4845 0 -2.0 1e-06 
0.0 -0.4844 0 -2.0 1e-06 
0.0 -0.4843 0 -2.0 1e-06 
0.0 -0.4842 0 -2.0 1e-06 
0.0 -0.4841 0 -2.0 1e-06 
0.0 -0.484 0 -2.0 1e-06 
0.0 -0.4839 0 -2.0 1e-06 
0.0 -0.4838 0 -2.0 1e-06 
0.0 -0.4837 0 -2.0 1e-06 
0.0 -0.4836 0 -2.0 1e-06 
0.0 -0.4835 0 -2.0 1e-06 
0.0 -0.4834 0 -2.0 1e-06 
0.0 -0.4833 0 -2.0 1e-06 
0.0 -0.4832 0 -2.0 1e-06 
0.0 -0.4831 0 -2.0 1e-06 
0.0 -0.483 0 -2.0 1e-06 
0.0 -0.4829 0 -2.0 1e-06 
0.0 -0.4828 0 -2.0 1e-06 
0.0 -0.4827 0 -2.0 1e-06 
0.0 -0.4826 0 -2.0 1e-06 
0.0 -0.4825 0 -2.0 1e-06 
0.0 -0.4824 0 -2.0 1e-06 
0.0 -0.4823 0 -2.0 1e-06 
0.0 -0.4822 0 -2.0 1e-06 
0.0 -0.4821 0 -2.0 1e-06 
0.0 -0.482 0 -2.0 1e-06 
0.0 -0.4819 0 -2.0 1e-06 
0.0 -0.4818 0 -2.0 1e-06 
0.0 -0.4817 0 -2.0 1e-06 
0.0 -0.4816 0 -2.0 1e-06 
0.0 -0.4815 0 -2.0 1e-06 
0.0 -0.4814 0 -2.0 1e-06 
0.0 -0.4813 0 -2.0 1e-06 
0.0 -0.4812 0 -2.0 1e-06 
0.0 -0.4811 0 -2.0 1e-06 
0.0 -0.481 0 -2.0 1e-06 
0.0 -0.4809 0 -2.0 1e-06 
0.0 -0.4808 0 -2.0 1e-06 
0.0 -0.4807 0 -2.0 1e-06 
0.0 -0.4806 0 -2.0 1e-06 
0.0 -0.4805 0 -2.0 1e-06 
0.0 -0.4804 0 -2.0 1e-06 
0.0 -0.4803 0 -2.0 1e-06 
0.0 -0.4802 0 -2.0 1e-06 
0.0 -0.4801 0 -2.0 1e-06 
0.0 -0.48 0 -2.0 1e-06 
0.0 -0.4799 0 -2.0 1e-06 
0.0 -0.4798 0 -2.0 1e-06 
0.0 -0.4797 0 -2.0 1e-06 
0.0 -0.4796 0 -2.0 1e-06 
0.0 -0.4795 0 -2.0 1e-06 
0.0 -0.4794 0 -2.0 1e-06 
0.0 -0.4793 0 -2.0 1e-06 
0.0 -0.4792 0 -2.0 1e-06 
0.0 -0.4791 0 -2.0 1e-06 
0.0 -0.479 0 -2.0 1e-06 
0.0 -0.4789 0 -2.0 1e-06 
0.0 -0.4788 0 -2.0 1e-06 
0.0 -0.4787 0 -2.0 1e-06 
0.0 -0.4786 0 -2.0 1e-06 
0.0 -0.4785 0 -2.0 1e-06 
0.0 -0.4784 0 -2.0 1e-06 
0.0 -0.4783 0 -2.0 1e-06 
0.0 -0.4782 0 -2.0 1e-06 
0.0 -0.4781 0 -2.0 1e-06 
0.0 -0.478 0 -2.0 1e-06 
0.0 -0.4779 0 -2.0 1e-06 
0.0 -0.4778 0 -2.0 1e-06 
0.0 -0.4777 0 -2.0 1e-06 
0.0 -0.4776 0 -2.0 1e-06 
0.0 -0.4775 0 -2.0 1e-06 
0.0 -0.4774 0 -2.0 1e-06 
0.0 -0.4773 0 -2.0 1e-06 
0.0 -0.4772 0 -2.0 1e-06 
0.0 -0.4771 0 -2.0 1e-06 
0.0 -0.477 0 -2.0 1e-06 
0.0 -0.4769 0 -2.0 1e-06 
0.0 -0.4768 0 -2.0 1e-06 
0.0 -0.4767 0 -2.0 1e-06 
0.0 -0.4766 0 -2.0 1e-06 
0.0 -0.4765 0 -2.0 1e-06 
0.0 -0.4764 0 -2.0 1e-06 
0.0 -0.4763 0 -2.0 1e-06 
0.0 -0.4762 0 -2.0 1e-06 
0.0 -0.4761 0 -2.0 1e-06 
0.0 -0.476 0 -2.0 1e-06 
0.0 -0.4759 0 -2.0 1e-06 
0.0 -0.4758 0 -2.0 1e-06 
0.0 -0.4757 0 -2.0 1e-06 
0.0 -0.4756 0 -2.0 1e-06 
0.0 -0.4755 0 -2.0 1e-06 
0.0 -0.4754 0 -2.0 1e-06 
0.0 -0.4753 0 -2.0 1e-06 
0.0 -0.4752 0 -2.0 1e-06 
0.0 -0.4751 0 -2.0 1e-06 
0.0 -0.475 0 -2.0 1e-06 
0.0 -0.4749 0 -2.0 1e-06 
0.0 -0.4748 0 -2.0 1e-06 
0.0 -0.4747 0 -2.0 1e-06 
0.0 -0.4746 0 -2.0 1e-06 
0.0 -0.4745 0 -2.0 1e-06 
0.0 -0.4744 0 -2.0 1e-06 
0.0 -0.4743 0 -2.0 1e-06 
0.0 -0.4742 0 -2.0 1e-06 
0.0 -0.4741 0 -2.0 1e-06 
0.0 -0.474 0 -2.0 1e-06 
0.0 -0.4739 0 -2.0 1e-06 
0.0 -0.4738 0 -2.0 1e-06 
0.0 -0.4737 0 -2.0 1e-06 
0.0 -0.4736 0 -2.0 1e-06 
0.0 -0.4735 0 -2.0 1e-06 
0.0 -0.4734 0 -2.0 1e-06 
0.0 -0.4733 0 -2.0 1e-06 
0.0 -0.4732 0 -2.0 1e-06 
0.0 -0.4731 0 -2.0 1e-06 
0.0 -0.473 0 -2.0 1e-06 
0.0 -0.4729 0 -2.0 1e-06 
0.0 -0.4728 0 -2.0 1e-06 
0.0 -0.4727 0 -2.0 1e-06 
0.0 -0.4726 0 -2.0 1e-06 
0.0 -0.4725 0 -2.0 1e-06 
0.0 -0.4724 0 -2.0 1e-06 
0.0 -0.4723 0 -2.0 1e-06 
0.0 -0.4722 0 -2.0 1e-06 
0.0 -0.4721 0 -2.0 1e-06 
0.0 -0.472 0 -2.0 1e-06 
0.0 -0.4719 0 -2.0 1e-06 
0.0 -0.4718 0 -2.0 1e-06 
0.0 -0.4717 0 -2.0 1e-06 
0.0 -0.4716 0 -2.0 1e-06 
0.0 -0.4715 0 -2.0 1e-06 
0.0 -0.4714 0 -2.0 1e-06 
0.0 -0.4713 0 -2.0 1e-06 
0.0 -0.4712 0 -2.0 1e-06 
0.0 -0.4711 0 -2.0 1e-06 
0.0 -0.471 0 -2.0 1e-06 
0.0 -0.4709 0 -2.0 1e-06 
0.0 -0.4708 0 -2.0 1e-06 
0.0 -0.4707 0 -2.0 1e-06 
0.0 -0.4706 0 -2.0 1e-06 
0.0 -0.4705 0 -2.0 1e-06 
0.0 -0.4704 0 -2.0 1e-06 
0.0 -0.4703 0 -2.0 1e-06 
0.0 -0.4702 0 -2.0 1e-06 
0.0 -0.4701 0 -2.0 1e-06 
0.0 -0.47 0 -2.0 1e-06 
0.0 -0.4699 0 -2.0 1e-06 
0.0 -0.4698 0 -2.0 1e-06 
0.0 -0.4697 0 -2.0 1e-06 
0.0 -0.4696 0 -2.0 1e-06 
0.0 -0.4695 0 -2.0 1e-06 
0.0 -0.4694 0 -2.0 1e-06 
0.0 -0.4693 0 -2.0 1e-06 
0.0 -0.4692 0 -2.0 1e-06 
0.0 -0.4691 0 -2.0 1e-06 
0.0 -0.469 0 -2.0 1e-06 
0.0 -0.4689 0 -2.0 1e-06 
0.0 -0.4688 0 -2.0 1e-06 
0.0 -0.4687 0 -2.0 1e-06 
0.0 -0.4686 0 -2.0 1e-06 
0.0 -0.4685 0 -2.0 1e-06 
0.0 -0.4684 0 -2.0 1e-06 
0.0 -0.4683 0 -2.0 1e-06 
0.0 -0.4682 0 -2.0 1e-06 
0.0 -0.4681 0 -2.0 1e-06 
0.0 -0.468 0 -2.0 1e-06 
0.0 -0.4679 0 -2.0 1e-06 
0.0 -0.4678 0 -2.0 1e-06 
0.0 -0.4677 0 -2.0 1e-06 
0.0 -0.4676 0 -2.0 1e-06 
0.0 -0.4675 0 -2.0 1e-06 
0.0 -0.4674 0 -2.0 1e-06 
0.0 -0.4673 0 -2.0 1e-06 
0.0 -0.4672 0 -2.0 1e-06 
0.0 -0.4671 0 -2.0 1e-06 
0.0 -0.467 0 -2.0 1e-06 
0.0 -0.4669 0 -2.0 1e-06 
0.0 -0.4668 0 -2.0 1e-06 
0.0 -0.4667 0 -2.0 1e-06 
0.0 -0.4666 0 -2.0 1e-06 
0.0 -0.4665 0 -2.0 1e-06 
0.0 -0.4664 0 -2.0 1e-06 
0.0 -0.4663 0 -2.0 1e-06 
0.0 -0.4662 0 -2.0 1e-06 
0.0 -0.4661 0 -2.0 1e-06 
0.0 -0.466 0 -2.0 1e-06 
0.0 -0.4659 0 -2.0 1e-06 
0.0 -0.4658 0 -2.0 1e-06 
0.0 -0.4657 0 -2.0 1e-06 
0.0 -0.4656 0 -2.0 1e-06 
0.0 -0.4655 0 -2.0 1e-06 
0.0 -0.4654 0 -2.0 1e-06 
0.0 -0.4653 0 -2.0 1e-06 
0.0 -0.4652 0 -2.0 1e-06 
0.0 -0.4651 0 -2.0 1e-06 
0.0 -0.465 0 -2.0 1e-06 
0.0 -0.4649 0 -2.0 1e-06 
0.0 -0.4648 0 -2.0 1e-06 
0.0 -0.4647 0 -2.0 1e-06 
0.0 -0.4646 0 -2.0 1e-06 
0.0 -0.4645 0 -2.0 1e-06 
0.0 -0.4644 0 -2.0 1e-06 
0.0 -0.4643 0 -2.0 1e-06 
0.0 -0.4642 0 -2.0 1e-06 
0.0 -0.4641 0 -2.0 1e-06 
0.0 -0.464 0 -2.0 1e-06 
0.0 -0.4639 0 -2.0 1e-06 
0.0 -0.4638 0 -2.0 1e-06 
0.0 -0.4637 0 -2.0 1e-06 
0.0 -0.4636 0 -2.0 1e-06 
0.0 -0.4635 0 -2.0 1e-06 
0.0 -0.4634 0 -2.0 1e-06 
0.0 -0.4633 0 -2.0 1e-06 
0.0 -0.4632 0 -2.0 1e-06 
0.0 -0.4631 0 -2.0 1e-06 
0.0 -0.463 0 -2.0 1e-06 
0.0 -0.4629 0 -2.0 1e-06 
0.0 -0.4628 0 -2.0 1e-06 
0.0 -0.4627 0 -2.0 1e-06 
0.0 -0.4626 0 -2.0 1e-06 
0.0 -0.4625 0 -2.0 1e-06 
0.0 -0.4624 0 -2.0 1e-06 
0.0 -0.4623 0 -2.0 1e-06 
0.0 -0.4622 0 -2.0 1e-06 
0.0 -0.4621 0 -2.0 1e-06 
0.0 -0.462 0 -2.0 1e-06 
0.0 -0.4619 0 -2.0 1e-06 
0.0 -0.4618 0 -2.0 1e-06 
0.0 -0.4617 0 -2.0 1e-06 
0.0 -0.4616 0 -2.0 1e-06 
0.0 -0.4615 0 -2.0 1e-06 
0.0 -0.4614 0 -2.0 1e-06 
0.0 -0.4613 0 -2.0 1e-06 
0.0 -0.4612 0 -2.0 1e-06 
0.0 -0.4611 0 -2.0 1e-06 
0.0 -0.461 0 -2.0 1e-06 
0.0 -0.4609 0 -2.0 1e-06 
0.0 -0.4608 0 -2.0 1e-06 
0.0 -0.4607 0 -2.0 1e-06 
0.0 -0.4606 0 -2.0 1e-06 
0.0 -0.4605 0 -2.0 1e-06 
0.0 -0.4604 0 -2.0 1e-06 
0.0 -0.4603 0 -2.0 1e-06 
0.0 -0.4602 0 -2.0 1e-06 
0.0 -0.4601 0 -2.0 1e-06 
0.0 -0.46 0 -2.0 1e-06 
0.0 -0.4599 0 -2.0 1e-06 
0.0 -0.4598 0 -2.0 1e-06 
0.0 -0.4597 0 -2.0 1e-06 
0.0 -0.4596 0 -2.0 1e-06 
0.0 -0.4595 0 -2.0 1e-06 
0.0 -0.4594 0 -2.0 1e-06 
0.0 -0.4593 0 -2.0 1e-06 
0.0 -0.4592 0 -2.0 1e-06 
0.0 -0.4591 0 -2.0 1e-06 
0.0 -0.459 0 -2.0 1e-06 
0.0 -0.4589 0 -2.0 1e-06 
0.0 -0.4588 0 -2.0 1e-06 
0.0 -0.4587 0 -2.0 1e-06 
0.0 -0.4586 0 -2.0 1e-06 
0.0 -0.4585 0 -2.0 1e-06 
0.0 -0.4584 0 -2.0 1e-06 
0.0 -0.4583 0 -2.0 1e-06 
0.0 -0.4582 0 -2.0 1e-06 
0.0 -0.4581 0 -2.0 1e-06 
0.0 -0.458 0 -2.0 1e-06 
0.0 -0.4579 0 -2.0 1e-06 
0.0 -0.4578 0 -2.0 1e-06 
0.0 -0.4577 0 -2.0 1e-06 
0.0 -0.4576 0 -2.0 1e-06 
0.0 -0.4575 0 -2.0 1e-06 
0.0 -0.4574 0 -2.0 1e-06 
0.0 -0.4573 0 -2.0 1e-06 
0.0 -0.4572 0 -2.0 1e-06 
0.0 -0.4571 0 -2.0 1e-06 
0.0 -0.457 0 -2.0 1e-06 
0.0 -0.4569 0 -2.0 1e-06 
0.0 -0.4568 0 -2.0 1e-06 
0.0 -0.4567 0 -2.0 1e-06 
0.0 -0.4566 0 -2.0 1e-06 
0.0 -0.4565 0 -2.0 1e-06 
0.0 -0.4564 0 -2.0 1e-06 
0.0 -0.4563 0 -2.0 1e-06 
0.0 -0.4562 0 -2.0 1e-06 
0.0 -0.4561 0 -2.0 1e-06 
0.0 -0.456 0 -2.0 1e-06 
0.0 -0.4559 0 -2.0 1e-06 
0.0 -0.4558 0 -2.0 1e-06 
0.0 -0.4557 0 -2.0 1e-06 
0.0 -0.4556 0 -2.0 1e-06 
0.0 -0.4555 0 -2.0 1e-06 
0.0 -0.4554 0 -2.0 1e-06 
0.0 -0.4553 0 -2.0 1e-06 
0.0 -0.4552 0 -2.0 1e-06 
0.0 -0.4551 0 -2.0 1e-06 
0.0 -0.455 0 -2.0 1e-06 
0.0 -0.4549 0 -2.0 1e-06 
0.0 -0.4548 0 -2.0 1e-06 
0.0 -0.4547 0 -2.0 1e-06 
0.0 -0.4546 0 -2.0 1e-06 
0.0 -0.4545 0 -2.0 1e-06 
0.0 -0.4544 0 -2.0 1e-06 
0.0 -0.4543 0 -2.0 1e-06 
0.0 -0.4542 0 -2.0 1e-06 
0.0 -0.4541 0 -2.0 1e-06 
0.0 -0.454 0 -2.0 1e-06 
0.0 -0.4539 0 -2.0 1e-06 
0.0 -0.4538 0 -2.0 1e-06 
0.0 -0.4537 0 -2.0 1e-06 
0.0 -0.4536 0 -2.0 1e-06 
0.0 -0.4535 0 -2.0 1e-06 
0.0 -0.4534 0 -2.0 1e-06 
0.0 -0.4533 0 -2.0 1e-06 
0.0 -0.4532 0 -2.0 1e-06 
0.0 -0.4531 0 -2.0 1e-06 
0.0 -0.453 0 -2.0 1e-06 
0.0 -0.4529 0 -2.0 1e-06 
0.0 -0.4528 0 -2.0 1e-06 
0.0 -0.4527 0 -2.0 1e-06 
0.0 -0.4526 0 -2.0 1e-06 
0.0 -0.4525 0 -2.0 1e-06 
0.0 -0.4524 0 -2.0 1e-06 
0.0 -0.4523 0 -2.0 1e-06 
0.0 -0.4522 0 -2.0 1e-06 
0.0 -0.4521 0 -2.0 1e-06 
0.0 -0.452 0 -2.0 1e-06 
0.0 -0.4519 0 -2.0 1e-06 
0.0 -0.4518 0 -2.0 1e-06 
0.0 -0.4517 0 -2.0 1e-06 
0.0 -0.4516 0 -2.0 1e-06 
0.0 -0.4515 0 -2.0 1e-06 
0.0 -0.4514 0 -2.0 1e-06 
0.0 -0.4513 0 -2.0 1e-06 
0.0 -0.4512 0 -2.0 1e-06 
0.0 -0.4511 0 -2.0 1e-06 
0.0 -0.451 0 -2.0 1e-06 
0.0 -0.4509 0 -2.0 1e-06 
0.0 -0.4508 0 -2.0 1e-06 
0.0 -0.4507 0 -2.0 1e-06 
0.0 -0.4506 0 -2.0 1e-06 
0.0 -0.4505 0 -2.0 1e-06 
0.0 -0.4504 0 -2.0 1e-06 
0.0 -0.4503 0 -2.0 1e-06 
0.0 -0.4502 0 -2.0 1e-06 
0.0 -0.4501 0 -2.0 1e-06 
0.0 -0.45 0 -2.0 1e-06 
0.0 -0.4499 0 -2.0 1e-06 
0.0 -0.4498 0 -2.0 1e-06 
0.0 -0.4497 0 -2.0 1e-06 
0.0 -0.4496 0 -2.0 1e-06 
0.0 -0.4495 0 -2.0 1e-06 
0.0 -0.4494 0 -2.0 1e-06 
0.0 -0.4493 0 -2.0 1e-06 
0.0 -0.4492 0 -2.0 1e-06 
0.0 -0.4491 0 -2.0 1e-06 
0.0 -0.449 0 -2.0 1e-06 
0.0 -0.4489 0 -2.0 1e-06 
0.0 -0.4488 0 -2.0 1e-06 
0.0 -0.4487 0 -2.0 1e-06 
0.0 -0.4486 0 -2.0 1e-06 
0.0 -0.4485 0 -2.0 1e-06 
0.0 -0.4484 0 -2.0 1e-06 
0.0 -0.4483 0 -2.0 1e-06 
0.0 -0.4482 0 -2.0 1e-06 
0.0 -0.4481 0 -2.0 1e-06 
0.0 -0.448 0 -2.0 1e-06 
0.0 -0.4479 0 -2.0 1e-06 
0.0 -0.4478 0 -2.0 1e-06 
0.0 -0.4477 0 -2.0 1e-06 
0.0 -0.4476 0 -2.0 1e-06 
0.0 -0.4475 0 -2.0 1e-06 
0.0 -0.4474 0 -2.0 1e-06 
0.0 -0.4473 0 -2.0 1e-06 
0.0 -0.4472 0 -2.0 1e-06 
0.0 -0.4471 0 -2.0 1e-06 
0.0 -0.447 0 -2.0 1e-06 
0.0 -0.4469 0 -2.0 1e-06 
0.0 -0.4468 0 -2.0 1e-06 
0.0 -0.4467 0 -2.0 1e-06 
0.0 -0.4466 0 -2.0 1e-06 
0.0 -0.4465 0 -2.0 1e-06 
0.0 -0.4464 0 -2.0 1e-06 
0.0 -0.4463 0 -2.0 1e-06 
0.0 -0.4462 0 -2.0 1e-06 
0.0 -0.4461 0 -2.0 1e-06 
0.0 -0.446 0 -2.0 1e-06 
0.0 -0.4459 0 -2.0 1e-06 
0.0 -0.4458 0 -2.0 1e-06 
0.0 -0.4457 0 -2.0 1e-06 
0.0 -0.4456 0 -2.0 1e-06 
0.0 -0.4455 0 -2.0 1e-06 
0.0 -0.4454 0 -2.0 1e-06 
0.0 -0.4453 0 -2.0 1e-06 
0.0 -0.4452 0 -2.0 1e-06 
0.0 -0.4451 0 -2.0 1e-06 
0.0 -0.445 0 -2.0 1e-06 
0.0 -0.4449 0 -2.0 1e-06 
0.0 -0.4448 0 -2.0 1e-06 
0.0 -0.4447 0 -2.0 1e-06 
0.0 -0.4446 0 -2.0 1e-06 
0.0 -0.4445 0 -2.0 1e-06 
0.0 -0.4444 0 -2.0 1e-06 
0.0 -0.4443 0 -2.0 1e-06 
0.0 -0.4442 0 -2.0 1e-06 
0.0 -0.4441 0 -2.0 1e-06 
0.0 -0.444 0 -2.0 1e-06 
0.0 -0.4439 0 -2.0 1e-06 
0.0 -0.4438 0 -2.0 1e-06 
0.0 -0.4437 0 -2.0 1e-06 
0.0 -0.4436 0 -2.0 1e-06 
0.0 -0.4435 0 -2.0 1e-06 
0.0 -0.4434 0 -2.0 1e-06 
0.0 -0.4433 0 -2.0 1e-06 
0.0 -0.4432 0 -2.0 1e-06 
0.0 -0.4431 0 -2.0 1e-06 
0.0 -0.443 0 -2.0 1e-06 
0.0 -0.4429 0 -2.0 1e-06 
0.0 -0.4428 0 -2.0 1e-06 
0.0 -0.4427 0 -2.0 1e-06 
0.0 -0.4426 0 -2.0 1e-06 
0.0 -0.4425 0 -2.0 1e-06 
0.0 -0.4424 0 -2.0 1e-06 
0.0 -0.4423 0 -2.0 1e-06 
0.0 -0.4422 0 -2.0 1e-06 
0.0 -0.4421 0 -2.0 1e-06 
0.0 -0.442 0 -2.0 1e-06 
0.0 -0.4419 0 -2.0 1e-06 
0.0 -0.4418 0 -2.0 1e-06 
0.0 -0.4417 0 -2.0 1e-06 
0.0 -0.4416 0 -2.0 1e-06 
0.0 -0.4415 0 -2.0 1e-06 
0.0 -0.4414 0 -2.0 1e-06 
0.0 -0.4413 0 -2.0 1e-06 
0.0 -0.4412 0 -2.0 1e-06 
0.0 -0.4411 0 -2.0 1e-06 
0.0 -0.441 0 -2.0 1e-06 
0.0 -0.4409 0 -2.0 1e-06 
0.0 -0.4408 0 -2.0 1e-06 
0.0 -0.4407 0 -2.0 1e-06 
0.0 -0.4406 0 -2.0 1e-06 
0.0 -0.4405 0 -2.0 1e-06 
0.0 -0.4404 0 -2.0 1e-06 
0.0 -0.4403 0 -2.0 1e-06 
0.0 -0.4402 0 -2.0 1e-06 
0.0 -0.4401 0 -2.0 1e-06 
0.0 -0.44 0 -2.0 1e-06 
0.0 -0.4399 0 -2.0 1e-06 
0.0 -0.4398 0 -2.0 1e-06 
0.0 -0.4397 0 -2.0 1e-06 
0.0 -0.4396 0 -2.0 1e-06 
0.0 -0.4395 0 -2.0 1e-06 
0.0 -0.4394 0 -2.0 1e-06 
0.0 -0.4393 0 -2.0 1e-06 
0.0 -0.4392 0 -2.0 1e-06 
0.0 -0.4391 0 -2.0 1e-06 
0.0 -0.439 0 -2.0 1e-06 
0.0 -0.4389 0 -2.0 1e-06 
0.0 -0.4388 0 -2.0 1e-06 
0.0 -0.4387 0 -2.0 1e-06 
0.0 -0.4386 0 -2.0 1e-06 
0.0 -0.4385 0 -2.0 1e-06 
0.0 -0.4384 0 -2.0 1e-06 
0.0 -0.4383 0 -2.0 1e-06 
0.0 -0.4382 0 -2.0 1e-06 
0.0 -0.4381 0 -2.0 1e-06 
0.0 -0.438 0 -2.0 1e-06 
0.0 -0.4379 0 -2.0 1e-06 
0.0 -0.4378 0 -2.0 1e-06 
0.0 -0.4377 0 -2.0 1e-06 
0.0 -0.4376 0 -2.0 1e-06 
0.0 -0.4375 0 -2.0 1e-06 
0.0 -0.4374 0 -2.0 1e-06 
0.0 -0.4373 0 -2.0 1e-06 
0.0 -0.4372 0 -2.0 1e-06 
0.0 -0.4371 0 -2.0 1e-06 
0.0 -0.437 0 -2.0 1e-06 
0.0 -0.4369 0 -2.0 1e-06 
0.0 -0.4368 0 -2.0 1e-06 
0.0 -0.4367 0 -2.0 1e-06 
0.0 -0.4366 0 -2.0 1e-06 
0.0 -0.4365 0 -2.0 1e-06 
0.0 -0.4364 0 -2.0 1e-06 
0.0 -0.4363 0 -2.0 1e-06 
0.0 -0.4362 0 -2.0 1e-06 
0.0 -0.4361 0 -2.0 1e-06 
0.0 -0.436 0 -2.0 1e-06 
0.0 -0.4359 0 -2.0 1e-06 
0.0 -0.4358 0 -2.0 1e-06 
0.0 -0.4357 0 -2.0 1e-06 
0.0 -0.4356 0 -2.0 1e-06 
0.0 -0.4355 0 -2.0 1e-06 
0.0 -0.4354 0 -2.0 1e-06 
0.0 -0.4353 0 -2.0 1e-06 
0.0 -0.4352 0 -2.0 1e-06 
0.0 -0.4351 0 -2.0 1e-06 
0.0 -0.435 0 -2.0 1e-06 
0.0 -0.4349 0 -2.0 1e-06 
0.0 -0.4348 0 -2.0 1e-06 
0.0 -0.4347 0 -2.0 1e-06 
0.0 -0.4346 0 -2.0 1e-06 
0.0 -0.4345 0 -2.0 1e-06 
0.0 -0.4344 0 -2.0 1e-06 
0.0 -0.4343 0 -2.0 1e-06 
0.0 -0.4342 0 -2.0 1e-06 
0.0 -0.4341 0 -2.0 1e-06 
0.0 -0.434 0 -2.0 1e-06 
0.0 -0.4339 0 -2.0 1e-06 
0.0 -0.4338 0 -2.0 1e-06 
0.0 -0.4337 0 -2.0 1e-06 
0.0 -0.4336 0 -2.0 1e-06 
0.0 -0.4335 0 -2.0 1e-06 
0.0 -0.4334 0 -2.0 1e-06 
0.0 -0.4333 0 -2.0 1e-06 
0.0 -0.4332 0 -2.0 1e-06 
0.0 -0.4331 0 -2.0 1e-06 
0.0 -0.433 0 -2.0 1e-06 
0.0 -0.4329 0 -2.0 1e-06 
0.0 -0.4328 0 -2.0 1e-06 
0.0 -0.4327 0 -2.0 1e-06 
0.0 -0.4326 0 -2.0 1e-06 
0.0 -0.4325 0 -2.0 1e-06 
0.0 -0.4324 0 -2.0 1e-06 
0.0 -0.4323 0 -2.0 1e-06 
0.0 -0.4322 0 -2.0 1e-06 
0.0 -0.4321 0 -2.0 1e-06 
0.0 -0.432 0 -2.0 1e-06 
0.0 -0.4319 0 -2.0 1e-06 
0.0 -0.4318 0 -2.0 1e-06 
0.0 -0.4317 0 -2.0 1e-06 
0.0 -0.4316 0 -2.0 1e-06 
0.0 -0.4315 0 -2.0 1e-06 
0.0 -0.4314 0 -2.0 1e-06 
0.0 -0.4313 0 -2.0 1e-06 
0.0 -0.4312 0 -2.0 1e-06 
0.0 -0.4311 0 -2.0 1e-06 
0.0 -0.431 0 -2.0 1e-06 
0.0 -0.4309 0 -2.0 1e-06 
0.0 -0.4308 0 -2.0 1e-06 
0.0 -0.4307 0 -2.0 1e-06 
0.0 -0.4306 0 -2.0 1e-06 
0.0 -0.4305 0 -2.0 1e-06 
0.0 -0.4304 0 -2.0 1e-06 
0.0 -0.4303 0 -2.0 1e-06 
0.0 -0.4302 0 -2.0 1e-06 
0.0 -0.4301 0 -2.0 1e-06 
0.0 -0.43 0 -2.0 1e-06 
0.0 -0.4299 0 -2.0 1e-06 
0.0 -0.4298 0 -2.0 1e-06 
0.0 -0.4297 0 -2.0 1e-06 
0.0 -0.4296 0 -2.0 1e-06 
0.0 -0.4295 0 -2.0 1e-06 
0.0 -0.4294 0 -2.0 1e-06 
0.0 -0.4293 0 -2.0 1e-06 
0.0 -0.4292 0 -2.0 1e-06 
0.0 -0.4291 0 -2.0 1e-06 
0.0 -0.429 0 -2.0 1e-06 
0.0 -0.4289 0 -2.0 1e-06 
0.0 -0.4288 0 -2.0 1e-06 
0.0 -0.4287 0 -2.0 1e-06 
0.0 -0.4286 0 -2.0 1e-06 
0.0 -0.4285 0 -2.0 1e-06 
0.0 -0.4284 0 -2.0 1e-06 
0.0 -0.4283 0 -2.0 1e-06 
0.0 -0.4282 0 -2.0 1e-06 
0.0 -0.4281 0 -2.0 1e-06 
0.0 -0.428 0 -2.0 1e-06 
0.0 -0.4279 0 -2.0 1e-06 
0.0 -0.4278 0 -2.0 1e-06 
0.0 -0.4277 0 -2.0 1e-06 
0.0 -0.4276 0 -2.0 1e-06 
0.0 -0.4275 0 -2.0 1e-06 
0.0 -0.4274 0 -2.0 1e-06 
0.0 -0.4273 0 -2.0 1e-06 
0.0 -0.4272 0 -2.0 1e-06 
0.0 -0.4271 0 -2.0 1e-06 
0.0 -0.427 0 -2.0 1e-06 
0.0 -0.4269 0 -2.0 1e-06 
0.0 -0.4268 0 -2.0 1e-06 
0.0 -0.4267 0 -2.0 1e-06 
0.0 -0.4266 0 -2.0 1e-06 
0.0 -0.4265 0 -2.0 1e-06 
0.0 -0.4264 0 -2.0 1e-06 
0.0 -0.4263 0 -2.0 1e-06 
0.0 -0.4262 0 -2.0 1e-06 
0.0 -0.4261 0 -2.0 1e-06 
0.0 -0.426 0 -2.0 1e-06 
0.0 -0.4259 0 -2.0 1e-06 
0.0 -0.4258 0 -2.0 1e-06 
0.0 -0.4257 0 -2.0 1e-06 
0.0 -0.4256 0 -2.0 1e-06 
0.0 -0.4255 0 -2.0 1e-06 
0.0 -0.4254 0 -2.0 1e-06 
0.0 -0.4253 0 -2.0 1e-06 
0.0 -0.4252 0 -2.0 1e-06 
0.0 -0.4251 0 -2.0 1e-06 
0.0 -0.425 0 -2.0 1e-06 
0.0 -0.4249 0 -2.0 1e-06 
0.0 -0.4248 0 -2.0 1e-06 
0.0 -0.4247 0 -2.0 1e-06 
0.0 -0.4246 0 -2.0 1e-06 
0.0 -0.4245 0 -2.0 1e-06 
0.0 -0.4244 0 -2.0 1e-06 
0.0 -0.4243 0 -2.0 1e-06 
0.0 -0.4242 0 -2.0 1e-06 
0.0 -0.4241 0 -2.0 1e-06 
0.0 -0.424 0 -2.0 1e-06 
0.0 -0.4239 0 -2.0 1e-06 
0.0 -0.4238 0 -2.0 1e-06 
0.0 -0.4237 0 -2.0 1e-06 
0.0 -0.4236 0 -2.0 1e-06 
0.0 -0.4235 0 -2.0 1e-06 
0.0 -0.4234 0 -2.0 1e-06 
0.0 -0.4233 0 -2.0 1e-06 
0.0 -0.4232 0 -2.0 1e-06 
0.0 -0.4231 0 -2.0 1e-06 
0.0 -0.423 0 -2.0 1e-06 
0.0 -0.4229 0 -2.0 1e-06 
0.0 -0.4228 0 -2.0 1e-06 
0.0 -0.4227 0 -2.0 1e-06 
0.0 -0.4226 0 -2.0 1e-06 
0.0 -0.4225 0 -2.0 1e-06 
0.0 -0.4224 0 -2.0 1e-06 
0.0 -0.4223 0 -2.0 1e-06 
0.0 -0.4222 0 -2.0 1e-06 
0.0 -0.4221 0 -2.0 1e-06 
0.0 -0.422 0 -2.0 1e-06 
0.0 -0.4219 0 -2.0 1e-06 
0.0 -0.4218 0 -2.0 1e-06 
0.0 -0.4217 0 -2.0 1e-06 
0.0 -0.4216 0 -2.0 1e-06 
0.0 -0.4215 0 -2.0 1e-06 
0.0 -0.4214 0 -2.0 1e-06 
0.0 -0.4213 0 -2.0 1e-06 
0.0 -0.4212 0 -2.0 1e-06 
0.0 -0.4211 0 -2.0 1e-06 
0.0 -0.421 0 -2.0 1e-06 
0.0 -0.4209 0 -2.0 1e-06 
0.0 -0.4208 0 -2.0 1e-06 
0.0 -0.4207 0 -2.0 1e-06 
0.0 -0.4206 0 -2.0 1e-06 
0.0 -0.4205 0 -2.0 1e-06 
0.0 -0.4204 0 -2.0 1e-06 
0.0 -0.4203 0 -2.0 1e-06 
0.0 -0.4202 0 -2.0 1e-06 
0.0 -0.4201 0 -2.0 1e-06 
0.0 -0.42 0 -2.0 1e-06 
0.0 -0.4199 0 -2.0 1e-06 
0.0 -0.4198 0 -2.0 1e-06 
0.0 -0.4197 0 -2.0 1e-06 
0.0 -0.4196 0 -2.0 1e-06 
0.0 -0.4195 0 -2.0 1e-06 
0.0 -0.4194 0 -2.0 1e-06 
0.0 -0.4193 0 -2.0 1e-06 
0.0 -0.4192 0 -2.0 1e-06 
0.0 -0.4191 0 -2.0 1e-06 
0.0 -0.419 0 -2.0 1e-06 
0.0 -0.4189 0 -2.0 1e-06 
0.0 -0.4188 0 -2.0 1e-06 
0.0 -0.4187 0 -2.0 1e-06 
0.0 -0.4186 0 -2.0 1e-06 
0.0 -0.4185 0 -2.0 1e-06 
0.0 -0.4184 0 -2.0 1e-06 
0.0 -0.4183 0 -2.0 1e-06 
0.0 -0.4182 0 -2.0 1e-06 
0.0 -0.4181 0 -2.0 1e-06 
0.0 -0.418 0 -2.0 1e-06 
0.0 -0.4179 0 -2.0 1e-06 
0.0 -0.4178 0 -2.0 1e-06 
0.0 -0.4177 0 -2.0 1e-06 
0.0 -0.4176 0 -2.0 1e-06 
0.0 -0.4175 0 -2.0 1e-06 
0.0 -0.4174 0 -2.0 1e-06 
0.0 -0.4173 0 -2.0 1e-06 
0.0 -0.4172 0 -2.0 1e-06 
0.0 -0.4171 0 -2.0 1e-06 
0.0 -0.417 0 -2.0 1e-06 
0.0 -0.4169 0 -2.0 1e-06 
0.0 -0.4168 0 -2.0 1e-06 
0.0 -0.4167 0 -2.0 1e-06 
0.0 -0.4166 0 -2.0 1e-06 
0.0 -0.4165 0 -2.0 1e-06 
0.0 -0.4164 0 -2.0 1e-06 
0.0 -0.4163 0 -2.0 1e-06 
0.0 -0.4162 0 -2.0 1e-06 
0.0 -0.4161 0 -2.0 1e-06 
0.0 -0.416 0 -2.0 1e-06 
0.0 -0.4159 0 -2.0 1e-06 
0.0 -0.4158 0 -2.0 1e-06 
0.0 -0.4157 0 -2.0 1e-06 
0.0 -0.4156 0 -2.0 1e-06 
0.0 -0.4155 0 -2.0 1e-06 
0.0 -0.4154 0 -2.0 1e-06 
0.0 -0.4153 0 -2.0 1e-06 
0.0 -0.4152 0 -2.0 1e-06 
0.0 -0.4151 0 -2.0 1e-06 
0.0 -0.415 0 -2.0 1e-06 
0.0 -0.4149 0 -2.0 1e-06 
0.0 -0.4148 0 -2.0 1e-06 
0.0 -0.4147 0 -2.0 1e-06 
0.0 -0.4146 0 -2.0 1e-06 
0.0 -0.4145 0 -2.0 1e-06 
0.0 -0.4144 0 -2.0 1e-06 
0.0 -0.4143 0 -2.0 1e-06 
0.0 -0.4142 0 -2.0 1e-06 
0.0 -0.4141 0 -2.0 1e-06 
0.0 -0.414 0 -2.0 1e-06 
0.0 -0.4139 0 -2.0 1e-06 
0.0 -0.4138 0 -2.0 1e-06 
0.0 -0.4137 0 -2.0 1e-06 
0.0 -0.4136 0 -2.0 1e-06 
0.0 -0.4135 0 -2.0 1e-06 
0.0 -0.4134 0 -2.0 1e-06 
0.0 -0.4133 0 -2.0 1e-06 
0.0 -0.4132 0 -2.0 1e-06 
0.0 -0.4131 0 -2.0 1e-06 
0.0 -0.413 0 -2.0 1e-06 
0.0 -0.4129 0 -2.0 1e-06 
0.0 -0.4128 0 -2.0 1e-06 
0.0 -0.4127 0 -2.0 1e-06 
0.0 -0.4126 0 -2.0 1e-06 
0.0 -0.4125 0 -2.0 1e-06 
0.0 -0.4124 0 -2.0 1e-06 
0.0 -0.4123 0 -2.0 1e-06 
0.0 -0.4122 0 -2.0 1e-06 
0.0 -0.4121 0 -2.0 1e-06 
0.0 -0.412 0 -2.0 1e-06 
0.0 -0.4119 0 -2.0 1e-06 
0.0 -0.4118 0 -2.0 1e-06 
0.0 -0.4117 0 -2.0 1e-06 
0.0 -0.4116 0 -2.0 1e-06 
0.0 -0.4115 0 -2.0 1e-06 
0.0 -0.4114 0 -2.0 1e-06 
0.0 -0.4113 0 -2.0 1e-06 
0.0 -0.4112 0 -2.0 1e-06 
0.0 -0.4111 0 -2.0 1e-06 
0.0 -0.411 0 -2.0 1e-06 
0.0 -0.4109 0 -2.0 1e-06 
0.0 -0.4108 0 -2.0 1e-06 
0.0 -0.4107 0 -2.0 1e-06 
0.0 -0.4106 0 -2.0 1e-06 
0.0 -0.4105 0 -2.0 1e-06 
0.0 -0.4104 0 -2.0 1e-06 
0.0 -0.4103 0 -2.0 1e-06 
0.0 -0.4102 0 -2.0 1e-06 
0.0 -0.4101 0 -2.0 1e-06 
0.0 -0.41 0 -2.0 1e-06 
0.0 -0.4099 0 -2.0 1e-06 
0.0 -0.4098 0 -2.0 1e-06 
0.0 -0.4097 0 -2.0 1e-06 
0.0 -0.4096 0 -2.0 1e-06 
0.0 -0.4095 0 -2.0 1e-06 
0.0 -0.4094 0 -2.0 1e-06 
0.0 -0.4093 0 -2.0 1e-06 
0.0 -0.4092 0 -2.0 1e-06 
0.0 -0.4091 0 -2.0 1e-06 
0.0 -0.409 0 -2.0 1e-06 
0.0 -0.4089 0 -2.0 1e-06 
0.0 -0.4088 0 -2.0 1e-06 
0.0 -0.4087 0 -2.0 1e-06 
0.0 -0.4086 0 -2.0 1e-06 
0.0 -0.4085 0 -2.0 1e-06 
0.0 -0.4084 0 -2.0 1e-06 
0.0 -0.4083 0 -2.0 1e-06 
0.0 -0.4082 0 -2.0 1e-06 
0.0 -0.4081 0 -2.0 1e-06 
0.0 -0.408 0 -2.0 1e-06 
0.0 -0.4079 0 -2.0 1e-06 
0.0 -0.4078 0 -2.0 1e-06 
0.0 -0.4077 0 -2.0 1e-06 
0.0 -0.4076 0 -2.0 1e-06 
0.0 -0.4075 0 -2.0 1e-06 
0.0 -0.4074 0 -2.0 1e-06 
0.0 -0.4073 0 -2.0 1e-06 
0.0 -0.4072 0 -2.0 1e-06 
0.0 -0.4071 0 -2.0 1e-06 
0.0 -0.407 0 -2.0 1e-06 
0.0 -0.4069 0 -2.0 1e-06 
0.0 -0.4068 0 -2.0 1e-06 
0.0 -0.4067 0 -2.0 1e-06 
0.0 -0.4066 0 -2.0 1e-06 
0.0 -0.4065 0 -2.0 1e-06 
0.0 -0.4064 0 -2.0 1e-06 
0.0 -0.4063 0 -2.0 1e-06 
0.0 -0.4062 0 -2.0 1e-06 
0.0 -0.4061 0 -2.0 1e-06 
0.0 -0.406 0 -2.0 1e-06 
0.0 -0.4059 0 -2.0 1e-06 
0.0 -0.4058 0 -2.0 1e-06 
0.0 -0.4057 0 -2.0 1e-06 
0.0 -0.4056 0 -2.0 1e-06 
0.0 -0.4055 0 -2.0 1e-06 
0.0 -0.4054 0 -2.0 1e-06 
0.0 -0.4053 0 -2.0 1e-06 
0.0 -0.4052 0 -2.0 1e-06 
0.0 -0.4051 0 -2.0 1e-06 
0.0 -0.405 0 -2.0 1e-06 
0.0 -0.4049 0 -2.0 1e-06 
0.0 -0.4048 0 -2.0 1e-06 
0.0 -0.4047 0 -2.0 1e-06 
0.0 -0.4046 0 -2.0 1e-06 
0.0 -0.4045 0 -2.0 1e-06 
0.0 -0.4044 0 -2.0 1e-06 
0.0 -0.4043 0 -2.0 1e-06 
0.0 -0.4042 0 -2.0 1e-06 
0.0 -0.4041 0 -2.0 1e-06 
0.0 -0.404 0 -2.0 1e-06 
0.0 -0.4039 0 -2.0 1e-06 
0.0 -0.4038 0 -2.0 1e-06 
0.0 -0.4037 0 -2.0 1e-06 
0.0 -0.4036 0 -2.0 1e-06 
0.0 -0.4035 0 -2.0 1e-06 
0.0 -0.4034 0 -2.0 1e-06 
0.0 -0.4033 0 -2.0 1e-06 
0.0 -0.4032 0 -2.0 1e-06 
0.0 -0.4031 0 -2.0 1e-06 
0.0 -0.403 0 -2.0 1e-06 
0.0 -0.4029 0 -2.0 1e-06 
0.0 -0.4028 0 -2.0 1e-06 
0.0 -0.4027 0 -2.0 1e-06 
0.0 -0.4026 0 -2.0 1e-06 
0.0 -0.4025 0 -2.0 1e-06 
0.0 -0.4024 0 -2.0 1e-06 
0.0 -0.4023 0 -2.0 1e-06 
0.0 -0.4022 0 -2.0 1e-06 
0.0 -0.4021 0 -2.0 1e-06 
0.0 -0.402 0 -2.0 1e-06 
0.0 -0.4019 0 -2.0 1e-06 
0.0 -0.4018 0 -2.0 1e-06 
0.0 -0.4017 0 -2.0 1e-06 
0.0 -0.4016 0 -2.0 1e-06 
0.0 -0.4015 0 -2.0 1e-06 
0.0 -0.4014 0 -2.0 1e-06 
0.0 -0.4013 0 -2.0 1e-06 
0.0 -0.4012 0 -2.0 1e-06 
0.0 -0.4011 0 -2.0 1e-06 
0.0 -0.401 0 -2.0 1e-06 
0.0 -0.4009 0 -2.0 1e-06 
0.0 -0.4008 0 -2.0 1e-06 
0.0 -0.4007 0 -2.0 1e-06 
0.0 -0.4006 0 -2.0 1e-06 
0.0 -0.4005 0 -2.0 1e-06 
0.0 -0.4004 0 -2.0 1e-06 
0.0 -0.4003 0 -2.0 1e-06 
0.0 -0.4002 0 -2.0 1e-06 
0.0 -0.4001 0 -2.0 1e-06 
0.0 -0.4 0 -2.0 1e-06 
0.0 -0.3999 0 -2.0 1e-06 
0.0 -0.3998 0 -2.0 1e-06 
0.0 -0.3997 0 -2.0 1e-06 
0.0 -0.3996 0 -2.0 1e-06 
0.0 -0.3995 0 -2.0 1e-06 
0.0 -0.3994 0 -2.0 1e-06 
0.0 -0.3993 0 -2.0 1e-06 
0.0 -0.3992 0 -2.0 1e-06 
0.0 -0.3991 0 -2.0 1e-06 
0.0 -0.399 0 -2.0 1e-06 
0.0 -0.3989 0 -2.0 1e-06 
0.0 -0.3988 0 -2.0 1e-06 
0.0 -0.3987 0 -2.0 1e-06 
0.0 -0.3986 0 -2.0 1e-06 
0.0 -0.3985 0 -2.0 1e-06 
0.0 -0.3984 0 -2.0 1e-06 
0.0 -0.3983 0 -2.0 1e-06 
0.0 -0.3982 0 -2.0 1e-06 
0.0 -0.3981 0 -2.0 1e-06 
0.0 -0.398 0 -2.0 1e-06 
0.0 -0.3979 0 -2.0 1e-06 
0.0 -0.3978 0 -2.0 1e-06 
0.0 -0.3977 0 -2.0 1e-06 
0.0 -0.3976 0 -2.0 1e-06 
0.0 -0.3975 0 -2.0 1e-06 
0.0 -0.3974 0 -2.0 1e-06 
0.0 -0.3973 0 -2.0 1e-06 
0.0 -0.3972 0 -2.0 1e-06 
0.0 -0.3971 0 -2.0 1e-06 
0.0 -0.397 0 -2.0 1e-06 
0.0 -0.3969 0 -2.0 1e-06 
0.0 -0.3968 0 -2.0 1e-06 
0.0 -0.3967 0 -2.0 1e-06 
0.0 -0.3966 0 -2.0 1e-06 
0.0 -0.3965 0 -2.0 1e-06 
0.0 -0.3964 0 -2.0 1e-06 
0.0 -0.3963 0 -2.0 1e-06 
0.0 -0.3962 0 -2.0 1e-06 
0.0 -0.3961 0 -2.0 1e-06 
0.0 -0.396 0 -2.0 1e-06 
0.0 -0.3959 0 -2.0 1e-06 
0.0 -0.3958 0 -2.0 1e-06 
0.0 -0.3957 0 -2.0 1e-06 
0.0 -0.3956 0 -2.0 1e-06 
0.0 -0.3955 0 -2.0 1e-06 
0.0 -0.3954 0 -2.0 1e-06 
0.0 -0.3953 0 -2.0 1e-06 
0.0 -0.3952 0 -2.0 1e-06 
0.0 -0.3951 0 -2.0 1e-06 
0.0 -0.395 0 -2.0 1e-06 
0.0 -0.3949 0 -2.0 1e-06 
0.0 -0.3948 0 -2.0 1e-06 
0.0 -0.3947 0 -2.0 1e-06 
0.0 -0.3946 0 -2.0 1e-06 
0.0 -0.3945 0 -2.0 1e-06 
0.0 -0.3944 0 -2.0 1e-06 
0.0 -0.3943 0 -2.0 1e-06 
0.0 -0.3942 0 -2.0 1e-06 
0.0 -0.3941 0 -2.0 1e-06 
0.0 -0.394 0 -2.0 1e-06 
0.0 -0.3939 0 -2.0 1e-06 
0.0 -0.3938 0 -2.0 1e-06 
0.0 -0.3937 0 -2.0 1e-06 
0.0 -0.3936 0 -2.0 1e-06 
0.0 -0.3935 0 -2.0 1e-06 
0.0 -0.3934 0 -2.0 1e-06 
0.0 -0.3933 0 -2.0 1e-06 
0.0 -0.3932 0 -2.0 1e-06 
0.0 -0.3931 0 -2.0 1e-06 
0.0 -0.393 0 -2.0 1e-06 
0.0 -0.3929 0 -2.0 1e-06 
0.0 -0.3928 0 -2.0 1e-06 
0.0 -0.3927 0 -2.0 1e-06 
0.0 -0.3926 0 -2.0 1e-06 
0.0 -0.3925 0 -2.0 1e-06 
0.0 -0.3924 0 -2.0 1e-06 
0.0 -0.3923 0 -2.0 1e-06 
0.0 -0.3922 0 -2.0 1e-06 
0.0 -0.3921 0 -2.0 1e-06 
0.0 -0.392 0 -2.0 1e-06 
0.0 -0.3919 0 -2.0 1e-06 
0.0 -0.3918 0 -2.0 1e-06 
0.0 -0.3917 0 -2.0 1e-06 
0.0 -0.3916 0 -2.0 1e-06 
0.0 -0.3915 0 -2.0 1e-06 
0.0 -0.3914 0 -2.0 1e-06 
0.0 -0.3913 0 -2.0 1e-06 
0.0 -0.3912 0 -2.0 1e-06 
0.0 -0.3911 0 -2.0 1e-06 
0.0 -0.391 0 -2.0 1e-06 
0.0 -0.3909 0 -2.0 1e-06 
0.0 -0.3908 0 -2.0 1e-06 
0.0 -0.3907 0 -2.0 1e-06 
0.0 -0.3906 0 -2.0 1e-06 
0.0 -0.3905 0 -2.0 1e-06 
0.0 -0.3904 0 -2.0 1e-06 
0.0 -0.3903 0 -2.0 1e-06 
0.0 -0.3902 0 -2.0 1e-06 
0.0 -0.3901 0 -2.0 1e-06 
0.0 -0.39 0 -2.0 1e-06 
0.0 -0.3899 0 -2.0 1e-06 
0.0 -0.3898 0 -2.0 1e-06 
0.0 -0.3897 0 -2.0 1e-06 
0.0 -0.3896 0 -2.0 1e-06 
0.0 -0.3895 0 -2.0 1e-06 
0.0 -0.3894 0 -2.0 1e-06 
0.0 -0.3893 0 -2.0 1e-06 
0.0 -0.3892 0 -2.0 1e-06 
0.0 -0.3891 0 -2.0 1e-06 
0.0 -0.389 0 -2.0 1e-06 
0.0 -0.3889 0 -2.0 1e-06 
0.0 -0.3888 0 -2.0 1e-06 
0.0 -0.3887 0 -2.0 1e-06 
0.0 -0.3886 0 -2.0 1e-06 
0.0 -0.3885 0 -2.0 1e-06 
0.0 -0.3884 0 -2.0 1e-06 
0.0 -0.3883 0 -2.0 1e-06 
0.0 -0.3882 0 -2.0 1e-06 
0.0 -0.3881 0 -2.0 1e-06 
0.0 -0.388 0 -2.0 1e-06 
0.0 -0.3879 0 -2.0 1e-06 
0.0 -0.3878 0 -2.0 1e-06 
0.0 -0.3877 0 -2.0 1e-06 
0.0 -0.3876 0 -2.0 1e-06 
0.0 -0.3875 0 -2.0 1e-06 
0.0 -0.3874 0 -2.0 1e-06 
0.0 -0.3873 0 -2.0 1e-06 
0.0 -0.3872 0 -2.0 1e-06 
0.0 -0.3871 0 -2.0 1e-06 
0.0 -0.387 0 -2.0 1e-06 
0.0 -0.3869 0 -2.0 1e-06 
0.0 -0.3868 0 -2.0 1e-06 
0.0 -0.3867 0 -2.0 1e-06 
0.0 -0.3866 0 -2.0 1e-06 
0.0 -0.3865 0 -2.0 1e-06 
0.0 -0.3864 0 -2.0 1e-06 
0.0 -0.3863 0 -2.0 1e-06 
0.0 -0.3862 0 -2.0 1e-06 
0.0 -0.3861 0 -2.0 1e-06 
0.0 -0.386 0 -2.0 1e-06 
0.0 -0.3859 0 -2.0 1e-06 
0.0 -0.3858 0 -2.0 1e-06 
0.0 -0.3857 0 -2.0 1e-06 
0.0 -0.3856 0 -2.0 1e-06 
0.0 -0.3855 0 -2.0 1e-06 
0.0 -0.3854 0 -2.0 1e-06 
0.0 -0.3853 0 -2.0 1e-06 
0.0 -0.3852 0 -2.0 1e-06 
0.0 -0.3851 0 -2.0 1e-06 
0.0 -0.385 0 -2.0 1e-06 
0.0 -0.3849 0 -2.0 1e-06 
0.0 -0.3848 0 -2.0 1e-06 
0.0 -0.3847 0 -2.0 1e-06 
0.0 -0.3846 0 -2.0 1e-06 
0.0 -0.3845 0 -2.0 1e-06 
0.0 -0.3844 0 -2.0 1e-06 
0.0 -0.3843 0 -2.0 1e-06 
0.0 -0.3842 0 -2.0 1e-06 
0.0 -0.3841 0 -2.0 1e-06 
0.0 -0.384 0 -2.0 1e-06 
0.0 -0.3839 0 -2.0 1e-06 
0.0 -0.3838 0 -2.0 1e-06 
0.0 -0.3837 0 -2.0 1e-06 
0.0 -0.3836 0 -2.0 1e-06 
0.0 -0.3835 0 -2.0 1e-06 
0.0 -0.3834 0 -2.0 1e-06 
0.0 -0.3833 0 -2.0 1e-06 
0.0 -0.3832 0 -2.0 1e-06 
0.0 -0.3831 0 -2.0 1e-06 
0.0 -0.383 0 -2.0 1e-06 
0.0 -0.3829 0 -2.0 1e-06 
0.0 -0.3828 0 -2.0 1e-06 
0.0 -0.3827 0 -2.0 1e-06 
0.0 -0.3826 0 -2.0 1e-06 
0.0 -0.3825 0 -2.0 1e-06 
0.0 -0.3824 0 -2.0 1e-06 
0.0 -0.3823 0 -2.0 1e-06 
0.0 -0.3822 0 -2.0 1e-06 
0.0 -0.3821 0 -2.0 1e-06 
0.0 -0.382 0 -2.0 1e-06 
0.0 -0.3819 0 -2.0 1e-06 
0.0 -0.3818 0 -2.0 1e-06 
0.0 -0.3817 0 -2.0 1e-06 
0.0 -0.3816 0 -2.0 1e-06 
0.0 -0.3815 0 -2.0 1e-06 
0.0 -0.3814 0 -2.0 1e-06 
0.0 -0.3813 0 -2.0 1e-06 
0.0 -0.3812 0 -2.0 1e-06 
0.0 -0.3811 0 -2.0 1e-06 
0.0 -0.381 0 -2.0 1e-06 
0.0 -0.3809 0 -2.0 1e-06 
0.0 -0.3808 0 -2.0 1e-06 
0.0 -0.3807 0 -2.0 1e-06 
0.0 -0.3806 0 -2.0 1e-06 
0.0 -0.3805 0 -2.0 1e-06 
0.0 -0.3804 0 -2.0 1e-06 
0.0 -0.3803 0 -2.0 1e-06 
0.0 -0.3802 0 -2.0 1e-06 
0.0 -0.3801 0 -2.0 1e-06 
0.0 -0.38 0 -2.0 1e-06 
0.0 -0.3799 0 -2.0 1e-06 
0.0 -0.3798 0 -2.0 1e-06 
0.0 -0.3797 0 -2.0 1e-06 
0.0 -0.3796 0 -2.0 1e-06 
0.0 -0.3795 0 -2.0 1e-06 
0.0 -0.3794 0 -2.0 1e-06 
0.0 -0.3793 0 -2.0 1e-06 
0.0 -0.3792 0 -2.0 1e-06 
0.0 -0.3791 0 -2.0 1e-06 
0.0 -0.379 0 -2.0 1e-06 
0.0 -0.3789 0 -2.0 1e-06 
0.0 -0.3788 0 -2.0 1e-06 
0.0 -0.3787 0 -2.0 1e-06 
0.0 -0.3786 0 -2.0 1e-06 
0.0 -0.3785 0 -2.0 1e-06 
0.0 -0.3784 0 -2.0 1e-06 
0.0 -0.3783 0 -2.0 1e-06 
0.0 -0.3782 0 -2.0 1e-06 
0.0 -0.3781 0 -2.0 1e-06 
0.0 -0.378 0 -2.0 1e-06 
0.0 -0.3779 0 -2.0 1e-06 
0.0 -0.3778 0 -2.0 1e-06 
0.0 -0.3777 0 -2.0 1e-06 
0.0 -0.3776 0 -2.0 1e-06 
0.0 -0.3775 0 -2.0 1e-06 
0.0 -0.3774 0 -2.0 1e-06 
0.0 -0.3773 0 -2.0 1e-06 
0.0 -0.3772 0 -2.0 1e-06 
0.0 -0.3771 0 -2.0 1e-06 
0.0 -0.377 0 -2.0 1e-06 
0.0 -0.3769 0 -2.0 1e-06 
0.0 -0.3768 0 -2.0 1e-06 
0.0 -0.3767 0 -2.0 1e-06 
0.0 -0.3766 0 -2.0 1e-06 
0.0 -0.3765 0 -2.0 1e-06 
0.0 -0.3764 0 -2.0 1e-06 
0.0 -0.3763 0 -2.0 1e-06 
0.0 -0.3762 0 -2.0 1e-06 
0.0 -0.3761 0 -2.0 1e-06 
0.0 -0.376 0 -2.0 1e-06 
0.0 -0.3759 0 -2.0 1e-06 
0.0 -0.3758 0 -2.0 1e-06 
0.0 -0.3757 0 -2.0 1e-06 
0.0 -0.3756 0 -2.0 1e-06 
0.0 -0.3755 0 -2.0 1e-06 
0.0 -0.3754 0 -2.0 1e-06 
0.0 -0.3753 0 -2.0 1e-06 
0.0 -0.3752 0 -2.0 1e-06 
0.0 -0.3751 0 -2.0 1e-06 
0.0 -0.375 0 -2.0 1e-06 
0.0 -0.3749 0 -2.0 1e-06 
0.0 -0.3748 0 -2.0 1e-06 
0.0 -0.3747 0 -2.0 1e-06 
0.0 -0.3746 0 -2.0 1e-06 
0.0 -0.3745 0 -2.0 1e-06 
0.0 -0.3744 0 -2.0 1e-06 
0.0 -0.3743 0 -2.0 1e-06 
0.0 -0.3742 0 -2.0 1e-06 
0.0 -0.3741 0 -2.0 1e-06 
0.0 -0.374 0 -2.0 1e-06 
0.0 -0.3739 0 -2.0 1e-06 
0.0 -0.3738 0 -2.0 1e-06 
0.0 -0.3737 0 -2.0 1e-06 
0.0 -0.3736 0 -2.0 1e-06 
0.0 -0.3735 0 -2.0 1e-06 
0.0 -0.3734 0 -2.0 1e-06 
0.0 -0.3733 0 -2.0 1e-06 
0.0 -0.3732 0 -2.0 1e-06 
0.0 -0.3731 0 -2.0 1e-06 
0.0 -0.373 0 -2.0 1e-06 
0.0 -0.3729 0 -2.0 1e-06 
0.0 -0.3728 0 -2.0 1e-06 
0.0 -0.3727 0 -2.0 1e-06 
0.0 -0.3726 0 -2.0 1e-06 
0.0 -0.3725 0 -2.0 1e-06 
0.0 -0.3724 0 -2.0 1e-06 
0.0 -0.3723 0 -2.0 1e-06 
0.0 -0.3722 0 -2.0 1e-06 
0.0 -0.3721 0 -2.0 1e-06 
0.0 -0.372 0 -2.0 1e-06 
0.0 -0.3719 0 -2.0 1e-06 
0.0 -0.3718 0 -2.0 1e-06 
0.0 -0.3717 0 -2.0 1e-06 
0.0 -0.3716 0 -2.0 1e-06 
0.0 -0.3715 0 -2.0 1e-06 
0.0 -0.3714 0 -2.0 1e-06 
0.0 -0.3713 0 -2.0 1e-06 
0.0 -0.3712 0 -2.0 1e-06 
0.0 -0.3711 0 -2.0 1e-06 
0.0 -0.371 0 -2.0 1e-06 
0.0 -0.3709 0 -2.0 1e-06 
0.0 -0.3708 0 -2.0 1e-06 
0.0 -0.3707 0 -2.0 1e-06 
0.0 -0.3706 0 -2.0 1e-06 
0.0 -0.3705 0 -2.0 1e-06 
0.0 -0.3704 0 -2.0 1e-06 
0.0 -0.3703 0 -2.0 1e-06 
0.0 -0.3702 0 -2.0 1e-06 
0.0 -0.3701 0 -2.0 1e-06 
0.0 -0.37 0 -2.0 1e-06 
0.0 -0.3699 0 -2.0 1e-06 
0.0 -0.3698 0 -2.0 1e-06 
0.0 -0.3697 0 -2.0 1e-06 
0.0 -0.3696 0 -2.0 1e-06 
0.0 -0.3695 0 -2.0 1e-06 
0.0 -0.3694 0 -2.0 1e-06 
0.0 -0.3693 0 -2.0 1e-06 
0.0 -0.3692 0 -2.0 1e-06 
0.0 -0.3691 0 -2.0 1e-06 
0.0 -0.369 0 -2.0 1e-06 
0.0 -0.3689 0 -2.0 1e-06 
0.0 -0.3688 0 -2.0 1e-06 
0.0 -0.3687 0 -2.0 1e-06 
0.0 -0.3686 0 -2.0 1e-06 
0.0 -0.3685 0 -2.0 1e-06 
0.0 -0.3684 0 -2.0 1e-06 
0.0 -0.3683 0 -2.0 1e-06 
0.0 -0.3682 0 -2.0 1e-06 
0.0 -0.3681 0 -2.0 1e-06 
0.0 -0.368 0 -2.0 1e-06 
0.0 -0.3679 0 -2.0 1e-06 
0.0 -0.3678 0 -2.0 1e-06 
0.0 -0.3677 0 -2.0 1e-06 
0.0 -0.3676 0 -2.0 1e-06 
0.0 -0.3675 0 -2.0 1e-06 
0.0 -0.3674 0 -2.0 1e-06 
0.0 -0.3673 0 -2.0 1e-06 
0.0 -0.3672 0 -2.0 1e-06 
0.0 -0.3671 0 -2.0 1e-06 
0.0 -0.367 0 -2.0 1e-06 
0.0 -0.3669 0 -2.0 1e-06 
0.0 -0.3668 0 -2.0 1e-06 
0.0 -0.3667 0 -2.0 1e-06 
0.0 -0.3666 0 -2.0 1e-06 
0.0 -0.3665 0 -2.0 1e-06 
0.0 -0.3664 0 -2.0 1e-06 
0.0 -0.3663 0 -2.0 1e-06 
0.0 -0.3662 0 -2.0 1e-06 
0.0 -0.3661 0 -2.0 1e-06 
0.0 -0.366 0 -2.0 1e-06 
0.0 -0.3659 0 -2.0 1e-06 
0.0 -0.3658 0 -2.0 1e-06 
0.0 -0.3657 0 -2.0 1e-06 
0.0 -0.3656 0 -2.0 1e-06 
0.0 -0.3655 0 -2.0 1e-06 
0.0 -0.3654 0 -2.0 1e-06 
0.0 -0.3653 0 -2.0 1e-06 
0.0 -0.3652 0 -2.0 1e-06 
0.0 -0.3651 0 -2.0 1e-06 
0.0 -0.365 0 -2.0 1e-06 
0.0 -0.3649 0 -2.0 1e-06 
0.0 -0.3648 0 -2.0 1e-06 
0.0 -0.3647 0 -2.0 1e-06 
0.0 -0.3646 0 -2.0 1e-06 
0.0 -0.3645 0 -2.0 1e-06 
0.0 -0.3644 0 -2.0 1e-06 
0.0 -0.3643 0 -2.0 1e-06 
0.0 -0.3642 0 -2.0 1e-06 
0.0 -0.3641 0 -2.0 1e-06 
0.0 -0.364 0 -2.0 1e-06 
0.0 -0.3639 0 -2.0 1e-06 
0.0 -0.3638 0 -2.0 1e-06 
0.0 -0.3637 0 -2.0 1e-06 
0.0 -0.3636 0 -2.0 1e-06 
0.0 -0.3635 0 -2.0 1e-06 
0.0 -0.3634 0 -2.0 1e-06 
0.0 -0.3633 0 -2.0 1e-06 
0.0 -0.3632 0 -2.0 1e-06 
0.0 -0.3631 0 -2.0 1e-06 
0.0 -0.363 0 -2.0 1e-06 
0.0 -0.3629 0 -2.0 1e-06 
0.0 -0.3628 0 -2.0 1e-06 
0.0 -0.3627 0 -2.0 1e-06 
0.0 -0.3626 0 -2.0 1e-06 
0.0 -0.3625 0 -2.0 1e-06 
0.0 -0.3624 0 -2.0 1e-06 
0.0 -0.3623 0 -2.0 1e-06 
0.0 -0.3622 0 -2.0 1e-06 
0.0 -0.3621 0 -2.0 1e-06 
0.0 -0.362 0 -2.0 1e-06 
0.0 -0.3619 0 -2.0 1e-06 
0.0 -0.3618 0 -2.0 1e-06 
0.0 -0.3617 0 -2.0 1e-06 
0.0 -0.3616 0 -2.0 1e-06 
0.0 -0.3615 0 -2.0 1e-06 
0.0 -0.3614 0 -2.0 1e-06 
0.0 -0.3613 0 -2.0 1e-06 
0.0 -0.3612 0 -2.0 1e-06 
0.0 -0.3611 0 -2.0 1e-06 
0.0 -0.361 0 -2.0 1e-06 
0.0 -0.3609 0 -2.0 1e-06 
0.0 -0.3608 0 -2.0 1e-06 
0.0 -0.3607 0 -2.0 1e-06 
0.0 -0.3606 0 -2.0 1e-06 
0.0 -0.3605 0 -2.0 1e-06 
0.0 -0.3604 0 -2.0 1e-06 
0.0 -0.3603 0 -2.0 1e-06 
0.0 -0.3602 0 -2.0 1e-06 
0.0 -0.3601 0 -2.0 1e-06 
0.0 -0.36 0 -2.0 1e-06 
0.0 -0.3599 0 -2.0 1e-06 
0.0 -0.3598 0 -2.0 1e-06 
0.0 -0.3597 0 -2.0 1e-06 
0.0 -0.3596 0 -2.0 1e-06 
0.0 -0.3595 0 -2.0 1e-06 
0.0 -0.3594 0 -2.0 1e-06 
0.0 -0.3593 0 -2.0 1e-06 
0.0 -0.3592 0 -2.0 1e-06 
0.0 -0.3591 0 -2.0 1e-06 
0.0 -0.359 0 -2.0 1e-06 
0.0 -0.3589 0 -2.0 1e-06 
0.0 -0.3588 0 -2.0 1e-06 
0.0 -0.3587 0 -2.0 1e-06 
0.0 -0.3586 0 -2.0 1e-06 
0.0 -0.3585 0 -2.0 1e-06 
0.0 -0.3584 0 -2.0 1e-06 
0.0 -0.3583 0 -2.0 1e-06 
0.0 -0.3582 0 -2.0 1e-06 
0.0 -0.3581 0 -2.0 1e-06 
0.0 -0.358 0 -2.0 1e-06 
0.0 -0.3579 0 -2.0 1e-06 
0.0 -0.3578 0 -2.0 1e-06 
0.0 -0.3577 0 -2.0 1e-06 
0.0 -0.3576 0 -2.0 1e-06 
0.0 -0.3575 0 -2.0 1e-06 
0.0 -0.3574 0 -2.0 1e-06 
0.0 -0.3573 0 -2.0 1e-06 
0.0 -0.3572 0 -2.0 1e-06 
0.0 -0.3571 0 -2.0 1e-06 
0.0 -0.357 0 -2.0 1e-06 
0.0 -0.3569 0 -2.0 1e-06 
0.0 -0.3568 0 -2.0 1e-06 
0.0 -0.3567 0 -2.0 1e-06 
0.0 -0.3566 0 -2.0 1e-06 
0.0 -0.3565 0 -2.0 1e-06 
0.0 -0.3564 0 -2.0 1e-06 
0.0 -0.3563 0 -2.0 1e-06 
0.0 -0.3562 0 -2.0 1e-06 
0.0 -0.3561 0 -2.0 1e-06 
0.0 -0.356 0 -2.0 1e-06 
0.0 -0.3559 0 -2.0 1e-06 
0.0 -0.3558 0 -2.0 1e-06 
0.0 -0.3557 0 -2.0 1e-06 
0.0 -0.3556 0 -2.0 1e-06 
0.0 -0.3555 0 -2.0 1e-06 
0.0 -0.3554 0 -2.0 1e-06 
0.0 -0.3553 0 -2.0 1e-06 
0.0 -0.3552 0 -2.0 1e-06 
0.0 -0.3551 0 -2.0 1e-06 
0.0 -0.355 0 -2.0 1e-06 
0.0 -0.3549 0 -2.0 1e-06 
0.0 -0.3548 0 -2.0 1e-06 
0.0 -0.3547 0 -2.0 1e-06 
0.0 -0.3546 0 -2.0 1e-06 
0.0 -0.3545 0 -2.0 1e-06 
0.0 -0.3544 0 -2.0 1e-06 
0.0 -0.3543 0 -2.0 1e-06 
0.0 -0.3542 0 -2.0 1e-06 
0.0 -0.3541 0 -2.0 1e-06 
0.0 -0.354 0 -2.0 1e-06 
0.0 -0.3539 0 -2.0 1e-06 
0.0 -0.3538 0 -2.0 1e-06 
0.0 -0.3537 0 -2.0 1e-06 
0.0 -0.3536 0 -2.0 1e-06 
0.0 -0.3535 0 -2.0 1e-06 
0.0 -0.3534 0 -2.0 1e-06 
0.0 -0.3533 0 -2.0 1e-06 
0.0 -0.3532 0 -2.0 1e-06 
0.0 -0.3531 0 -2.0 1e-06 
0.0 -0.353 0 -2.0 1e-06 
0.0 -0.3529 0 -2.0 1e-06 
0.0 -0.3528 0 -2.0 1e-06 
0.0 -0.3527 0 -2.0 1e-06 
0.0 -0.3526 0 -2.0 1e-06 
0.0 -0.3525 0 -2.0 1e-06 
0.0 -0.3524 0 -2.0 1e-06 
0.0 -0.3523 0 -2.0 1e-06 
0.0 -0.3522 0 -2.0 1e-06 
0.0 -0.3521 0 -2.0 1e-06 
0.0 -0.352 0 -2.0 1e-06 
0.0 -0.3519 0 -2.0 1e-06 
0.0 -0.3518 0 -2.0 1e-06 
0.0 -0.3517 0 -2.0 1e-06 
0.0 -0.3516 0 -2.0 1e-06 
0.0 -0.3515 0 -2.0 1e-06 
0.0 -0.3514 0 -2.0 1e-06 
0.0 -0.3513 0 -2.0 1e-06 
0.0 -0.3512 0 -2.0 1e-06 
0.0 -0.3511 0 -2.0 1e-06 
0.0 -0.351 0 -2.0 1e-06 
0.0 -0.3509 0 -2.0 1e-06 
0.0 -0.3508 0 -2.0 1e-06 
0.0 -0.3507 0 -2.0 1e-06 
0.0 -0.3506 0 -2.0 1e-06 
0.0 -0.3505 0 -2.0 1e-06 
0.0 -0.3504 0 -2.0 1e-06 
0.0 -0.3503 0 -2.0 1e-06 
0.0 -0.3502 0 -2.0 1e-06 
0.0 -0.3501 0 -2.0 1e-06 
0.0 -0.35 0 -2.0 1e-06 
0.0 -0.3499 0 -2.0 1e-06 
0.0 -0.3498 0 -2.0 1e-06 
0.0 -0.3497 0 -2.0 1e-06 
0.0 -0.3496 0 -2.0 1e-06 
0.0 -0.3495 0 -2.0 1e-06 
0.0 -0.3494 0 -2.0 1e-06 
0.0 -0.3493 0 -2.0 1e-06 
0.0 -0.3492 0 -2.0 1e-06 
0.0 -0.3491 0 -2.0 1e-06 
0.0 -0.349 0 -2.0 1e-06 
0.0 -0.3489 0 -2.0 1e-06 
0.0 -0.3488 0 -2.0 1e-06 
0.0 -0.3487 0 -2.0 1e-06 
0.0 -0.3486 0 -2.0 1e-06 
0.0 -0.3485 0 -2.0 1e-06 
0.0 -0.3484 0 -2.0 1e-06 
0.0 -0.3483 0 -2.0 1e-06 
0.0 -0.3482 0 -2.0 1e-06 
0.0 -0.3481 0 -2.0 1e-06 
0.0 -0.348 0 -2.0 1e-06 
0.0 -0.3479 0 -2.0 1e-06 
0.0 -0.3478 0 -2.0 1e-06 
0.0 -0.3477 0 -2.0 1e-06 
0.0 -0.3476 0 -2.0 1e-06 
0.0 -0.3475 0 -2.0 1e-06 
0.0 -0.3474 0 -2.0 1e-06 
0.0 -0.3473 0 -2.0 1e-06 
0.0 -0.3472 0 -2.0 1e-06 
0.0 -0.3471 0 -2.0 1e-06 
0.0 -0.347 0 -2.0 1e-06 
0.0 -0.3469 0 -2.0 1e-06 
0.0 -0.3468 0 -2.0 1e-06 
0.0 -0.3467 0 -2.0 1e-06 
0.0 -0.3466 0 -2.0 1e-06 
0.0 -0.3465 0 -2.0 1e-06 
0.0 -0.3464 0 -2.0 1e-06 
0.0 -0.3463 0 -2.0 1e-06 
0.0 -0.3462 0 -2.0 1e-06 
0.0 -0.3461 0 -2.0 1e-06 
0.0 -0.346 0 -2.0 1e-06 
0.0 -0.3459 0 -2.0 1e-06 
0.0 -0.3458 0 -2.0 1e-06 
0.0 -0.3457 0 -2.0 1e-06 
0.0 -0.3456 0 -2.0 1e-06 
0.0 -0.3455 0 -2.0 1e-06 
0.0 -0.3454 0 -2.0 1e-06 
0.0 -0.3453 0 -2.0 1e-06 
0.0 -0.3452 0 -2.0 1e-06 
0.0 -0.3451 0 -2.0 1e-06 
0.0 -0.345 0 -2.0 1e-06 
0.0 -0.3449 0 -2.0 1e-06 
0.0 -0.3448 0 -2.0 1e-06 
0.0 -0.3447 0 -2.0 1e-06 
0.0 -0.3446 0 -2.0 1e-06 
0.0 -0.3445 0 -2.0 1e-06 
0.0 -0.3444 0 -2.0 1e-06 
0.0 -0.3443 0 -2.0 1e-06 
0.0 -0.3442 0 -2.0 1e-06 
0.0 -0.3441 0 -2.0 1e-06 
0.0 -0.344 0 -2.0 1e-06 
0.0 -0.3439 0 -2.0 1e-06 
0.0 -0.3438 0 -2.0 1e-06 
0.0 -0.3437 0 -2.0 1e-06 
0.0 -0.3436 0 -2.0 1e-06 
0.0 -0.3435 0 -2.0 1e-06 
0.0 -0.3434 0 -2.0 1e-06 
0.0 -0.3433 0 -2.0 1e-06 
0.0 -0.3432 0 -2.0 1e-06 
0.0 -0.3431 0 -2.0 1e-06 
0.0 -0.343 0 -2.0 1e-06 
0.0 -0.3429 0 -2.0 1e-06 
0.0 -0.3428 0 -2.0 1e-06 
0.0 -0.3427 0 -2.0 1e-06 
0.0 -0.3426 0 -2.0 1e-06 
0.0 -0.3425 0 -2.0 1e-06 
0.0 -0.3424 0 -2.0 1e-06 
0.0 -0.3423 0 -2.0 1e-06 
0.0 -0.3422 0 -2.0 1e-06 
0.0 -0.3421 0 -2.0 1e-06 
0.0 -0.342 0 -2.0 1e-06 
0.0 -0.3419 0 -2.0 1e-06 
0.0 -0.3418 0 -2.0 1e-06 
0.0 -0.3417 0 -2.0 1e-06 
0.0 -0.3416 0 -2.0 1e-06 
0.0 -0.3415 0 -2.0 1e-06 
0.0 -0.3414 0 -2.0 1e-06 
0.0 -0.3413 0 -2.0 1e-06 
0.0 -0.3412 0 -2.0 1e-06 
0.0 -0.3411 0 -2.0 1e-06 
0.0 -0.341 0 -2.0 1e-06 
0.0 -0.3409 0 -2.0 1e-06 
0.0 -0.3408 0 -2.0 1e-06 
0.0 -0.3407 0 -2.0 1e-06 
0.0 -0.3406 0 -2.0 1e-06 
0.0 -0.3405 0 -2.0 1e-06 
0.0 -0.3404 0 -2.0 1e-06 
0.0 -0.3403 0 -2.0 1e-06 
0.0 -0.3402 0 -2.0 1e-06 
0.0 -0.3401 0 -2.0 1e-06 
0.0 -0.34 0 -2.0 1e-06 
0.0 -0.3399 0 -2.0 1e-06 
0.0 -0.3398 0 -2.0 1e-06 
0.0 -0.3397 0 -2.0 1e-06 
0.0 -0.3396 0 -2.0 1e-06 
0.0 -0.3395 0 -2.0 1e-06 
0.0 -0.3394 0 -2.0 1e-06 
0.0 -0.3393 0 -2.0 1e-06 
0.0 -0.3392 0 -2.0 1e-06 
0.0 -0.3391 0 -2.0 1e-06 
0.0 -0.339 0 -2.0 1e-06 
0.0 -0.3389 0 -2.0 1e-06 
0.0 -0.3388 0 -2.0 1e-06 
0.0 -0.3387 0 -2.0 1e-06 
0.0 -0.3386 0 -2.0 1e-06 
0.0 -0.3385 0 -2.0 1e-06 
0.0 -0.3384 0 -2.0 1e-06 
0.0 -0.3383 0 -2.0 1e-06 
0.0 -0.3382 0 -2.0 1e-06 
0.0 -0.3381 0 -2.0 1e-06 
0.0 -0.338 0 -2.0 1e-06 
0.0 -0.3379 0 -2.0 1e-06 
0.0 -0.3378 0 -2.0 1e-06 
0.0 -0.3377 0 -2.0 1e-06 
0.0 -0.3376 0 -2.0 1e-06 
0.0 -0.3375 0 -2.0 1e-06 
0.0 -0.3374 0 -2.0 1e-06 
0.0 -0.3373 0 -2.0 1e-06 
0.0 -0.3372 0 -2.0 1e-06 
0.0 -0.3371 0 -2.0 1e-06 
0.0 -0.337 0 -2.0 1e-06 
0.0 -0.3369 0 -2.0 1e-06 
0.0 -0.3368 0 -2.0 1e-06 
0.0 -0.3367 0 -2.0 1e-06 
0.0 -0.3366 0 -2.0 1e-06 
0.0 -0.3365 0 -2.0 1e-06 
0.0 -0.3364 0 -2.0 1e-06 
0.0 -0.3363 0 -2.0 1e-06 
0.0 -0.3362 0 -2.0 1e-06 
0.0 -0.3361 0 -2.0 1e-06 
0.0 -0.336 0 -2.0 1e-06 
0.0 -0.3359 0 -2.0 1e-06 
0.0 -0.3358 0 -2.0 1e-06 
0.0 -0.3357 0 -2.0 1e-06 
0.0 -0.3356 0 -2.0 1e-06 
0.0 -0.3355 0 -2.0 1e-06 
0.0 -0.3354 0 -2.0 1e-06 
0.0 -0.3353 0 -2.0 1e-06 
0.0 -0.3352 0 -2.0 1e-06 
0.0 -0.3351 0 -2.0 1e-06 
0.0 -0.335 0 -2.0 1e-06 
0.0 -0.3349 0 -2.0 1e-06 
0.0 -0.3348 0 -2.0 1e-06 
0.0 -0.3347 0 -2.0 1e-06 
0.0 -0.3346 0 -2.0 1e-06 
0.0 -0.3345 0 -2.0 1e-06 
0.0 -0.3344 0 -2.0 1e-06 
0.0 -0.3343 0 -2.0 1e-06 
0.0 -0.3342 0 -2.0 1e-06 
0.0 -0.3341 0 -2.0 1e-06 
0.0 -0.334 0 -2.0 1e-06 
0.0 -0.3339 0 -2.0 1e-06 
0.0 -0.3338 0 -2.0 1e-06 
0.0 -0.3337 0 -2.0 1e-06 
0.0 -0.3336 0 -2.0 1e-06 
0.0 -0.3335 0 -2.0 1e-06 
0.0 -0.3334 0 -2.0 1e-06 
0.0 -0.3333 0 -2.0 1e-06 
0.0 -0.3332 0 -2.0 1e-06 
0.0 -0.3331 0 -2.0 1e-06 
0.0 -0.333 0 -2.0 1e-06 
0.0 -0.3329 0 -2.0 1e-06 
0.0 -0.3328 0 -2.0 1e-06 
0.0 -0.3327 0 -2.0 1e-06 
0.0 -0.3326 0 -2.0 1e-06 
0.0 -0.3325 0 -2.0 1e-06 
0.0 -0.3324 0 -2.0 1e-06 
0.0 -0.3323 0 -2.0 1e-06 
0.0 -0.3322 0 -2.0 1e-06 
0.0 -0.3321 0 -2.0 1e-06 
0.0 -0.332 0 -2.0 1e-06 
0.0 -0.3319 0 -2.0 1e-06 
0.0 -0.3318 0 -2.0 1e-06 
0.0 -0.3317 0 -2.0 1e-06 
0.0 -0.3316 0 -2.0 1e-06 
0.0 -0.3315 0 -2.0 1e-06 
0.0 -0.3314 0 -2.0 1e-06 
0.0 -0.3313 0 -2.0 1e-06 
0.0 -0.3312 0 -2.0 1e-06 
0.0 -0.3311 0 -2.0 1e-06 
0.0 -0.331 0 -2.0 1e-06 
0.0 -0.3309 0 -2.0 1e-06 
0.0 -0.3308 0 -2.0 1e-06 
0.0 -0.3307 0 -2.0 1e-06 
0.0 -0.3306 0 -2.0 1e-06 
0.0 -0.3305 0 -2.0 1e-06 
0.0 -0.3304 0 -2.0 1e-06 
0.0 -0.3303 0 -2.0 1e-06 
0.0 -0.3302 0 -2.0 1e-06 
0.0 -0.3301 0 -2.0 1e-06 
0.0 -0.33 0 -2.0 1e-06 
0.0 -0.3299 0 -2.0 1e-06 
0.0 -0.3298 0 -2.0 1e-06 
0.0 -0.3297 0 -2.0 1e-06 
0.0 -0.3296 0 -2.0 1e-06 
0.0 -0.3295 0 -2.0 1e-06 
0.0 -0.3294 0 -2.0 1e-06 
0.0 -0.3293 0 -2.0 1e-06 
0.0 -0.3292 0 -2.0 1e-06 
0.0 -0.3291 0 -2.0 1e-06 
0.0 -0.329 0 -2.0 1e-06 
0.0 -0.3289 0 -2.0 1e-06 
0.0 -0.3288 0 -2.0 1e-06 
0.0 -0.3287 0 -2.0 1e-06 
0.0 -0.3286 0 -2.0 1e-06 
0.0 -0.3285 0 -2.0 1e-06 
0.0 -0.3284 0 -2.0 1e-06 
0.0 -0.3283 0 -2.0 1e-06 
0.0 -0.3282 0 -2.0 1e-06 
0.0 -0.3281 0 -2.0 1e-06 
0.0 -0.328 0 -2.0 1e-06 
0.0 -0.3279 0 -2.0 1e-06 
0.0 -0.3278 0 -2.0 1e-06 
0.0 -0.3277 0 -2.0 1e-06 
0.0 -0.3276 0 -2.0 1e-06 
0.0 -0.3275 0 -2.0 1e-06 
0.0 -0.3274 0 -2.0 1e-06 
0.0 -0.3273 0 -2.0 1e-06 
0.0 -0.3272 0 -2.0 1e-06 
0.0 -0.3271 0 -2.0 1e-06 
0.0 -0.327 0 -2.0 1e-06 
0.0 -0.3269 0 -2.0 1e-06 
0.0 -0.3268 0 -2.0 1e-06 
0.0 -0.3267 0 -2.0 1e-06 
0.0 -0.3266 0 -2.0 1e-06 
0.0 -0.3265 0 -2.0 1e-06 
0.0 -0.3264 0 -2.0 1e-06 
0.0 -0.3263 0 -2.0 1e-06 
0.0 -0.3262 0 -2.0 1e-06 
0.0 -0.3261 0 -2.0 1e-06 
0.0 -0.326 0 -2.0 1e-06 
0.0 -0.3259 0 -2.0 1e-06 
0.0 -0.3258 0 -2.0 1e-06 
0.0 -0.3257 0 -2.0 1e-06 
0.0 -0.3256 0 -2.0 1e-06 
0.0 -0.3255 0 -2.0 1e-06 
0.0 -0.3254 0 -2.0 1e-06 
0.0 -0.3253 0 -2.0 1e-06 
0.0 -0.3252 0 -2.0 1e-06 
0.0 -0.3251 0 -2.0 1e-06 
0.0 -0.325 0 -2.0 1e-06 
0.0 -0.3249 0 -2.0 1e-06 
0.0 -0.3248 0 -2.0 1e-06 
0.0 -0.3247 0 -2.0 1e-06 
0.0 -0.3246 0 -2.0 1e-06 
0.0 -0.3245 0 -2.0 1e-06 
0.0 -0.3244 0 -2.0 1e-06 
0.0 -0.3243 0 -2.0 1e-06 
0.0 -0.3242 0 -2.0 1e-06 
0.0 -0.3241 0 -2.0 1e-06 
0.0 -0.324 0 -2.0 1e-06 
0.0 -0.3239 0 -2.0 1e-06 
0.0 -0.3238 0 -2.0 1e-06 
0.0 -0.3237 0 -2.0 1e-06 
0.0 -0.3236 0 -2.0 1e-06 
0.0 -0.3235 0 -2.0 1e-06 
0.0 -0.3234 0 -2.0 1e-06 
0.0 -0.3233 0 -2.0 1e-06 
0.0 -0.3232 0 -2.0 1e-06 
0.0 -0.3231 0 -2.0 1e-06 
0.0 -0.323 0 -2.0 1e-06 
0.0 -0.3229 0 -2.0 1e-06 
0.0 -0.3228 0 -2.0 1e-06 
0.0 -0.3227 0 -2.0 1e-06 
0.0 -0.3226 0 -2.0 1e-06 
0.0 -0.3225 0 -2.0 1e-06 
0.0 -0.3224 0 -2.0 1e-06 
0.0 -0.3223 0 -2.0 1e-06 
0.0 -0.3222 0 -2.0 1e-06 
0.0 -0.3221 0 -2.0 1e-06 
0.0 -0.322 0 -2.0 1e-06 
0.0 -0.3219 0 -2.0 1e-06 
0.0 -0.3218 0 -2.0 1e-06 
0.0 -0.3217 0 -2.0 1e-06 
0.0 -0.3216 0 -2.0 1e-06 
0.0 -0.3215 0 -2.0 1e-06 
0.0 -0.3214 0 -2.0 1e-06 
0.0 -0.3213 0 -2.0 1e-06 
0.0 -0.3212 0 -2.0 1e-06 
0.0 -0.3211 0 -2.0 1e-06 
0.0 -0.321 0 -2.0 1e-06 
0.0 -0.3209 0 -2.0 1e-06 
0.0 -0.3208 0 -2.0 1e-06 
0.0 -0.3207 0 -2.0 1e-06 
0.0 -0.3206 0 -2.0 1e-06 
0.0 -0.3205 0 -2.0 1e-06 
0.0 -0.3204 0 -2.0 1e-06 
0.0 -0.3203 0 -2.0 1e-06 
0.0 -0.3202 0 -2.0 1e-06 
0.0 -0.3201 0 -2.0 1e-06 
0.0 -0.32 0 -2.0 1e-06 
0.0 -0.3199 0 -2.0 1e-06 
0.0 -0.3198 0 -2.0 1e-06 
0.0 -0.3197 0 -2.0 1e-06 
0.0 -0.3196 0 -2.0 1e-06 
0.0 -0.3195 0 -2.0 1e-06 
0.0 -0.3194 0 -2.0 1e-06 
0.0 -0.3193 0 -2.0 1e-06 
0.0 -0.3192 0 -2.0 1e-06 
0.0 -0.3191 0 -2.0 1e-06 
0.0 -0.319 0 -2.0 1e-06 
0.0 -0.3189 0 -2.0 1e-06 
0.0 -0.3188 0 -2.0 1e-06 
0.0 -0.3187 0 -2.0 1e-06 
0.0 -0.3186 0 -2.0 1e-06 
0.0 -0.3185 0 -2.0 1e-06 
0.0 -0.3184 0 -2.0 1e-06 
0.0 -0.3183 0 -2.0 1e-06 
0.0 -0.3182 0 -2.0 1e-06 
0.0 -0.3181 0 -2.0 1e-06 
0.0 -0.318 0 -2.0 1e-06 
0.0 -0.3179 0 -2.0 1e-06 
0.0 -0.3178 0 -2.0 1e-06 
0.0 -0.3177 0 -2.0 1e-06 
0.0 -0.3176 0 -2.0 1e-06 
0.0 -0.3175 0 -2.0 1e-06 
0.0 -0.3174 0 -2.0 1e-06 
0.0 -0.3173 0 -2.0 1e-06 
0.0 -0.3172 0 -2.0 1e-06 
0.0 -0.3171 0 -2.0 1e-06 
0.0 -0.317 0 -2.0 1e-06 
0.0 -0.3169 0 -2.0 1e-06 
0.0 -0.3168 0 -2.0 1e-06 
0.0 -0.3167 0 -2.0 1e-06 
0.0 -0.3166 0 -2.0 1e-06 
0.0 -0.3165 0 -2.0 1e-06 
0.0 -0.3164 0 -2.0 1e-06 
0.0 -0.3163 0 -2.0 1e-06 
0.0 -0.3162 0 -2.0 1e-06 
0.0 -0.3161 0 -2.0 1e-06 
0.0 -0.316 0 -2.0 1e-06 
0.0 -0.3159 0 -2.0 1e-06 
0.0 -0.3158 0 -2.0 1e-06 
0.0 -0.3157 0 -2.0 1e-06 
0.0 -0.3156 0 -2.0 1e-06 
0.0 -0.3155 0 -2.0 1e-06 
0.0 -0.3154 0 -2.0 1e-06 
0.0 -0.3153 0 -2.0 1e-06 
0.0 -0.3152 0 -2.0 1e-06 
0.0 -0.3151 0 -2.0 1e-06 
0.0 -0.315 0 -2.0 1e-06 
0.0 -0.3149 0 -2.0 1e-06 
0.0 -0.3148 0 -2.0 1e-06 
0.0 -0.3147 0 -2.0 1e-06 
0.0 -0.3146 0 -2.0 1e-06 
0.0 -0.3145 0 -2.0 1e-06 
0.0 -0.3144 0 -2.0 1e-06 
0.0 -0.3143 0 -2.0 1e-06 
0.0 -0.3142 0 -2.0 1e-06 
0.0 -0.3141 0 -2.0 1e-06 
0.0 -0.314 0 -2.0 1e-06 
0.0 -0.3139 0 -2.0 1e-06 
0.0 -0.3138 0 -2.0 1e-06 
0.0 -0.3137 0 -2.0 1e-06 
0.0 -0.3136 0 -2.0 1e-06 
0.0 -0.3135 0 -2.0 1e-06 
0.0 -0.3134 0 -2.0 1e-06 
0.0 -0.3133 0 -2.0 1e-06 
0.0 -0.3132 0 -2.0 1e-06 
0.0 -0.3131 0 -2.0 1e-06 
0.0 -0.313 0 -2.0 1e-06 
0.0 -0.3129 0 -2.0 1e-06 
0.0 -0.3128 0 -2.0 1e-06 
0.0 -0.3127 0 -2.0 1e-06 
0.0 -0.3126 0 -2.0 1e-06 
0.0 -0.3125 0 -2.0 1e-06 
0.0 -0.3124 0 -2.0 1e-06 
0.0 -0.3123 0 -2.0 1e-06 
0.0 -0.3122 0 -2.0 1e-06 
0.0 -0.3121 0 -2.0 1e-06 
0.0 -0.312 0 -2.0 1e-06 
0.0 -0.3119 0 -2.0 1e-06 
0.0 -0.3118 0 -2.0 1e-06 
0.0 -0.3117 0 -2.0 1e-06 
0.0 -0.3116 0 -2.0 1e-06 
0.0 -0.3115 0 -2.0 1e-06 
0.0 -0.3114 0 -2.0 1e-06 
0.0 -0.3113 0 -2.0 1e-06 
0.0 -0.3112 0 -2.0 1e-06 
0.0 -0.3111 0 -2.0 1e-06 
0.0 -0.311 0 -2.0 1e-06 
0.0 -0.3109 0 -2.0 1e-06 
0.0 -0.3108 0 -2.0 1e-06 
0.0 -0.3107 0 -2.0 1e-06 
0.0 -0.3106 0 -2.0 1e-06 
0.0 -0.3105 0 -2.0 1e-06 
0.0 -0.3104 0 -2.0 1e-06 
0.0 -0.3103 0 -2.0 1e-06 
0.0 -0.3102 0 -2.0 1e-06 
0.0 -0.3101 0 -2.0 1e-06 
0.0 -0.31 0 -2.0 1e-06 
0.0 -0.3099 0 -2.0 1e-06 
0.0 -0.3098 0 -2.0 1e-06 
0.0 -0.3097 0 -2.0 1e-06 
0.0 -0.3096 0 -2.0 1e-06 
0.0 -0.3095 0 -2.0 1e-06 
0.0 -0.3094 0 -2.0 1e-06 
0.0 -0.3093 0 -2.0 1e-06 
0.0 -0.3092 0 -2.0 1e-06 
0.0 -0.3091 0 -2.0 1e-06 
0.0 -0.309 0 -2.0 1e-06 
0.0 -0.3089 0 -2.0 1e-06 
0.0 -0.3088 0 -2.0 1e-06 
0.0 -0.3087 0 -2.0 1e-06 
0.0 -0.3086 0 -2.0 1e-06 
0.0 -0.3085 0 -2.0 1e-06 
0.0 -0.3084 0 -2.0 1e-06 
0.0 -0.3083 0 -2.0 1e-06 
0.0 -0.3082 0 -2.0 1e-06 
0.0 -0.3081 0 -2.0 1e-06 
0.0 -0.308 0 -2.0 1e-06 
0.0 -0.3079 0 -2.0 1e-06 
0.0 -0.3078 0 -2.0 1e-06 
0.0 -0.3077 0 -2.0 1e-06 
0.0 -0.3076 0 -2.0 1e-06 
0.0 -0.3075 0 -2.0 1e-06 
0.0 -0.3074 0 -2.0 1e-06 
0.0 -0.3073 0 -2.0 1e-06 
0.0 -0.3072 0 -2.0 1e-06 
0.0 -0.3071 0 -2.0 1e-06 
0.0 -0.307 0 -2.0 1e-06 
0.0 -0.3069 0 -2.0 1e-06 
0.0 -0.3068 0 -2.0 1e-06 
0.0 -0.3067 0 -2.0 1e-06 
0.0 -0.3066 0 -2.0 1e-06 
0.0 -0.3065 0 -2.0 1e-06 
0.0 -0.3064 0 -2.0 1e-06 
0.0 -0.3063 0 -2.0 1e-06 
0.0 -0.3062 0 -2.0 1e-06 
0.0 -0.3061 0 -2.0 1e-06 
0.0 -0.306 0 -2.0 1e-06 
0.0 -0.3059 0 -2.0 1e-06 
0.0 -0.3058 0 -2.0 1e-06 
0.0 -0.3057 0 -2.0 1e-06 
0.0 -0.3056 0 -2.0 1e-06 
0.0 -0.3055 0 -2.0 1e-06 
0.0 -0.3054 0 -2.0 1e-06 
0.0 -0.3053 0 -2.0 1e-06 
0.0 -0.3052 0 -2.0 1e-06 
0.0 -0.3051 0 -2.0 1e-06 
0.0 -0.305 0 -2.0 1e-06 
0.0 -0.3049 0 -2.0 1e-06 
0.0 -0.3048 0 -2.0 1e-06 
0.0 -0.3047 0 -2.0 1e-06 
0.0 -0.3046 0 -2.0 1e-06 
0.0 -0.3045 0 -2.0 1e-06 
0.0 -0.3044 0 -2.0 1e-06 
0.0 -0.3043 0 -2.0 1e-06 
0.0 -0.3042 0 -2.0 1e-06 
0.0 -0.3041 0 -2.0 1e-06 
0.0 -0.304 0 -2.0 1e-06 
0.0 -0.3039 0 -2.0 1e-06 
0.0 -0.3038 0 -2.0 1e-06 
0.0 -0.3037 0 -2.0 1e-06 
0.0 -0.3036 0 -2.0 1e-06 
0.0 -0.3035 0 -2.0 1e-06 
0.0 -0.3034 0 -2.0 1e-06 
0.0 -0.3033 0 -2.0 1e-06 
0.0 -0.3032 0 -2.0 1e-06 
0.0 -0.3031 0 -2.0 1e-06 
0.0 -0.303 0 -2.0 1e-06 
0.0 -0.3029 0 -2.0 1e-06 
0.0 -0.3028 0 -2.0 1e-06 
0.0 -0.3027 0 -2.0 1e-06 
0.0 -0.3026 0 -2.0 1e-06 
0.0 -0.3025 0 -2.0 1e-06 
0.0 -0.3024 0 -2.0 1e-06 
0.0 -0.3023 0 -2.0 1e-06 
0.0 -0.3022 0 -2.0 1e-06 
0.0 -0.3021 0 -2.0 1e-06 
0.0 -0.302 0 -2.0 1e-06 
0.0 -0.3019 0 -2.0 1e-06 
0.0 -0.3018 0 -2.0 1e-06 
0.0 -0.3017 0 -2.0 1e-06 
0.0 -0.3016 0 -2.0 1e-06 
0.0 -0.3015 0 -2.0 1e-06 
0.0 -0.3014 0 -2.0 1e-06 
0.0 -0.3013 0 -2.0 1e-06 
0.0 -0.3012 0 -2.0 1e-06 
0.0 -0.3011 0 -2.0 1e-06 
0.0 -0.301 0 -2.0 1e-06 
0.0 -0.3009 0 -2.0 1e-06 
0.0 -0.3008 0 -2.0 1e-06 
0.0 -0.3007 0 -2.0 1e-06 
0.0 -0.3006 0 -2.0 1e-06 
0.0 -0.3005 0 -2.0 1e-06 
0.0 -0.3004 0 -2.0 1e-06 
0.0 -0.3003 0 -2.0 1e-06 
0.0 -0.3002 0 -2.0 1e-06 
0.0 -0.3001 0 -2.0 1e-06 
0.0 -0.3 0 -2.0 1e-06 
0.0 -0.2999 0 -2.0 1e-06 
0.0 -0.2998 0 -2.0 1e-06 
0.0 -0.2997 0 -2.0 1e-06 
0.0 -0.2996 0 -2.0 1e-06 
0.0 -0.2995 0 -2.0 1e-06 
0.0 -0.2994 0 -2.0 1e-06 
0.0 -0.2993 0 -2.0 1e-06 
0.0 -0.2992 0 -2.0 1e-06 
0.0 -0.2991 0 -2.0 1e-06 
0.0 -0.299 0 -2.0 1e-06 
0.0 -0.2989 0 -2.0 1e-06 
0.0 -0.2988 0 -2.0 1e-06 
0.0 -0.2987 0 -2.0 1e-06 
0.0 -0.2986 0 -2.0 1e-06 
0.0 -0.2985 0 -2.0 1e-06 
0.0 -0.2984 0 -2.0 1e-06 
0.0 -0.2983 0 -2.0 1e-06 
0.0 -0.2982 0 -2.0 1e-06 
0.0 -0.2981 0 -2.0 1e-06 
0.0 -0.298 0 -2.0 1e-06 
0.0 -0.2979 0 -2.0 1e-06 
0.0 -0.2978 0 -2.0 1e-06 
0.0 -0.2977 0 -2.0 1e-06 
0.0 -0.2976 0 -2.0 1e-06 
0.0 -0.2975 0 -2.0 1e-06 
0.0 -0.2974 0 -2.0 1e-06 
0.0 -0.2973 0 -2.0 1e-06 
0.0 -0.2972 0 -2.0 1e-06 
0.0 -0.2971 0 -2.0 1e-06 
0.0 -0.297 0 -2.0 1e-06 
0.0 -0.2969 0 -2.0 1e-06 
0.0 -0.2968 0 -2.0 1e-06 
0.0 -0.2967 0 -2.0 1e-06 
0.0 -0.2966 0 -2.0 1e-06 
0.0 -0.2965 0 -2.0 1e-06 
0.0 -0.2964 0 -2.0 1e-06 
0.0 -0.2963 0 -2.0 1e-06 
0.0 -0.2962 0 -2.0 1e-06 
0.0 -0.2961 0 -2.0 1e-06 
0.0 -0.296 0 -2.0 1e-06 
0.0 -0.2959 0 -2.0 1e-06 
0.0 -0.2958 0 -2.0 1e-06 
0.0 -0.2957 0 -2.0 1e-06 
0.0 -0.2956 0 -2.0 1e-06 
0.0 -0.2955 0 -2.0 1e-06 
0.0 -0.2954 0 -2.0 1e-06 
0.0 -0.2953 0 -2.0 1e-06 
0.0 -0.2952 0 -2.0 1e-06 
0.0 -0.2951 0 -2.0 1e-06 
0.0 -0.295 0 -2.0 1e-06 
0.0 -0.2949 0 -2.0 1e-06 
0.0 -0.2948 0 -2.0 1e-06 
0.0 -0.2947 0 -2.0 1e-06 
0.0 -0.2946 0 -2.0 1e-06 
0.0 -0.2945 0 -2.0 1e-06 
0.0 -0.2944 0 -2.0 1e-06 
0.0 -0.2943 0 -2.0 1e-06 
0.0 -0.2942 0 -2.0 1e-06 
0.0 -0.2941 0 -2.0 1e-06 
0.0 -0.294 0 -2.0 1e-06 
0.0 -0.2939 0 -2.0 1e-06 
0.0 -0.2938 0 -2.0 1e-06 
0.0 -0.2937 0 -2.0 1e-06 
0.0 -0.2936 0 -2.0 1e-06 
0.0 -0.2935 0 -2.0 1e-06 
0.0 -0.2934 0 -2.0 1e-06 
0.0 -0.2933 0 -2.0 1e-06 
0.0 -0.2932 0 -2.0 1e-06 
0.0 -0.2931 0 -2.0 1e-06 
0.0 -0.293 0 -2.0 1e-06 
0.0 -0.2929 0 -2.0 1e-06 
0.0 -0.2928 0 -2.0 1e-06 
0.0 -0.2927 0 -2.0 1e-06 
0.0 -0.2926 0 -2.0 1e-06 
0.0 -0.2925 0 -2.0 1e-06 
0.0 -0.2924 0 -2.0 1e-06 
0.0 -0.2923 0 -2.0 1e-06 
0.0 -0.2922 0 -2.0 1e-06 
0.0 -0.2921 0 -2.0 1e-06 
0.0 -0.292 0 -2.0 1e-06 
0.0 -0.2919 0 -2.0 1e-06 
0.0 -0.2918 0 -2.0 1e-06 
0.0 -0.2917 0 -2.0 1e-06 
0.0 -0.2916 0 -2.0 1e-06 
0.0 -0.2915 0 -2.0 1e-06 
0.0 -0.2914 0 -2.0 1e-06 
0.0 -0.2913 0 -2.0 1e-06 
0.0 -0.2912 0 -2.0 1e-06 
0.0 -0.2911 0 -2.0 1e-06 
0.0 -0.291 0 -2.0 1e-06 
0.0 -0.2909 0 -2.0 1e-06 
0.0 -0.2908 0 -2.0 1e-06 
0.0 -0.2907 0 -2.0 1e-06 
0.0 -0.2906 0 -2.0 1e-06 
0.0 -0.2905 0 -2.0 1e-06 
0.0 -0.2904 0 -2.0 1e-06 
0.0 -0.2903 0 -2.0 1e-06 
0.0 -0.2902 0 -2.0 1e-06 
0.0 -0.2901 0 -2.0 1e-06 
0.0 -0.29 0 -2.0 1e-06 
0.0 -0.2899 0 -2.0 1e-06 
0.0 -0.2898 0 -2.0 1e-06 
0.0 -0.2897 0 -2.0 1e-06 
0.0 -0.2896 0 -2.0 1e-06 
0.0 -0.2895 0 -2.0 1e-06 
0.0 -0.2894 0 -2.0 1e-06 
0.0 -0.2893 0 -2.0 1e-06 
0.0 -0.2892 0 -2.0 1e-06 
0.0 -0.2891 0 -2.0 1e-06 
0.0 -0.289 0 -2.0 1e-06 
0.0 -0.2889 0 -2.0 1e-06 
0.0 -0.2888 0 -2.0 1e-06 
0.0 -0.2887 0 -2.0 1e-06 
0.0 -0.2886 0 -2.0 1e-06 
0.0 -0.2885 0 -2.0 1e-06 
0.0 -0.2884 0 -2.0 1e-06 
0.0 -0.2883 0 -2.0 1e-06 
0.0 -0.2882 0 -2.0 1e-06 
0.0 -0.2881 0 -2.0 1e-06 
0.0 -0.288 0 -2.0 1e-06 
0.0 -0.2879 0 -2.0 1e-06 
0.0 -0.2878 0 -2.0 1e-06 
0.0 -0.2877 0 -2.0 1e-06 
0.0 -0.2876 0 -2.0 1e-06 
0.0 -0.2875 0 -2.0 1e-06 
0.0 -0.2874 0 -2.0 1e-06 
0.0 -0.2873 0 -2.0 1e-06 
0.0 -0.2872 0 -2.0 1e-06 
0.0 -0.2871 0 -2.0 1e-06 
0.0 -0.287 0 -2.0 1e-06 
0.0 -0.2869 0 -2.0 1e-06 
0.0 -0.2868 0 -2.0 1e-06 
0.0 -0.2867 0 -2.0 1e-06 
0.0 -0.2866 0 -2.0 1e-06 
0.0 -0.2865 0 -2.0 1e-06 
0.0 -0.2864 0 -2.0 1e-06 
0.0 -0.2863 0 -2.0 1e-06 
0.0 -0.2862 0 -2.0 1e-06 
0.0 -0.2861 0 -2.0 1e-06 
0.0 -0.286 0 -2.0 1e-06 
0.0 -0.2859 0 -2.0 1e-06 
0.0 -0.2858 0 -2.0 1e-06 
0.0 -0.2857 0 -2.0 1e-06 
0.0 -0.2856 0 -2.0 1e-06 
0.0 -0.2855 0 -2.0 1e-06 
0.0 -0.2854 0 -2.0 1e-06 
0.0 -0.2853 0 -2.0 1e-06 
0.0 -0.2852 0 -2.0 1e-06 
0.0 -0.2851 0 -2.0 1e-06 
0.0 -0.285 0 -2.0 1e-06 
0.0 -0.2849 0 -2.0 1e-06 
0.0 -0.2848 0 -2.0 1e-06 
0.0 -0.2847 0 -2.0 1e-06 
0.0 -0.2846 0 -2.0 1e-06 
0.0 -0.2845 0 -2.0 1e-06 
0.0 -0.2844 0 -2.0 1e-06 
0.0 -0.2843 0 -2.0 1e-06 
0.0 -0.2842 0 -2.0 1e-06 
0.0 -0.2841 0 -2.0 1e-06 
0.0 -0.284 0 -2.0 1e-06 
0.0 -0.2839 0 -2.0 1e-06 
0.0 -0.2838 0 -2.0 1e-06 
0.0 -0.2837 0 -2.0 1e-06 
0.0 -0.2836 0 -2.0 1e-06 
0.0 -0.2835 0 -2.0 1e-06 
0.0 -0.2834 0 -2.0 1e-06 
0.0 -0.2833 0 -2.0 1e-06 
0.0 -0.2832 0 -2.0 1e-06 
0.0 -0.2831 0 -2.0 1e-06 
0.0 -0.283 0 -2.0 1e-06 
0.0 -0.2829 0 -2.0 1e-06 
0.0 -0.2828 0 -2.0 1e-06 
0.0 -0.2827 0 -2.0 1e-06 
0.0 -0.2826 0 -2.0 1e-06 
0.0 -0.2825 0 -2.0 1e-06 
0.0 -0.2824 0 -2.0 1e-06 
0.0 -0.2823 0 -2.0 1e-06 
0.0 -0.2822 0 -2.0 1e-06 
0.0 -0.2821 0 -2.0 1e-06 
0.0 -0.282 0 -2.0 1e-06 
0.0 -0.2819 0 -2.0 1e-06 
0.0 -0.2818 0 -2.0 1e-06 
0.0 -0.2817 0 -2.0 1e-06 
0.0 -0.2816 0 -2.0 1e-06 
0.0 -0.2815 0 -2.0 1e-06 
0.0 -0.2814 0 -2.0 1e-06 
0.0 -0.2813 0 -2.0 1e-06 
0.0 -0.2812 0 -2.0 1e-06 
0.0 -0.2811 0 -2.0 1e-06 
0.0 -0.281 0 -2.0 1e-06 
0.0 -0.2809 0 -2.0 1e-06 
0.0 -0.2808 0 -2.0 1e-06 
0.0 -0.2807 0 -2.0 1e-06 
0.0 -0.2806 0 -2.0 1e-06 
0.0 -0.2805 0 -2.0 1e-06 
0.0 -0.2804 0 -2.0 1e-06 
0.0 -0.2803 0 -2.0 1e-06 
0.0 -0.2802 0 -2.0 1e-06 
0.0 -0.2801 0 -2.0 1e-06 
0.0 -0.28 0 -2.0 1e-06 
0.0 -0.2799 0 -2.0 1e-06 
0.0 -0.2798 0 -2.0 1e-06 
0.0 -0.2797 0 -2.0 1e-06 
0.0 -0.2796 0 -2.0 1e-06 
0.0 -0.2795 0 -2.0 1e-06 
0.0 -0.2794 0 -2.0 1e-06 
0.0 -0.2793 0 -2.0 1e-06 
0.0 -0.2792 0 -2.0 1e-06 
0.0 -0.2791 0 -2.0 1e-06 
0.0 -0.279 0 -2.0 1e-06 
0.0 -0.2789 0 -2.0 1e-06 
0.0 -0.2788 0 -2.0 1e-06 
0.0 -0.2787 0 -2.0 1e-06 
0.0 -0.2786 0 -2.0 1e-06 
0.0 -0.2785 0 -2.0 1e-06 
0.0 -0.2784 0 -2.0 1e-06 
0.0 -0.2783 0 -2.0 1e-06 
0.0 -0.2782 0 -2.0 1e-06 
0.0 -0.2781 0 -2.0 1e-06 
0.0 -0.278 0 -2.0 1e-06 
0.0 -0.2779 0 -2.0 1e-06 
0.0 -0.2778 0 -2.0 1e-06 
0.0 -0.2777 0 -2.0 1e-06 
0.0 -0.2776 0 -2.0 1e-06 
0.0 -0.2775 0 -2.0 1e-06 
0.0 -0.2774 0 -2.0 1e-06 
0.0 -0.2773 0 -2.0 1e-06 
0.0 -0.2772 0 -2.0 1e-06 
0.0 -0.2771 0 -2.0 1e-06 
0.0 -0.277 0 -2.0 1e-06 
0.0 -0.2769 0 -2.0 1e-06 
0.0 -0.2768 0 -2.0 1e-06 
0.0 -0.2767 0 -2.0 1e-06 
0.0 -0.2766 0 -2.0 1e-06 
0.0 -0.2765 0 -2.0 1e-06 
0.0 -0.2764 0 -2.0 1e-06 
0.0 -0.2763 0 -2.0 1e-06 
0.0 -0.2762 0 -2.0 1e-06 
0.0 -0.2761 0 -2.0 1e-06 
0.0 -0.276 0 -2.0 1e-06 
0.0 -0.2759 0 -2.0 1e-06 
0.0 -0.2758 0 -2.0 1e-06 
0.0 -0.2757 0 -2.0 1e-06 
0.0 -0.2756 0 -2.0 1e-06 
0.0 -0.2755 0 -2.0 1e-06 
0.0 -0.2754 0 -2.0 1e-06 
0.0 -0.2753 0 -2.0 1e-06 
0.0 -0.2752 0 -2.0 1e-06 
0.0 -0.2751 0 -2.0 1e-06 
0.0 -0.275 0 -2.0 1e-06 
0.0 -0.2749 0 -2.0 1e-06 
0.0 -0.2748 0 -2.0 1e-06 
0.0 -0.2747 0 -2.0 1e-06 
0.0 -0.2746 0 -2.0 1e-06 
0.0 -0.2745 0 -2.0 1e-06 
0.0 -0.2744 0 -2.0 1e-06 
0.0 -0.2743 0 -2.0 1e-06 
0.0 -0.2742 0 -2.0 1e-06 
0.0 -0.2741 0 -2.0 1e-06 
0.0 -0.274 0 -2.0 1e-06 
0.0 -0.2739 0 -2.0 1e-06 
0.0 -0.2738 0 -2.0 1e-06 
0.0 -0.2737 0 -2.0 1e-06 
0.0 -0.2736 0 -2.0 1e-06 
0.0 -0.2735 0 -2.0 1e-06 
0.0 -0.2734 0 -2.0 1e-06 
0.0 -0.2733 0 -2.0 1e-06 
0.0 -0.2732 0 -2.0 1e-06 
0.0 -0.2731 0 -2.0 1e-06 
0.0 -0.273 0 -2.0 1e-06 
0.0 -0.2729 0 -2.0 1e-06 
0.0 -0.2728 0 -2.0 1e-06 
0.0 -0.2727 0 -2.0 1e-06 
0.0 -0.2726 0 -2.0 1e-06 
0.0 -0.2725 0 -2.0 1e-06 
0.0 -0.2724 0 -2.0 1e-06 
0.0 -0.2723 0 -2.0 1e-06 
0.0 -0.2722 0 -2.0 1e-06 
0.0 -0.2721 0 -2.0 1e-06 
0.0 -0.272 0 -2.0 1e-06 
0.0 -0.2719 0 -2.0 1e-06 
0.0 -0.2718 0 -2.0 1e-06 
0.0 -0.2717 0 -2.0 1e-06 
0.0 -0.2716 0 -2.0 1e-06 
0.0 -0.2715 0 -2.0 1e-06 
0.0 -0.2714 0 -2.0 1e-06 
0.0 -0.2713 0 -2.0 1e-06 
0.0 -0.2712 0 -2.0 1e-06 
0.0 -0.2711 0 -2.0 1e-06 
0.0 -0.271 0 -2.0 1e-06 
0.0 -0.2709 0 -2.0 1e-06 
0.0 -0.2708 0 -2.0 1e-06 
0.0 -0.2707 0 -2.0 1e-06 
0.0 -0.2706 0 -2.0 1e-06 
0.0 -0.2705 0 -2.0 1e-06 
0.0 -0.2704 0 -2.0 1e-06 
0.0 -0.2703 0 -2.0 1e-06 
0.0 -0.2702 0 -2.0 1e-06 
0.0 -0.2701 0 -2.0 1e-06 
0.0 -0.27 0 -2.0 1e-06 
0.0 -0.2699 0 -2.0 1e-06 
0.0 -0.2698 0 -2.0 1e-06 
0.0 -0.2697 0 -2.0 1e-06 
0.0 -0.2696 0 -2.0 1e-06 
0.0 -0.2695 0 -2.0 1e-06 
0.0 -0.2694 0 -2.0 1e-06 
0.0 -0.2693 0 -2.0 1e-06 
0.0 -0.2692 0 -2.0 1e-06 
0.0 -0.2691 0 -2.0 1e-06 
0.0 -0.269 0 -2.0 1e-06 
0.0 -0.2689 0 -2.0 1e-06 
0.0 -0.2688 0 -2.0 1e-06 
0.0 -0.2687 0 -2.0 1e-06 
0.0 -0.2686 0 -2.0 1e-06 
0.0 -0.2685 0 -2.0 1e-06 
0.0 -0.2684 0 -2.0 1e-06 
0.0 -0.2683 0 -2.0 1e-06 
0.0 -0.2682 0 -2.0 1e-06 
0.0 -0.2681 0 -2.0 1e-06 
0.0 -0.268 0 -2.0 1e-06 
0.0 -0.2679 0 -2.0 1e-06 
0.0 -0.2678 0 -2.0 1e-06 
0.0 -0.2677 0 -2.0 1e-06 
0.0 -0.2676 0 -2.0 1e-06 
0.0 -0.2675 0 -2.0 1e-06 
0.0 -0.2674 0 -2.0 1e-06 
0.0 -0.2673 0 -2.0 1e-06 
0.0 -0.2672 0 -2.0 1e-06 
0.0 -0.2671 0 -2.0 1e-06 
0.0 -0.267 0 -2.0 1e-06 
0.0 -0.2669 0 -2.0 1e-06 
0.0 -0.2668 0 -2.0 1e-06 
0.0 -0.2667 0 -2.0 1e-06 
0.0 -0.2666 0 -2.0 1e-06 
0.0 -0.2665 0 -2.0 1e-06 
0.0 -0.2664 0 -2.0 1e-06 
0.0 -0.2663 0 -2.0 1e-06 
0.0 -0.2662 0 -2.0 1e-06 
0.0 -0.2661 0 -2.0 1e-06 
0.0 -0.266 0 -2.0 1e-06 
0.0 -0.2659 0 -2.0 1e-06 
0.0 -0.2658 0 -2.0 1e-06 
0.0 -0.2657 0 -2.0 1e-06 
0.0 -0.2656 0 -2.0 1e-06 
0.0 -0.2655 0 -2.0 1e-06 
0.0 -0.2654 0 -2.0 1e-06 
0.0 -0.2653 0 -2.0 1e-06 
0.0 -0.2652 0 -2.0 1e-06 
0.0 -0.2651 0 -2.0 1e-06 
0.0 -0.265 0 -2.0 1e-06 
0.0 -0.2649 0 -2.0 1e-06 
0.0 -0.2648 0 -2.0 1e-06 
0.0 -0.2647 0 -2.0 1e-06 
0.0 -0.2646 0 -2.0 1e-06 
0.0 -0.2645 0 -2.0 1e-06 
0.0 -0.2644 0 -2.0 1e-06 
0.0 -0.2643 0 -2.0 1e-06 
0.0 -0.2642 0 -2.0 1e-06 
0.0 -0.2641 0 -2.0 1e-06 
0.0 -0.264 0 -2.0 1e-06 
0.0 -0.2639 0 -2.0 1e-06 
0.0 -0.2638 0 -2.0 1e-06 
0.0 -0.2637 0 -2.0 1e-06 
0.0 -0.2636 0 -2.0 1e-06 
0.0 -0.2635 0 -2.0 1e-06 
0.0 -0.2634 0 -2.0 1e-06 
0.0 -0.2633 0 -2.0 1e-06 
0.0 -0.2632 0 -2.0 1e-06 
0.0 -0.2631 0 -2.0 1e-06 
0.0 -0.263 0 -2.0 1e-06 
0.0 -0.2629 0 -2.0 1e-06 
0.0 -0.2628 0 -2.0 1e-06 
0.0 -0.2627 0 -2.0 1e-06 
0.0 -0.2626 0 -2.0 1e-06 
0.0 -0.2625 0 -2.0 1e-06 
0.0 -0.2624 0 -2.0 1e-06 
0.0 -0.2623 0 -2.0 1e-06 
0.0 -0.2622 0 -2.0 1e-06 
0.0 -0.2621 0 -2.0 1e-06 
0.0 -0.262 0 -2.0 1e-06 
0.0 -0.2619 0 -2.0 1e-06 
0.0 -0.2618 0 -2.0 1e-06 
0.0 -0.2617 0 -2.0 1e-06 
0.0 -0.2616 0 -2.0 1e-06 
0.0 -0.2615 0 -2.0 1e-06 
0.0 -0.2614 0 -2.0 1e-06 
0.0 -0.2613 0 -2.0 1e-06 
0.0 -0.2612 0 -2.0 1e-06 
0.0 -0.2611 0 -2.0 1e-06 
0.0 -0.261 0 -2.0 1e-06 
0.0 -0.2609 0 -2.0 1e-06 
0.0 -0.2608 0 -2.0 1e-06 
0.0 -0.2607 0 -2.0 1e-06 
0.0 -0.2606 0 -2.0 1e-06 
0.0 -0.2605 0 -2.0 1e-06 
0.0 -0.2604 0 -2.0 1e-06 
0.0 -0.2603 0 -2.0 1e-06 
0.0 -0.2602 0 -2.0 1e-06 
0.0 -0.2601 0 -2.0 1e-06 
0.0 -0.26 0 -2.0 1e-06 
0.0 -0.2599 0 -2.0 1e-06 
0.0 -0.2598 0 -2.0 1e-06 
0.0 -0.2597 0 -2.0 1e-06 
0.0 -0.2596 0 -2.0 1e-06 
0.0 -0.2595 0 -2.0 1e-06 
0.0 -0.2594 0 -2.0 1e-06 
0.0 -0.2593 0 -2.0 1e-06 
0.0 -0.2592 0 -2.0 1e-06 
0.0 -0.2591 0 -2.0 1e-06 
0.0 -0.259 0 -2.0 1e-06 
0.0 -0.2589 0 -2.0 1e-06 
0.0 -0.2588 0 -2.0 1e-06 
0.0 -0.2587 0 -2.0 1e-06 
0.0 -0.2586 0 -2.0 1e-06 
0.0 -0.2585 0 -2.0 1e-06 
0.0 -0.2584 0 -2.0 1e-06 
0.0 -0.2583 0 -2.0 1e-06 
0.0 -0.2582 0 -2.0 1e-06 
0.0 -0.2581 0 -2.0 1e-06 
0.0 -0.258 0 -2.0 1e-06 
0.0 -0.2579 0 -2.0 1e-06 
0.0 -0.2578 0 -2.0 1e-06 
0.0 -0.2577 0 -2.0 1e-06 
0.0 -0.2576 0 -2.0 1e-06 
0.0 -0.2575 0 -2.0 1e-06 
0.0 -0.2574 0 -2.0 1e-06 
0.0 -0.2573 0 -2.0 1e-06 
0.0 -0.2572 0 -2.0 1e-06 
0.0 -0.2571 0 -2.0 1e-06 
0.0 -0.257 0 -2.0 1e-06 
0.0 -0.2569 0 -2.0 1e-06 
0.0 -0.2568 0 -2.0 1e-06 
0.0 -0.2567 0 -2.0 1e-06 
0.0 -0.2566 0 -2.0 1e-06 
0.0 -0.2565 0 -2.0 1e-06 
0.0 -0.2564 0 -2.0 1e-06 
0.0 -0.2563 0 -2.0 1e-06 
0.0 -0.2562 0 -2.0 1e-06 
0.0 -0.2561 0 -2.0 1e-06 
0.0 -0.256 0 -2.0 1e-06 
0.0 -0.2559 0 -2.0 1e-06 
0.0 -0.2558 0 -2.0 1e-06 
0.0 -0.2557 0 -2.0 1e-06 
0.0 -0.2556 0 -2.0 1e-06 
0.0 -0.2555 0 -2.0 1e-06 
0.0 -0.2554 0 -2.0 1e-06 
0.0 -0.2553 0 -2.0 1e-06 
0.0 -0.2552 0 -2.0 1e-06 
0.0 -0.2551 0 -2.0 1e-06 
0.0 -0.255 0 -2.0 1e-06 
0.0 -0.2549 0 -2.0 1e-06 
0.0 -0.2548 0 -2.0 1e-06 
0.0 -0.2547 0 -2.0 1e-06 
0.0 -0.2546 0 -2.0 1e-06 
0.0 -0.2545 0 -2.0 1e-06 
0.0 -0.2544 0 -2.0 1e-06 
0.0 -0.2543 0 -2.0 1e-06 
0.0 -0.2542 0 -2.0 1e-06 
0.0 -0.2541 0 -2.0 1e-06 
0.0 -0.254 0 -2.0 1e-06 
0.0 -0.2539 0 -2.0 1e-06 
0.0 -0.2538 0 -2.0 1e-06 
0.0 -0.2537 0 -2.0 1e-06 
0.0 -0.2536 0 -2.0 1e-06 
0.0 -0.2535 0 -2.0 1e-06 
0.0 -0.2534 0 -2.0 1e-06 
0.0 -0.2533 0 -2.0 1e-06 
0.0 -0.2532 0 -2.0 1e-06 
0.0 -0.2531 0 -2.0 1e-06 
0.0 -0.253 0 -2.0 1e-06 
0.0 -0.2529 0 -2.0 1e-06 
0.0 -0.2528 0 -2.0 1e-06 
0.0 -0.2527 0 -2.0 1e-06 
0.0 -0.2526 0 -2.0 1e-06 
0.0 -0.2525 0 -2.0 1e-06 
0.0 -0.2524 0 -2.0 1e-06 
0.0 -0.2523 0 -2.0 1e-06 
0.0 -0.2522 0 -2.0 1e-06 
0.0 -0.2521 0 -2.0 1e-06 
0.0 -0.252 0 -2.0 1e-06 
0.0 -0.2519 0 -2.0 1e-06 
0.0 -0.2518 0 -2.0 1e-06 
0.0 -0.2517 0 -2.0 1e-06 
0.0 -0.2516 0 -2.0 1e-06 
0.0 -0.2515 0 -2.0 1e-06 
0.0 -0.2514 0 -2.0 1e-06 
0.0 -0.2513 0 -2.0 1e-06 
0.0 -0.2512 0 -2.0 1e-06 
0.0 -0.2511 0 -2.0 1e-06 
0.0 -0.251 0 -2.0 1e-06 
0.0 -0.2509 0 -2.0 1e-06 
0.0 -0.2508 0 -2.0 1e-06 
0.0 -0.2507 0 -2.0 1e-06 
0.0 -0.2506 0 -2.0 1e-06 
0.0 -0.2505 0 -2.0 1e-06 
0.0 -0.2504 0 -2.0 1e-06 
0.0 -0.2503 0 -2.0 1e-06 
0.0 -0.2502 0 -2.0 1e-06 
0.0 -0.2501 0 -2.0 1e-06 
0.0 -0.25 0 -2.0 1e-06 
0.0 -0.2499 0 -2.0 1e-06 
0.0 -0.2498 0 -2.0 1e-06 
0.0 -0.2497 0 -2.0 1e-06 
0.0 -0.2496 0 -2.0 1e-06 
0.0 -0.2495 0 -2.0 1e-06 
0.0 -0.2494 0 -2.0 1e-06 
0.0 -0.2493 0 -2.0 1e-06 
0.0 -0.2492 0 -2.0 1e-06 
0.0 -0.2491 0 -2.0 1e-06 
0.0 -0.249 0 -2.0 1e-06 
0.0 -0.2489 0 -2.0 1e-06 
0.0 -0.2488 0 -2.0 1e-06 
0.0 -0.2487 0 -2.0 1e-06 
0.0 -0.2486 0 -2.0 1e-06 
0.0 -0.2485 0 -2.0 1e-06 
0.0 -0.2484 0 -2.0 1e-06 
0.0 -0.2483 0 -2.0 1e-06 
0.0 -0.2482 0 -2.0 1e-06 
0.0 -0.2481 0 -2.0 1e-06 
0.0 -0.248 0 -2.0 1e-06 
0.0 -0.2479 0 -2.0 1e-06 
0.0 -0.2478 0 -2.0 1e-06 
0.0 -0.2477 0 -2.0 1e-06 
0.0 -0.2476 0 -2.0 1e-06 
0.0 -0.2475 0 -2.0 1e-06 
0.0 -0.2474 0 -2.0 1e-06 
0.0 -0.2473 0 -2.0 1e-06 
0.0 -0.2472 0 -2.0 1e-06 
0.0 -0.2471 0 -2.0 1e-06 
0.0 -0.247 0 -2.0 1e-06 
0.0 -0.2469 0 -2.0 1e-06 
0.0 -0.2468 0 -2.0 1e-06 
0.0 -0.2467 0 -2.0 1e-06 
0.0 -0.2466 0 -2.0 1e-06 
0.0 -0.2465 0 -2.0 1e-06 
0.0 -0.2464 0 -2.0 1e-06 
0.0 -0.2463 0 -2.0 1e-06 
0.0 -0.2462 0 -2.0 1e-06 
0.0 -0.2461 0 -2.0 1e-06 
0.0 -0.246 0 -2.0 1e-06 
0.0 -0.2459 0 -2.0 1e-06 
0.0 -0.2458 0 -2.0 1e-06 
0.0 -0.2457 0 -2.0 1e-06 
0.0 -0.2456 0 -2.0 1e-06 
0.0 -0.2455 0 -2.0 1e-06 
0.0 -0.2454 0 -2.0 1e-06 
0.0 -0.2453 0 -2.0 1e-06 
0.0 -0.2452 0 -2.0 1e-06 
0.0 -0.2451 0 -2.0 1e-06 
0.0 -0.245 0 -2.0 1e-06 
0.0 -0.2449 0 -2.0 1e-06 
0.0 -0.2448 0 -2.0 1e-06 
0.0 -0.2447 0 -2.0 1e-06 
0.0 -0.2446 0 -2.0 1e-06 
0.0 -0.2445 0 -2.0 1e-06 
0.0 -0.2444 0 -2.0 1e-06 
0.0 -0.2443 0 -2.0 1e-06 
0.0 -0.2442 0 -2.0 1e-06 
0.0 -0.2441 0 -2.0 1e-06 
0.0 -0.244 0 -2.0 1e-06 
0.0 -0.2439 0 -2.0 1e-06 
0.0 -0.2438 0 -2.0 1e-06 
0.0 -0.2437 0 -2.0 1e-06 
0.0 -0.2436 0 -2.0 1e-06 
0.0 -0.2435 0 -2.0 1e-06 
0.0 -0.2434 0 -2.0 1e-06 
0.0 -0.2433 0 -2.0 1e-06 
0.0 -0.2432 0 -2.0 1e-06 
0.0 -0.2431 0 -2.0 1e-06 
0.0 -0.243 0 -2.0 1e-06 
0.0 -0.2429 0 -2.0 1e-06 
0.0 -0.2428 0 -2.0 1e-06 
0.0 -0.2427 0 -2.0 1e-06 
0.0 -0.2426 0 -2.0 1e-06 
0.0 -0.2425 0 -2.0 1e-06 
0.0 -0.2424 0 -2.0 1e-06 
0.0 -0.2423 0 -2.0 1e-06 
0.0 -0.2422 0 -2.0 1e-06 
0.0 -0.2421 0 -2.0 1e-06 
0.0 -0.242 0 -2.0 1e-06 
0.0 -0.2419 0 -2.0 1e-06 
0.0 -0.2418 0 -2.0 1e-06 
0.0 -0.2417 0 -2.0 1e-06 
0.0 -0.2416 0 -2.0 1e-06 
0.0 -0.2415 0 -2.0 1e-06 
0.0 -0.2414 0 -2.0 1e-06 
0.0 -0.2413 0 -2.0 1e-06 
0.0 -0.2412 0 -2.0 1e-06 
0.0 -0.2411 0 -2.0 1e-06 
0.0 -0.241 0 -2.0 1e-06 
0.0 -0.2409 0 -2.0 1e-06 
0.0 -0.2408 0 -2.0 1e-06 
0.0 -0.2407 0 -2.0 1e-06 
0.0 -0.2406 0 -2.0 1e-06 
0.0 -0.2405 0 -2.0 1e-06 
0.0 -0.2404 0 -2.0 1e-06 
0.0 -0.2403 0 -2.0 1e-06 
0.0 -0.2402 0 -2.0 1e-06 
0.0 -0.2401 0 -2.0 1e-06 
0.0 -0.24 0 -2.0 1e-06 
0.0 -0.2399 0 -2.0 1e-06 
0.0 -0.2398 0 -2.0 1e-06 
0.0 -0.2397 0 -2.0 1e-06 
0.0 -0.2396 0 -2.0 1e-06 
0.0 -0.2395 0 -2.0 1e-06 
0.0 -0.2394 0 -2.0 1e-06 
0.0 -0.2393 0 -2.0 1e-06 
0.0 -0.2392 0 -2.0 1e-06 
0.0 -0.2391 0 -2.0 1e-06 
0.0 -0.239 0 -2.0 1e-06 
0.0 -0.2389 0 -2.0 1e-06 
0.0 -0.2388 0 -2.0 1e-06 
0.0 -0.2387 0 -2.0 1e-06 
0.0 -0.2386 0 -2.0 1e-06 
0.0 -0.2385 0 -2.0 1e-06 
0.0 -0.2384 0 -2.0 1e-06 
0.0 -0.2383 0 -2.0 1e-06 
0.0 -0.2382 0 -2.0 1e-06 
0.0 -0.2381 0 -2.0 1e-06 
0.0 -0.238 0 -2.0 1e-06 
0.0 -0.2379 0 -2.0 1e-06 
0.0 -0.2378 0 -2.0 1e-06 
0.0 -0.2377 0 -2.0 1e-06 
0.0 -0.2376 0 -2.0 1e-06 
0.0 -0.2375 0 -2.0 1e-06 
0.0 -0.2374 0 -2.0 1e-06 
0.0 -0.2373 0 -2.0 1e-06 
0.0 -0.2372 0 -2.0 1e-06 
0.0 -0.2371 0 -2.0 1e-06 
0.0 -0.237 0 -2.0 1e-06 
0.0 -0.2369 0 -2.0 1e-06 
0.0 -0.2368 0 -2.0 1e-06 
0.0 -0.2367 0 -2.0 1e-06 
0.0 -0.2366 0 -2.0 1e-06 
0.0 -0.2365 0 -2.0 1e-06 
0.0 -0.2364 0 -2.0 1e-06 
0.0 -0.2363 0 -2.0 1e-06 
0.0 -0.2362 0 -2.0 1e-06 
0.0 -0.2361 0 -2.0 1e-06 
0.0 -0.236 0 -2.0 1e-06 
0.0 -0.2359 0 -2.0 1e-06 
0.0 -0.2358 0 -2.0 1e-06 
0.0 -0.2357 0 -2.0 1e-06 
0.0 -0.2356 0 -2.0 1e-06 
0.0 -0.2355 0 -2.0 1e-06 
0.0 -0.2354 0 -2.0 1e-06 
0.0 -0.2353 0 -2.0 1e-06 
0.0 -0.2352 0 -2.0 1e-06 
0.0 -0.2351 0 -2.0 1e-06 
0.0 -0.235 0 -2.0 1e-06 
0.0 -0.2349 0 -2.0 1e-06 
0.0 -0.2348 0 -2.0 1e-06 
0.0 -0.2347 0 -2.0 1e-06 
0.0 -0.2346 0 -2.0 1e-06 
0.0 -0.2345 0 -2.0 1e-06 
0.0 -0.2344 0 -2.0 1e-06 
0.0 -0.2343 0 -2.0 1e-06 
0.0 -0.2342 0 -2.0 1e-06 
0.0 -0.2341 0 -2.0 1e-06 
0.0 -0.234 0 -2.0 1e-06 
0.0 -0.2339 0 -2.0 1e-06 
0.0 -0.2338 0 -2.0 1e-06 
0.0 -0.2337 0 -2.0 1e-06 
0.0 -0.2336 0 -2.0 1e-06 
0.0 -0.2335 0 -2.0 1e-06 
0.0 -0.2334 0 -2.0 1e-06 
0.0 -0.2333 0 -2.0 1e-06 
0.0 -0.2332 0 -2.0 1e-06 
0.0 -0.2331 0 -2.0 1e-06 
0.0 -0.233 0 -2.0 1e-06 
0.0 -0.2329 0 -2.0 1e-06 
0.0 -0.2328 0 -2.0 1e-06 
0.0 -0.2327 0 -2.0 1e-06 
0.0 -0.2326 0 -2.0 1e-06 
0.0 -0.2325 0 -2.0 1e-06 
0.0 -0.2324 0 -2.0 1e-06 
0.0 -0.2323 0 -2.0 1e-06 
0.0 -0.2322 0 -2.0 1e-06 
0.0 -0.2321 0 -2.0 1e-06 
0.0 -0.232 0 -2.0 1e-06 
0.0 -0.2319 0 -2.0 1e-06 
0.0 -0.2318 0 -2.0 1e-06 
0.0 -0.2317 0 -2.0 1e-06 
0.0 -0.2316 0 -2.0 1e-06 
0.0 -0.2315 0 -2.0 1e-06 
0.0 -0.2314 0 -2.0 1e-06 
0.0 -0.2313 0 -2.0 1e-06 
0.0 -0.2312 0 -2.0 1e-06 
0.0 -0.2311 0 -2.0 1e-06 
0.0 -0.231 0 -2.0 1e-06 
0.0 -0.2309 0 -2.0 1e-06 
0.0 -0.2308 0 -2.0 1e-06 
0.0 -0.2307 0 -2.0 1e-06 
0.0 -0.2306 0 -2.0 1e-06 
0.0 -0.2305 0 -2.0 1e-06 
0.0 -0.2304 0 -2.0 1e-06 
0.0 -0.2303 0 -2.0 1e-06 
0.0 -0.2302 0 -2.0 1e-06 
0.0 -0.2301 0 -2.0 1e-06 
0.0 -0.23 0 -2.0 1e-06 
0.0 -0.2299 0 -2.0 1e-06 
0.0 -0.2298 0 -2.0 1e-06 
0.0 -0.2297 0 -2.0 1e-06 
0.0 -0.2296 0 -2.0 1e-06 
0.0 -0.2295 0 -2.0 1e-06 
0.0 -0.2294 0 -2.0 1e-06 
0.0 -0.2293 0 -2.0 1e-06 
0.0 -0.2292 0 -2.0 1e-06 
0.0 -0.2291 0 -2.0 1e-06 
0.0 -0.229 0 -2.0 1e-06 
0.0 -0.2289 0 -2.0 1e-06 
0.0 -0.2288 0 -2.0 1e-06 
0.0 -0.2287 0 -2.0 1e-06 
0.0 -0.2286 0 -2.0 1e-06 
0.0 -0.2285 0 -2.0 1e-06 
0.0 -0.2284 0 -2.0 1e-06 
0.0 -0.2283 0 -2.0 1e-06 
0.0 -0.2282 0 -2.0 1e-06 
0.0 -0.2281 0 -2.0 1e-06 
0.0 -0.228 0 -2.0 1e-06 
0.0 -0.2279 0 -2.0 1e-06 
0.0 -0.2278 0 -2.0 1e-06 
0.0 -0.2277 0 -2.0 1e-06 
0.0 -0.2276 0 -2.0 1e-06 
0.0 -0.2275 0 -2.0 1e-06 
0.0 -0.2274 0 -2.0 1e-06 
0.0 -0.2273 0 -2.0 1e-06 
0.0 -0.2272 0 -2.0 1e-06 
0.0 -0.2271 0 -2.0 1e-06 
0.0 -0.227 0 -2.0 1e-06 
0.0 -0.2269 0 -2.0 1e-06 
0.0 -0.2268 0 -2.0 1e-06 
0.0 -0.2267 0 -2.0 1e-06 
0.0 -0.2266 0 -2.0 1e-06 
0.0 -0.2265 0 -2.0 1e-06 
0.0 -0.2264 0 -2.0 1e-06 
0.0 -0.2263 0 -2.0 1e-06 
0.0 -0.2262 0 -2.0 1e-06 
0.0 -0.2261 0 -2.0 1e-06 
0.0 -0.226 0 -2.0 1e-06 
0.0 -0.2259 0 -2.0 1e-06 
0.0 -0.2258 0 -2.0 1e-06 
0.0 -0.2257 0 -2.0 1e-06 
0.0 -0.2256 0 -2.0 1e-06 
0.0 -0.2255 0 -2.0 1e-06 
0.0 -0.2254 0 -2.0 1e-06 
0.0 -0.2253 0 -2.0 1e-06 
0.0 -0.2252 0 -2.0 1e-06 
0.0 -0.2251 0 -2.0 1e-06 
0.0 -0.225 0 -2.0 1e-06 
0.0 -0.2249 0 -2.0 1e-06 
0.0 -0.2248 0 -2.0 1e-06 
0.0 -0.2247 0 -2.0 1e-06 
0.0 -0.2246 0 -2.0 1e-06 
0.0 -0.2245 0 -2.0 1e-06 
0.0 -0.2244 0 -2.0 1e-06 
0.0 -0.2243 0 -2.0 1e-06 
0.0 -0.2242 0 -2.0 1e-06 
0.0 -0.2241 0 -2.0 1e-06 
0.0 -0.224 0 -2.0 1e-06 
0.0 -0.2239 0 -2.0 1e-06 
0.0 -0.2238 0 -2.0 1e-06 
0.0 -0.2237 0 -2.0 1e-06 
0.0 -0.2236 0 -2.0 1e-06 
0.0 -0.2235 0 -2.0 1e-06 
0.0 -0.2234 0 -2.0 1e-06 
0.0 -0.2233 0 -2.0 1e-06 
0.0 -0.2232 0 -2.0 1e-06 
0.0 -0.2231 0 -2.0 1e-06 
0.0 -0.223 0 -2.0 1e-06 
0.0 -0.2229 0 -2.0 1e-06 
0.0 -0.2228 0 -2.0 1e-06 
0.0 -0.2227 0 -2.0 1e-06 
0.0 -0.2226 0 -2.0 1e-06 
0.0 -0.2225 0 -2.0 1e-06 
0.0 -0.2224 0 -2.0 1e-06 
0.0 -0.2223 0 -2.0 1e-06 
0.0 -0.2222 0 -2.0 1e-06 
0.0 -0.2221 0 -2.0 1e-06 
0.0 -0.222 0 -2.0 1e-06 
0.0 -0.2219 0 -2.0 1e-06 
0.0 -0.2218 0 -2.0 1e-06 
0.0 -0.2217 0 -2.0 1e-06 
0.0 -0.2216 0 -2.0 1e-06 
0.0 -0.2215 0 -2.0 1e-06 
0.0 -0.2214 0 -2.0 1e-06 
0.0 -0.2213 0 -2.0 1e-06 
0.0 -0.2212 0 -2.0 1e-06 
0.0 -0.2211 0 -2.0 1e-06 
0.0 -0.221 0 -2.0 1e-06 
0.0 -0.2209 0 -2.0 1e-06 
0.0 -0.2208 0 -2.0 1e-06 
0.0 -0.2207 0 -2.0 1e-06 
0.0 -0.2206 0 -2.0 1e-06 
0.0 -0.2205 0 -2.0 1e-06 
0.0 -0.2204 0 -2.0 1e-06 
0.0 -0.2203 0 -2.0 1e-06 
0.0 -0.2202 0 -2.0 1e-06 
0.0 -0.2201 0 -2.0 1e-06 
0.0 -0.22 0 -2.0 1e-06 
0.0 -0.2199 0 -2.0 1e-06 
0.0 -0.2198 0 -2.0 1e-06 
0.0 -0.2197 0 -2.0 1e-06 
0.0 -0.2196 0 -2.0 1e-06 
0.0 -0.2195 0 -2.0 1e-06 
0.0 -0.2194 0 -2.0 1e-06 
0.0 -0.2193 0 -2.0 1e-06 
0.0 -0.2192 0 -2.0 1e-06 
0.0 -0.2191 0 -2.0 1e-06 
0.0 -0.219 0 -2.0 1e-06 
0.0 -0.2189 0 -2.0 1e-06 
0.0 -0.2188 0 -2.0 1e-06 
0.0 -0.2187 0 -2.0 1e-06 
0.0 -0.2186 0 -2.0 1e-06 
0.0 -0.2185 0 -2.0 1e-06 
0.0 -0.2184 0 -2.0 1e-06 
0.0 -0.2183 0 -2.0 1e-06 
0.0 -0.2182 0 -2.0 1e-06 
0.0 -0.2181 0 -2.0 1e-06 
0.0 -0.218 0 -2.0 1e-06 
0.0 -0.2179 0 -2.0 1e-06 
0.0 -0.2178 0 -2.0 1e-06 
0.0 -0.2177 0 -2.0 1e-06 
0.0 -0.2176 0 -2.0 1e-06 
0.0 -0.2175 0 -2.0 1e-06 
0.0 -0.2174 0 -2.0 1e-06 
0.0 -0.2173 0 -2.0 1e-06 
0.0 -0.2172 0 -2.0 1e-06 
0.0 -0.2171 0 -2.0 1e-06 
0.0 -0.217 0 -2.0 1e-06 
0.0 -0.2169 0 -2.0 1e-06 
0.0 -0.2168 0 -2.0 1e-06 
0.0 -0.2167 0 -2.0 1e-06 
0.0 -0.2166 0 -2.0 1e-06 
0.0 -0.2165 0 -2.0 1e-06 
0.0 -0.2164 0 -2.0 1e-06 
0.0 -0.2163 0 -2.0 1e-06 
0.0 -0.2162 0 -2.0 1e-06 
0.0 -0.2161 0 -2.0 1e-06 
0.0 -0.216 0 -2.0 1e-06 
0.0 -0.2159 0 -2.0 1e-06 
0.0 -0.2158 0 -2.0 1e-06 
0.0 -0.2157 0 -2.0 1e-06 
0.0 -0.2156 0 -2.0 1e-06 
0.0 -0.2155 0 -2.0 1e-06 
0.0 -0.2154 0 -2.0 1e-06 
0.0 -0.2153 0 -2.0 1e-06 
0.0 -0.2152 0 -2.0 1e-06 
0.0 -0.2151 0 -2.0 1e-06 
0.0 -0.215 0 -2.0 1e-06 
0.0 -0.2149 0 -2.0 1e-06 
0.0 -0.2148 0 -2.0 1e-06 
0.0 -0.2147 0 -2.0 1e-06 
0.0 -0.2146 0 -2.0 1e-06 
0.0 -0.2145 0 -2.0 1e-06 
0.0 -0.2144 0 -2.0 1e-06 
0.0 -0.2143 0 -2.0 1e-06 
0.0 -0.2142 0 -2.0 1e-06 
0.0 -0.2141 0 -2.0 1e-06 
0.0 -0.214 0 -2.0 1e-06 
0.0 -0.2139 0 -2.0 1e-06 
0.0 -0.2138 0 -2.0 1e-06 
0.0 -0.2137 0 -2.0 1e-06 
0.0 -0.2136 0 -2.0 1e-06 
0.0 -0.2135 0 -2.0 1e-06 
0.0 -0.2134 0 -2.0 1e-06 
0.0 -0.2133 0 -2.0 1e-06 
0.0 -0.2132 0 -2.0 1e-06 
0.0 -0.2131 0 -2.0 1e-06 
0.0 -0.213 0 -2.0 1e-06 
0.0 -0.2129 0 -2.0 1e-06 
0.0 -0.2128 0 -2.0 1e-06 
0.0 -0.2127 0 -2.0 1e-06 
0.0 -0.2126 0 -2.0 1e-06 
0.0 -0.2125 0 -2.0 1e-06 
0.0 -0.2124 0 -2.0 1e-06 
0.0 -0.2123 0 -2.0 1e-06 
0.0 -0.2122 0 -2.0 1e-06 
0.0 -0.2121 0 -2.0 1e-06 
0.0 -0.212 0 -2.0 1e-06 
0.0 -0.2119 0 -2.0 1e-06 
0.0 -0.2118 0 -2.0 1e-06 
0.0 -0.2117 0 -2.0 1e-06 
0.0 -0.2116 0 -2.0 1e-06 
0.0 -0.2115 0 -2.0 1e-06 
0.0 -0.2114 0 -2.0 1e-06 
0.0 -0.2113 0 -2.0 1e-06 
0.0 -0.2112 0 -2.0 1e-06 
0.0 -0.2111 0 -2.0 1e-06 
0.0 -0.211 0 -2.0 1e-06 
0.0 -0.2109 0 -2.0 1e-06 
0.0 -0.2108 0 -2.0 1e-06 
0.0 -0.2107 0 -2.0 1e-06 
0.0 -0.2106 0 -2.0 1e-06 
0.0 -0.2105 0 -2.0 1e-06 
0.0 -0.2104 0 -2.0 1e-06 
0.0 -0.2103 0 -2.0 1e-06 
0.0 -0.2102 0 -2.0 1e-06 
0.0 -0.2101 0 -2.0 1e-06 
0.0 -0.21 0 -2.0 1e-06 
0.0 -0.2099 0 -2.0 1e-06 
0.0 -0.2098 0 -2.0 1e-06 
0.0 -0.2097 0 -2.0 1e-06 
0.0 -0.2096 0 -2.0 1e-06 
0.0 -0.2095 0 -2.0 1e-06 
0.0 -0.2094 0 -2.0 1e-06 
0.0 -0.2093 0 -2.0 1e-06 
0.0 -0.2092 0 -2.0 1e-06 
0.0 -0.2091 0 -2.0 1e-06 
0.0 -0.209 0 -2.0 1e-06 
0.0 -0.2089 0 -2.0 1e-06 
0.0 -0.2088 0 -2.0 1e-06 
0.0 -0.2087 0 -2.0 1e-06 
0.0 -0.2086 0 -2.0 1e-06 
0.0 -0.2085 0 -2.0 1e-06 
0.0 -0.2084 0 -2.0 1e-06 
0.0 -0.2083 0 -2.0 1e-06 
0.0 -0.2082 0 -2.0 1e-06 
0.0 -0.2081 0 -2.0 1e-06 
0.0 -0.208 0 -2.0 1e-06 
0.0 -0.2079 0 -2.0 1e-06 
0.0 -0.2078 0 -2.0 1e-06 
0.0 -0.2077 0 -2.0 1e-06 
0.0 -0.2076 0 -2.0 1e-06 
0.0 -0.2075 0 -2.0 1e-06 
0.0 -0.2074 0 -2.0 1e-06 
0.0 -0.2073 0 -2.0 1e-06 
0.0 -0.2072 0 -2.0 1e-06 
0.0 -0.2071 0 -2.0 1e-06 
0.0 -0.207 0 -2.0 1e-06 
0.0 -0.2069 0 -2.0 1e-06 
0.0 -0.2068 0 -2.0 1e-06 
0.0 -0.2067 0 -2.0 1e-06 
0.0 -0.2066 0 -2.0 1e-06 
0.0 -0.2065 0 -2.0 1e-06 
0.0 -0.2064 0 -2.0 1e-06 
0.0 -0.2063 0 -2.0 1e-06 
0.0 -0.2062 0 -2.0 1e-06 
0.0 -0.2061 0 -2.0 1e-06 
0.0 -0.206 0 -2.0 1e-06 
0.0 -0.2059 0 -2.0 1e-06 
0.0 -0.2058 0 -2.0 1e-06 
0.0 -0.2057 0 -2.0 1e-06 
0.0 -0.2056 0 -2.0 1e-06 
0.0 -0.2055 0 -2.0 1e-06 
0.0 -0.2054 0 -2.0 1e-06 
0.0 -0.2053 0 -2.0 1e-06 
0.0 -0.2052 0 -2.0 1e-06 
0.0 -0.2051 0 -2.0 1e-06 
0.0 -0.205 0 -2.0 1e-06 
0.0 -0.2049 0 -2.0 1e-06 
0.0 -0.2048 0 -2.0 1e-06 
0.0 -0.2047 0 -2.0 1e-06 
0.0 -0.2046 0 -2.0 1e-06 
0.0 -0.2045 0 -2.0 1e-06 
0.0 -0.2044 0 -2.0 1e-06 
0.0 -0.2043 0 -2.0 1e-06 
0.0 -0.2042 0 -2.0 1e-06 
0.0 -0.2041 0 -2.0 1e-06 
0.0 -0.204 0 -2.0 1e-06 
0.0 -0.2039 0 -2.0 1e-06 
0.0 -0.2038 0 -2.0 1e-06 
0.0 -0.2037 0 -2.0 1e-06 
0.0 -0.2036 0 -2.0 1e-06 
0.0 -0.2035 0 -2.0 1e-06 
0.0 -0.2034 0 -2.0 1e-06 
0.0 -0.2033 0 -2.0 1e-06 
0.0 -0.2032 0 -2.0 1e-06 
0.0 -0.2031 0 -2.0 1e-06 
0.0 -0.203 0 -2.0 1e-06 
0.0 -0.2029 0 -2.0 1e-06 
0.0 -0.2028 0 -2.0 1e-06 
0.0 -0.2027 0 -2.0 1e-06 
0.0 -0.2026 0 -2.0 1e-06 
0.0 -0.2025 0 -2.0 1e-06 
0.0 -0.2024 0 -2.0 1e-06 
0.0 -0.2023 0 -2.0 1e-06 
0.0 -0.2022 0 -2.0 1e-06 
0.0 -0.2021 0 -2.0 1e-06 
0.0 -0.202 0 -2.0 1e-06 
0.0 -0.2019 0 -2.0 1e-06 
0.0 -0.2018 0 -2.0 1e-06 
0.0 -0.2017 0 -2.0 1e-06 
0.0 -0.2016 0 -2.0 1e-06 
0.0 -0.2015 0 -2.0 1e-06 
0.0 -0.2014 0 -2.0 1e-06 
0.0 -0.2013 0 -2.0 1e-06 
0.0 -0.2012 0 -2.0 1e-06 
0.0 -0.2011 0 -2.0 1e-06 
0.0 -0.201 0 -2.0 1e-06 
0.0 -0.2009 0 -2.0 1e-06 
0.0 -0.2008 0 -2.0 1e-06 
0.0 -0.2007 0 -2.0 1e-06 
0.0 -0.2006 0 -2.0 1e-06 
0.0 -0.2005 0 -2.0 1e-06 
0.0 -0.2004 0 -2.0 1e-06 
0.0 -0.2003 0 -2.0 1e-06 
0.0 -0.2002 0 -2.0 1e-06 
0.0 -0.2001 0 -2.0 1e-06 
0.0 -0.2 0 -2.0 1e-06 
0.0 -0.1999 0 -2.0 1e-06 
0.0 -0.1998 0 -2.0 1e-06 
0.0 -0.1997 0 -2.0 1e-06 
0.0 -0.1996 0 -2.0 1e-06 
0.0 -0.1995 0 -2.0 1e-06 
0.0 -0.1994 0 -2.0 1e-06 
0.0 -0.1993 0 -2.0 1e-06 
0.0 -0.1992 0 -2.0 1e-06 
0.0 -0.1991 0 -2.0 1e-06 
0.0 -0.199 0 -2.0 1e-06 
0.0 -0.1989 0 -2.0 1e-06 
0.0 -0.1988 0 -2.0 1e-06 
0.0 -0.1987 0 -2.0 1e-06 
0.0 -0.1986 0 -2.0 1e-06 
0.0 -0.1985 0 -2.0 1e-06 
0.0 -0.1984 0 -2.0 1e-06 
0.0 -0.1983 0 -2.0 1e-06 
0.0 -0.1982 0 -2.0 1e-06 
0.0 -0.1981 0 -2.0 1e-06 
0.0 -0.198 0 -2.0 1e-06 
0.0 -0.1979 0 -2.0 1e-06 
0.0 -0.1978 0 -2.0 1e-06 
0.0 -0.1977 0 -2.0 1e-06 
0.0 -0.1976 0 -2.0 1e-06 
0.0 -0.1975 0 -2.0 1e-06 
0.0 -0.1974 0 -2.0 1e-06 
0.0 -0.1973 0 -2.0 1e-06 
0.0 -0.1972 0 -2.0 1e-06 
0.0 -0.1971 0 -2.0 1e-06 
0.0 -0.197 0 -2.0 1e-06 
0.0 -0.1969 0 -2.0 1e-06 
0.0 -0.1968 0 -2.0 1e-06 
0.0 -0.1967 0 -2.0 1e-06 
0.0 -0.1966 0 -2.0 1e-06 
0.0 -0.1965 0 -2.0 1e-06 
0.0 -0.1964 0 -2.0 1e-06 
0.0 -0.1963 0 -2.0 1e-06 
0.0 -0.1962 0 -2.0 1e-06 
0.0 -0.1961 0 -2.0 1e-06 
0.0 -0.196 0 -2.0 1e-06 
0.0 -0.1959 0 -2.0 1e-06 
0.0 -0.1958 0 -2.0 1e-06 
0.0 -0.1957 0 -2.0 1e-06 
0.0 -0.1956 0 -2.0 1e-06 
0.0 -0.1955 0 -2.0 1e-06 
0.0 -0.1954 0 -2.0 1e-06 
0.0 -0.1953 0 -2.0 1e-06 
0.0 -0.1952 0 -2.0 1e-06 
0.0 -0.1951 0 -2.0 1e-06 
0.0 -0.195 0 -2.0 1e-06 
0.0 -0.1949 0 -2.0 1e-06 
0.0 -0.1948 0 -2.0 1e-06 
0.0 -0.1947 0 -2.0 1e-06 
0.0 -0.1946 0 -2.0 1e-06 
0.0 -0.1945 0 -2.0 1e-06 
0.0 -0.1944 0 -2.0 1e-06 
0.0 -0.1943 0 -2.0 1e-06 
0.0 -0.1942 0 -2.0 1e-06 
0.0 -0.1941 0 -2.0 1e-06 
0.0 -0.194 0 -2.0 1e-06 
0.0 -0.1939 0 -2.0 1e-06 
0.0 -0.1938 0 -2.0 1e-06 
0.0 -0.1937 0 -2.0 1e-06 
0.0 -0.1936 0 -2.0 1e-06 
0.0 -0.1935 0 -2.0 1e-06 
0.0 -0.1934 0 -2.0 1e-06 
0.0 -0.1933 0 -2.0 1e-06 
0.0 -0.1932 0 -2.0 1e-06 
0.0 -0.1931 0 -2.0 1e-06 
0.0 -0.193 0 -2.0 1e-06 
0.0 -0.1929 0 -2.0 1e-06 
0.0 -0.1928 0 -2.0 1e-06 
0.0 -0.1927 0 -2.0 1e-06 
0.0 -0.1926 0 -2.0 1e-06 
0.0 -0.1925 0 -2.0 1e-06 
0.0 -0.1924 0 -2.0 1e-06 
0.0 -0.1923 0 -2.0 1e-06 
0.0 -0.1922 0 -2.0 1e-06 
0.0 -0.1921 0 -2.0 1e-06 
0.0 -0.192 0 -2.0 1e-06 
0.0 -0.1919 0 -2.0 1e-06 
0.0 -0.1918 0 -2.0 1e-06 
0.0 -0.1917 0 -2.0 1e-06 
0.0 -0.1916 0 -2.0 1e-06 
0.0 -0.1915 0 -2.0 1e-06 
0.0 -0.1914 0 -2.0 1e-06 
0.0 -0.1913 0 -2.0 1e-06 
0.0 -0.1912 0 -2.0 1e-06 
0.0 -0.1911 0 -2.0 1e-06 
0.0 -0.191 0 -2.0 1e-06 
0.0 -0.1909 0 -2.0 1e-06 
0.0 -0.1908 0 -2.0 1e-06 
0.0 -0.1907 0 -2.0 1e-06 
0.0 -0.1906 0 -2.0 1e-06 
0.0 -0.1905 0 -2.0 1e-06 
0.0 -0.1904 0 -2.0 1e-06 
0.0 -0.1903 0 -2.0 1e-06 
0.0 -0.1902 0 -2.0 1e-06 
0.0 -0.1901 0 -2.0 1e-06 
0.0 -0.19 0 -2.0 1e-06 
0.0 -0.1899 0 -2.0 1e-06 
0.0 -0.1898 0 -2.0 1e-06 
0.0 -0.1897 0 -2.0 1e-06 
0.0 -0.1896 0 -2.0 1e-06 
0.0 -0.1895 0 -2.0 1e-06 
0.0 -0.1894 0 -2.0 1e-06 
0.0 -0.1893 0 -2.0 1e-06 
0.0 -0.1892 0 -2.0 1e-06 
0.0 -0.1891 0 -2.0 1e-06 
0.0 -0.189 0 -2.0 1e-06 
0.0 -0.1889 0 -2.0 1e-06 
0.0 -0.1888 0 -2.0 1e-06 
0.0 -0.1887 0 -2.0 1e-06 
0.0 -0.1886 0 -2.0 1e-06 
0.0 -0.1885 0 -2.0 1e-06 
0.0 -0.1884 0 -2.0 1e-06 
0.0 -0.1883 0 -2.0 1e-06 
0.0 -0.1882 0 -2.0 1e-06 
0.0 -0.1881 0 -2.0 1e-06 
0.0 -0.188 0 -2.0 1e-06 
0.0 -0.1879 0 -2.0 1e-06 
0.0 -0.1878 0 -2.0 1e-06 
0.0 -0.1877 0 -2.0 1e-06 
0.0 -0.1876 0 -2.0 1e-06 
0.0 -0.1875 0 -2.0 1e-06 
0.0 -0.1874 0 -2.0 1e-06 
0.0 -0.1873 0 -2.0 1e-06 
0.0 -0.1872 0 -2.0 1e-06 
0.0 -0.1871 0 -2.0 1e-06 
0.0 -0.187 0 -2.0 1e-06 
0.0 -0.1869 0 -2.0 1e-06 
0.0 -0.1868 0 -2.0 1e-06 
0.0 -0.1867 0 -2.0 1e-06 
0.0 -0.1866 0 -2.0 1e-06 
0.0 -0.1865 0 -2.0 1e-06 
0.0 -0.1864 0 -2.0 1e-06 
0.0 -0.1863 0 -2.0 1e-06 
0.0 -0.1862 0 -2.0 1e-06 
0.0 -0.1861 0 -2.0 1e-06 
0.0 -0.186 0 -2.0 1e-06 
0.0 -0.1859 0 -2.0 1e-06 
0.0 -0.1858 0 -2.0 1e-06 
0.0 -0.1857 0 -2.0 1e-06 
0.0 -0.1856 0 -2.0 1e-06 
0.0 -0.1855 0 -2.0 1e-06 
0.0 -0.1854 0 -2.0 1e-06 
0.0 -0.1853 0 -2.0 1e-06 
0.0 -0.1852 0 -2.0 1e-06 
0.0 -0.1851 0 -2.0 1e-06 
0.0 -0.185 0 -2.0 1e-06 
0.0 -0.1849 0 -2.0 1e-06 
0.0 -0.1848 0 -2.0 1e-06 
0.0 -0.1847 0 -2.0 1e-06 
0.0 -0.1846 0 -2.0 1e-06 
0.0 -0.1845 0 -2.0 1e-06 
0.0 -0.1844 0 -2.0 1e-06 
0.0 -0.1843 0 -2.0 1e-06 
0.0 -0.1842 0 -2.0 1e-06 
0.0 -0.1841 0 -2.0 1e-06 
0.0 -0.184 0 -2.0 1e-06 
0.0 -0.1839 0 -2.0 1e-06 
0.0 -0.1838 0 -2.0 1e-06 
0.0 -0.1837 0 -2.0 1e-06 
0.0 -0.1836 0 -2.0 1e-06 
0.0 -0.1835 0 -2.0 1e-06 
0.0 -0.1834 0 -2.0 1e-06 
0.0 -0.1833 0 -2.0 1e-06 
0.0 -0.1832 0 -2.0 1e-06 
0.0 -0.1831 0 -2.0 1e-06 
0.0 -0.183 0 -2.0 1e-06 
0.0 -0.1829 0 -2.0 1e-06 
0.0 -0.1828 0 -2.0 1e-06 
0.0 -0.1827 0 -2.0 1e-06 
0.0 -0.1826 0 -2.0 1e-06 
0.0 -0.1825 0 -2.0 1e-06 
0.0 -0.1824 0 -2.0 1e-06 
0.0 -0.1823 0 -2.0 1e-06 
0.0 -0.1822 0 -2.0 1e-06 
0.0 -0.1821 0 -2.0 1e-06 
0.0 -0.182 0 -2.0 1e-06 
0.0 -0.1819 0 -2.0 1e-06 
0.0 -0.1818 0 -2.0 1e-06 
0.0 -0.1817 0 -2.0 1e-06 
0.0 -0.1816 0 -2.0 1e-06 
0.0 -0.1815 0 -2.0 1e-06 
0.0 -0.1814 0 -2.0 1e-06 
0.0 -0.1813 0 -2.0 1e-06 
0.0 -0.1812 0 -2.0 1e-06 
0.0 -0.1811 0 -2.0 1e-06 
0.0 -0.181 0 -2.0 1e-06 
0.0 -0.1809 0 -2.0 1e-06 
0.0 -0.1808 0 -2.0 1e-06 
0.0 -0.1807 0 -2.0 1e-06 
0.0 -0.1806 0 -2.0 1e-06 
0.0 -0.1805 0 -2.0 1e-06 
0.0 -0.1804 0 -2.0 1e-06 
0.0 -0.1803 0 -2.0 1e-06 
0.0 -0.1802 0 -2.0 1e-06 
0.0 -0.1801 0 -2.0 1e-06 
0.0 -0.18 0 -2.0 1e-06 
0.0 -0.1799 0 -2.0 1e-06 
0.0 -0.1798 0 -2.0 1e-06 
0.0 -0.1797 0 -2.0 1e-06 
0.0 -0.1796 0 -2.0 1e-06 
0.0 -0.1795 0 -2.0 1e-06 
0.0 -0.1794 0 -2.0 1e-06 
0.0 -0.1793 0 -2.0 1e-06 
0.0 -0.1792 0 -2.0 1e-06 
0.0 -0.1791 0 -2.0 1e-06 
0.0 -0.179 0 -2.0 1e-06 
0.0 -0.1789 0 -2.0 1e-06 
0.0 -0.1788 0 -2.0 1e-06 
0.0 -0.1787 0 -2.0 1e-06 
0.0 -0.1786 0 -2.0 1e-06 
0.0 -0.1785 0 -2.0 1e-06 
0.0 -0.1784 0 -2.0 1e-06 
0.0 -0.1783 0 -2.0 1e-06 
0.0 -0.1782 0 -2.0 1e-06 
0.0 -0.1781 0 -2.0 1e-06 
0.0 -0.178 0 -2.0 1e-06 
0.0 -0.1779 0 -2.0 1e-06 
0.0 -0.1778 0 -2.0 1e-06 
0.0 -0.1777 0 -2.0 1e-06 
0.0 -0.1776 0 -2.0 1e-06 
0.0 -0.1775 0 -2.0 1e-06 
0.0 -0.1774 0 -2.0 1e-06 
0.0 -0.1773 0 -2.0 1e-06 
0.0 -0.1772 0 -2.0 1e-06 
0.0 -0.1771 0 -2.0 1e-06 
0.0 -0.177 0 -2.0 1e-06 
0.0 -0.1769 0 -2.0 1e-06 
0.0 -0.1768 0 -2.0 1e-06 
0.0 -0.1767 0 -2.0 1e-06 
0.0 -0.1766 0 -2.0 1e-06 
0.0 -0.1765 0 -2.0 1e-06 
0.0 -0.1764 0 -2.0 1e-06 
0.0 -0.1763 0 -2.0 1e-06 
0.0 -0.1762 0 -2.0 1e-06 
0.0 -0.1761 0 -2.0 1e-06 
0.0 -0.176 0 -2.0 1e-06 
0.0 -0.1759 0 -2.0 1e-06 
0.0 -0.1758 0 -2.0 1e-06 
0.0 -0.1757 0 -2.0 1e-06 
0.0 -0.1756 0 -2.0 1e-06 
0.0 -0.1755 0 -2.0 1e-06 
0.0 -0.1754 0 -2.0 1e-06 
0.0 -0.1753 0 -2.0 1e-06 
0.0 -0.1752 0 -2.0 1e-06 
0.0 -0.1751 0 -2.0 1e-06 
0.0 -0.175 0 -2.0 1e-06 
0.0 -0.1749 0 -2.0 1e-06 
0.0 -0.1748 0 -2.0 1e-06 
0.0 -0.1747 0 -2.0 1e-06 
0.0 -0.1746 0 -2.0 1e-06 
0.0 -0.1745 0 -2.0 1e-06 
0.0 -0.1744 0 -2.0 1e-06 
0.0 -0.1743 0 -2.0 1e-06 
0.0 -0.1742 0 -2.0 1e-06 
0.0 -0.1741 0 -2.0 1e-06 
0.0 -0.174 0 -2.0 1e-06 
0.0 -0.1739 0 -2.0 1e-06 
0.0 -0.1738 0 -2.0 1e-06 
0.0 -0.1737 0 -2.0 1e-06 
0.0 -0.1736 0 -2.0 1e-06 
0.0 -0.1735 0 -2.0 1e-06 
0.0 -0.1734 0 -2.0 1e-06 
0.0 -0.1733 0 -2.0 1e-06 
0.0 -0.1732 0 -2.0 1e-06 
0.0 -0.1731 0 -2.0 1e-06 
0.0 -0.173 0 -2.0 1e-06 
0.0 -0.1729 0 -2.0 1e-06 
0.0 -0.1728 0 -2.0 1e-06 
0.0 -0.1727 0 -2.0 1e-06 
0.0 -0.1726 0 -2.0 1e-06 
0.0 -0.1725 0 -2.0 1e-06 
0.0 -0.1724 0 -2.0 1e-06 
0.0 -0.1723 0 -2.0 1e-06 
0.0 -0.1722 0 -2.0 1e-06 
0.0 -0.1721 0 -2.0 1e-06 
0.0 -0.172 0 -2.0 1e-06 
0.0 -0.1719 0 -2.0 1e-06 
0.0 -0.1718 0 -2.0 1e-06 
0.0 -0.1717 0 -2.0 1e-06 
0.0 -0.1716 0 -2.0 1e-06 
0.0 -0.1715 0 -2.0 1e-06 
0.0 -0.1714 0 -2.0 1e-06 
0.0 -0.1713 0 -2.0 1e-06 
0.0 -0.1712 0 -2.0 1e-06 
0.0 -0.1711 0 -2.0 1e-06 
0.0 -0.171 0 -2.0 1e-06 
0.0 -0.1709 0 -2.0 1e-06 
0.0 -0.1708 0 -2.0 1e-06 
0.0 -0.1707 0 -2.0 1e-06 
0.0 -0.1706 0 -2.0 1e-06 
0.0 -0.1705 0 -2.0 1e-06 
0.0 -0.1704 0 -2.0 1e-06 
0.0 -0.1703 0 -2.0 1e-06 
0.0 -0.1702 0 -2.0 1e-06 
0.0 -0.1701 0 -2.0 1e-06 
0.0 -0.17 0 -2.0 1e-06 
0.0 -0.1699 0 -2.0 1e-06 
0.0 -0.1698 0 -2.0 1e-06 
0.0 -0.1697 0 -2.0 1e-06 
0.0 -0.1696 0 -2.0 1e-06 
0.0 -0.1695 0 -2.0 1e-06 
0.0 -0.1694 0 -2.0 1e-06 
0.0 -0.1693 0 -2.0 1e-06 
0.0 -0.1692 0 -2.0 1e-06 
0.0 -0.1691 0 -2.0 1e-06 
0.0 -0.169 0 -2.0 1e-06 
0.0 -0.1689 0 -2.0 1e-06 
0.0 -0.1688 0 -2.0 1e-06 
0.0 -0.1687 0 -2.0 1e-06 
0.0 -0.1686 0 -2.0 1e-06 
0.0 -0.1685 0 -2.0 1e-06 
0.0 -0.1684 0 -2.0 1e-06 
0.0 -0.1683 0 -2.0 1e-06 
0.0 -0.1682 0 -2.0 1e-06 
0.0 -0.1681 0 -2.0 1e-06 
0.0 -0.168 0 -2.0 1e-06 
0.0 -0.1679 0 -2.0 1e-06 
0.0 -0.1678 0 -2.0 1e-06 
0.0 -0.1677 0 -2.0 1e-06 
0.0 -0.1676 0 -2.0 1e-06 
0.0 -0.1675 0 -2.0 1e-06 
0.0 -0.1674 0 -2.0 1e-06 
0.0 -0.1673 0 -2.0 1e-06 
0.0 -0.1672 0 -2.0 1e-06 
0.0 -0.1671 0 -2.0 1e-06 
0.0 -0.167 0 -2.0 1e-06 
0.0 -0.1669 0 -2.0 1e-06 
0.0 -0.1668 0 -2.0 1e-06 
0.0 -0.1667 0 -2.0 1e-06 
0.0 -0.1666 0 -2.0 1e-06 
0.0 -0.1665 0 -2.0 1e-06 
0.0 -0.1664 0 -2.0 1e-06 
0.0 -0.1663 0 -2.0 1e-06 
0.0 -0.1662 0 -2.0 1e-06 
0.0 -0.1661 0 -2.0 1e-06 
0.0 -0.166 0 -2.0 1e-06 
0.0 -0.1659 0 -2.0 1e-06 
0.0 -0.1658 0 -2.0 1e-06 
0.0 -0.1657 0 -2.0 1e-06 
0.0 -0.1656 0 -2.0 1e-06 
0.0 -0.1655 0 -2.0 1e-06 
0.0 -0.1654 0 -2.0 1e-06 
0.0 -0.1653 0 -2.0 1e-06 
0.0 -0.1652 0 -2.0 1e-06 
0.0 -0.1651 0 -2.0 1e-06 
0.0 -0.165 0 -2.0 1e-06 
0.0 -0.1649 0 -2.0 1e-06 
0.0 -0.1648 0 -2.0 1e-06 
0.0 -0.1647 0 -2.0 1e-06 
0.0 -0.1646 0 -2.0 1e-06 
0.0 -0.1645 0 -2.0 1e-06 
0.0 -0.1644 0 -2.0 1e-06 
0.0 -0.1643 0 -2.0 1e-06 
0.0 -0.1642 0 -2.0 1e-06 
0.0 -0.1641 0 -2.0 1e-06 
0.0 -0.164 0 -2.0 1e-06 
0.0 -0.1639 0 -2.0 1e-06 
0.0 -0.1638 0 -2.0 1e-06 
0.0 -0.1637 0 -2.0 1e-06 
0.0 -0.1636 0 -2.0 1e-06 
0.0 -0.1635 0 -2.0 1e-06 
0.0 -0.1634 0 -2.0 1e-06 
0.0 -0.1633 0 -2.0 1e-06 
0.0 -0.1632 0 -2.0 1e-06 
0.0 -0.1631 0 -2.0 1e-06 
0.0 -0.163 0 -2.0 1e-06 
0.0 -0.1629 0 -2.0 1e-06 
0.0 -0.1628 0 -2.0 1e-06 
0.0 -0.1627 0 -2.0 1e-06 
0.0 -0.1626 0 -2.0 1e-06 
0.0 -0.1625 0 -2.0 1e-06 
0.0 -0.1624 0 -2.0 1e-06 
0.0 -0.1623 0 -2.0 1e-06 
0.0 -0.1622 0 -2.0 1e-06 
0.0 -0.1621 0 -2.0 1e-06 
0.0 -0.162 0 -2.0 1e-06 
0.0 -0.1619 0 -2.0 1e-06 
0.0 -0.1618 0 -2.0 1e-06 
0.0 -0.1617 0 -2.0 1e-06 
0.0 -0.1616 0 -2.0 1e-06 
0.0 -0.1615 0 -2.0 1e-06 
0.0 -0.1614 0 -2.0 1e-06 
0.0 -0.1613 0 -2.0 1e-06 
0.0 -0.1612 0 -2.0 1e-06 
0.0 -0.1611 0 -2.0 1e-06 
0.0 -0.161 0 -2.0 1e-06 
0.0 -0.1609 0 -2.0 1e-06 
0.0 -0.1608 0 -2.0 1e-06 
0.0 -0.1607 0 -2.0 1e-06 
0.0 -0.1606 0 -2.0 1e-06 
0.0 -0.1605 0 -2.0 1e-06 
0.0 -0.1604 0 -2.0 1e-06 
0.0 -0.1603 0 -2.0 1e-06 
0.0 -0.1602 0 -2.0 1e-06 
0.0 -0.1601 0 -2.0 1e-06 
0.0 -0.16 0 -2.0 1e-06 
0.0 -0.1599 0 -2.0 1e-06 
0.0 -0.1598 0 -2.0 1e-06 
0.0 -0.1597 0 -2.0 1e-06 
0.0 -0.1596 0 -2.0 1e-06 
0.0 -0.1595 0 -2.0 1e-06 
0.0 -0.1594 0 -2.0 1e-06 
0.0 -0.1593 0 -2.0 1e-06 
0.0 -0.1592 0 -2.0 1e-06 
0.0 -0.1591 0 -2.0 1e-06 
0.0 -0.159 0 -2.0 1e-06 
0.0 -0.1589 0 -2.0 1e-06 
0.0 -0.1588 0 -2.0 1e-06 
0.0 -0.1587 0 -2.0 1e-06 
0.0 -0.1586 0 -2.0 1e-06 
0.0 -0.1585 0 -2.0 1e-06 
0.0 -0.1584 0 -2.0 1e-06 
0.0 -0.1583 0 -2.0 1e-06 
0.0 -0.1582 0 -2.0 1e-06 
0.0 -0.1581 0 -2.0 1e-06 
0.0 -0.158 0 -2.0 1e-06 
0.0 -0.1579 0 -2.0 1e-06 
0.0 -0.1578 0 -2.0 1e-06 
0.0 -0.1577 0 -2.0 1e-06 
0.0 -0.1576 0 -2.0 1e-06 
0.0 -0.1575 0 -2.0 1e-06 
0.0 -0.1574 0 -2.0 1e-06 
0.0 -0.1573 0 -2.0 1e-06 
0.0 -0.1572 0 -2.0 1e-06 
0.0 -0.1571 0 -2.0 1e-06 
0.0 -0.157 0 -2.0 1e-06 
0.0 -0.1569 0 -2.0 1e-06 
0.0 -0.1568 0 -2.0 1e-06 
0.0 -0.1567 0 -2.0 1e-06 
0.0 -0.1566 0 -2.0 1e-06 
0.0 -0.1565 0 -2.0 1e-06 
0.0 -0.1564 0 -2.0 1e-06 
0.0 -0.1563 0 -2.0 1e-06 
0.0 -0.1562 0 -2.0 1e-06 
0.0 -0.1561 0 -2.0 1e-06 
0.0 -0.156 0 -2.0 1e-06 
0.0 -0.1559 0 -2.0 1e-06 
0.0 -0.1558 0 -2.0 1e-06 
0.0 -0.1557 0 -2.0 1e-06 
0.0 -0.1556 0 -2.0 1e-06 
0.0 -0.1555 0 -2.0 1e-06 
0.0 -0.1554 0 -2.0 1e-06 
0.0 -0.1553 0 -2.0 1e-06 
0.0 -0.1552 0 -2.0 1e-06 
0.0 -0.1551 0 -2.0 1e-06 
0.0 -0.155 0 -2.0 1e-06 
0.0 -0.1549 0 -2.0 1e-06 
0.0 -0.1548 0 -2.0 1e-06 
0.0 -0.1547 0 -2.0 1e-06 
0.0 -0.1546 0 -2.0 1e-06 
0.0 -0.1545 0 -2.0 1e-06 
0.0 -0.1544 0 -2.0 1e-06 
0.0 -0.1543 0 -2.0 1e-06 
0.0 -0.1542 0 -2.0 1e-06 
0.0 -0.1541 0 -2.0 1e-06 
0.0 -0.154 0 -2.0 1e-06 
0.0 -0.1539 0 -2.0 1e-06 
0.0 -0.1538 0 -2.0 1e-06 
0.0 -0.1537 0 -2.0 1e-06 
0.0 -0.1536 0 -2.0 1e-06 
0.0 -0.1535 0 -2.0 1e-06 
0.0 -0.1534 0 -2.0 1e-06 
0.0 -0.1533 0 -2.0 1e-06 
0.0 -0.1532 0 -2.0 1e-06 
0.0 -0.1531 0 -2.0 1e-06 
0.0 -0.153 0 -2.0 1e-06 
0.0 -0.1529 0 -2.0 1e-06 
0.0 -0.1528 0 -2.0 1e-06 
0.0 -0.1527 0 -2.0 1e-06 
0.0 -0.1526 0 -2.0 1e-06 
0.0 -0.1525 0 -2.0 1e-06 
0.0 -0.1524 0 -2.0 1e-06 
0.0 -0.1523 0 -2.0 1e-06 
0.0 -0.1522 0 -2.0 1e-06 
0.0 -0.1521 0 -2.0 1e-06 
0.0 -0.152 0 -2.0 1e-06 
0.0 -0.1519 0 -2.0 1e-06 
0.0 -0.1518 0 -2.0 1e-06 
0.0 -0.1517 0 -2.0 1e-06 
0.0 -0.1516 0 -2.0 1e-06 
0.0 -0.1515 0 -2.0 1e-06 
0.0 -0.1514 0 -2.0 1e-06 
0.0 -0.1513 0 -2.0 1e-06 
0.0 -0.1512 0 -2.0 1e-06 
0.0 -0.1511 0 -2.0 1e-06 
0.0 -0.151 0 -2.0 1e-06 
0.0 -0.1509 0 -2.0 1e-06 
0.0 -0.1508 0 -2.0 1e-06 
0.0 -0.1507 0 -2.0 1e-06 
0.0 -0.1506 0 -2.0 1e-06 
0.0 -0.1505 0 -2.0 1e-06 
0.0 -0.1504 0 -2.0 1e-06 
0.0 -0.1503 0 -2.0 1e-06 
0.0 -0.1502 0 -2.0 1e-06 
0.0 -0.1501 0 -2.0 1e-06 
0.0 -0.15 0 -2.0 1e-06 
0.0 -0.1499 0 -2.0 1e-06 
0.0 -0.1498 0 -2.0 1e-06 
0.0 -0.1497 0 -2.0 1e-06 
0.0 -0.1496 0 -2.0 1e-06 
0.0 -0.1495 0 -2.0 1e-06 
0.0 -0.1494 0 -2.0 1e-06 
0.0 -0.1493 0 -2.0 1e-06 
0.0 -0.1492 0 -2.0 1e-06 
0.0 -0.1491 0 -2.0 1e-06 
0.0 -0.149 0 -2.0 1e-06 
0.0 -0.1489 0 -2.0 1e-06 
0.0 -0.1488 0 -2.0 1e-06 
0.0 -0.1487 0 -2.0 1e-06 
0.0 -0.1486 0 -2.0 1e-06 
0.0 -0.1485 0 -2.0 1e-06 
0.0 -0.1484 0 -2.0 1e-06 
0.0 -0.1483 0 -2.0 1e-06 
0.0 -0.1482 0 -2.0 1e-06 
0.0 -0.1481 0 -2.0 1e-06 
0.0 -0.148 0 -2.0 1e-06 
0.0 -0.1479 0 -2.0 1e-06 
0.0 -0.1478 0 -2.0 1e-06 
0.0 -0.1477 0 -2.0 1e-06 
0.0 -0.1476 0 -2.0 1e-06 
0.0 -0.1475 0 -2.0 1e-06 
0.0 -0.1474 0 -2.0 1e-06 
0.0 -0.1473 0 -2.0 1e-06 
0.0 -0.1472 0 -2.0 1e-06 
0.0 -0.1471 0 -2.0 1e-06 
0.0 -0.147 0 -2.0 1e-06 
0.0 -0.1469 0 -2.0 1e-06 
0.0 -0.1468 0 -2.0 1e-06 
0.0 -0.1467 0 -2.0 1e-06 
0.0 -0.1466 0 -2.0 1e-06 
0.0 -0.1465 0 -2.0 1e-06 
0.0 -0.1464 0 -2.0 1e-06 
0.0 -0.1463 0 -2.0 1e-06 
0.0 -0.1462 0 -2.0 1e-06 
0.0 -0.1461 0 -2.0 1e-06 
0.0 -0.146 0 -2.0 1e-06 
0.0 -0.1459 0 -2.0 1e-06 
0.0 -0.1458 0 -2.0 1e-06 
0.0 -0.1457 0 -2.0 1e-06 
0.0 -0.1456 0 -2.0 1e-06 
0.0 -0.1455 0 -2.0 1e-06 
0.0 -0.1454 0 -2.0 1e-06 
0.0 -0.1453 0 -2.0 1e-06 
0.0 -0.1452 0 -2.0 1e-06 
0.0 -0.1451 0 -2.0 1e-06 
0.0 -0.145 0 -2.0 1e-06 
0.0 -0.1449 0 -2.0 1e-06 
0.0 -0.1448 0 -2.0 1e-06 
0.0 -0.1447 0 -2.0 1e-06 
0.0 -0.1446 0 -2.0 1e-06 
0.0 -0.1445 0 -2.0 1e-06 
0.0 -0.1444 0 -2.0 1e-06 
0.0 -0.1443 0 -2.0 1e-06 
0.0 -0.1442 0 -2.0 1e-06 
0.0 -0.1441 0 -2.0 1e-06 
0.0 -0.144 0 -2.0 1e-06 
0.0 -0.1439 0 -2.0 1e-06 
0.0 -0.1438 0 -2.0 1e-06 
0.0 -0.1437 0 -2.0 1e-06 
0.0 -0.1436 0 -2.0 1e-06 
0.0 -0.1435 0 -2.0 1e-06 
0.0 -0.1434 0 -2.0 1e-06 
0.0 -0.1433 0 -2.0 1e-06 
0.0 -0.1432 0 -2.0 1e-06 
0.0 -0.1431 0 -2.0 1e-06 
0.0 -0.143 0 -2.0 1e-06 
0.0 -0.1429 0 -2.0 1e-06 
0.0 -0.1428 0 -2.0 1e-06 
0.0 -0.1427 0 -2.0 1e-06 
0.0 -0.1426 0 -2.0 1e-06 
0.0 -0.1425 0 -2.0 1e-06 
0.0 -0.1424 0 -2.0 1e-06 
0.0 -0.1423 0 -2.0 1e-06 
0.0 -0.1422 0 -2.0 1e-06 
0.0 -0.1421 0 -2.0 1e-06 
0.0 -0.142 0 -2.0 1e-06 
0.0 -0.1419 0 -2.0 1e-06 
0.0 -0.1418 0 -2.0 1e-06 
0.0 -0.1417 0 -2.0 1e-06 
0.0 -0.1416 0 -2.0 1e-06 
0.0 -0.1415 0 -2.0 1e-06 
0.0 -0.1414 0 -2.0 1e-06 
0.0 -0.1413 0 -2.0 1e-06 
0.0 -0.1412 0 -2.0 1e-06 
0.0 -0.1411 0 -2.0 1e-06 
0.0 -0.141 0 -2.0 1e-06 
0.0 -0.1409 0 -2.0 1e-06 
0.0 -0.1408 0 -2.0 1e-06 
0.0 -0.1407 0 -2.0 1e-06 
0.0 -0.1406 0 -2.0 1e-06 
0.0 -0.1405 0 -2.0 1e-06 
0.0 -0.1404 0 -2.0 1e-06 
0.0 -0.1403 0 -2.0 1e-06 
0.0 -0.1402 0 -2.0 1e-06 
0.0 -0.1401 0 -2.0 1e-06 
0.0 -0.14 0 -2.0 1e-06 
0.0 -0.1399 0 -2.0 1e-06 
0.0 -0.1398 0 -2.0 1e-06 
0.0 -0.1397 0 -2.0 1e-06 
0.0 -0.1396 0 -2.0 1e-06 
0.0 -0.1395 0 -2.0 1e-06 
0.0 -0.1394 0 -2.0 1e-06 
0.0 -0.1393 0 -2.0 1e-06 
0.0 -0.1392 0 -2.0 1e-06 
0.0 -0.1391 0 -2.0 1e-06 
0.0 -0.139 0 -2.0 1e-06 
0.0 -0.1389 0 -2.0 1e-06 
0.0 -0.1388 0 -2.0 1e-06 
0.0 -0.1387 0 -2.0 1e-06 
0.0 -0.1386 0 -2.0 1e-06 
0.0 -0.1385 0 -2.0 1e-06 
0.0 -0.1384 0 -2.0 1e-06 
0.0 -0.1383 0 -2.0 1e-06 
0.0 -0.1382 0 -2.0 1e-06 
0.0 -0.1381 0 -2.0 1e-06 
0.0 -0.138 0 -2.0 1e-06 
0.0 -0.1379 0 -2.0 1e-06 
0.0 -0.1378 0 -2.0 1e-06 
0.0 -0.1377 0 -2.0 1e-06 
0.0 -0.1376 0 -2.0 1e-06 
0.0 -0.1375 0 -2.0 1e-06 
0.0 -0.1374 0 -2.0 1e-06 
0.0 -0.1373 0 -2.0 1e-06 
0.0 -0.1372 0 -2.0 1e-06 
0.0 -0.1371 0 -2.0 1e-06 
0.0 -0.137 0 -2.0 1e-06 
0.0 -0.1369 0 -2.0 1e-06 
0.0 -0.1368 0 -2.0 1e-06 
0.0 -0.1367 0 -2.0 1e-06 
0.0 -0.1366 0 -2.0 1e-06 
0.0 -0.1365 0 -2.0 1e-06 
0.0 -0.1364 0 -2.0 1e-06 
0.0 -0.1363 0 -2.0 1e-06 
0.0 -0.1362 0 -2.0 1e-06 
0.0 -0.1361 0 -2.0 1e-06 
0.0 -0.136 0 -2.0 1e-06 
0.0 -0.1359 0 -2.0 1e-06 
0.0 -0.1358 0 -2.0 1e-06 
0.0 -0.1357 0 -2.0 1e-06 
0.0 -0.1356 0 -2.0 1e-06 
0.0 -0.1355 0 -2.0 1e-06 
0.0 -0.1354 0 -2.0 1e-06 
0.0 -0.1353 0 -2.0 1e-06 
0.0 -0.1352 0 -2.0 1e-06 
0.0 -0.1351 0 -2.0 1e-06 
0.0 -0.135 0 -2.0 1e-06 
0.0 -0.1349 0 -2.0 1e-06 
0.0 -0.1348 0 -2.0 1e-06 
0.0 -0.1347 0 -2.0 1e-06 
0.0 -0.1346 0 -2.0 1e-06 
0.0 -0.1345 0 -2.0 1e-06 
0.0 -0.1344 0 -2.0 1e-06 
0.0 -0.1343 0 -2.0 1e-06 
0.0 -0.1342 0 -2.0 1e-06 
0.0 -0.1341 0 -2.0 1e-06 
0.0 -0.134 0 -2.0 1e-06 
0.0 -0.1339 0 -2.0 1e-06 
0.0 -0.1338 0 -2.0 1e-06 
0.0 -0.1337 0 -2.0 1e-06 
0.0 -0.1336 0 -2.0 1e-06 
0.0 -0.1335 0 -2.0 1e-06 
0.0 -0.1334 0 -2.0 1e-06 
0.0 -0.1333 0 -2.0 1e-06 
0.0 -0.1332 0 -2.0 1e-06 
0.0 -0.1331 0 -2.0 1e-06 
0.0 -0.133 0 -2.0 1e-06 
0.0 -0.1329 0 -2.0 1e-06 
0.0 -0.1328 0 -2.0 1e-06 
0.0 -0.1327 0 -2.0 1e-06 
0.0 -0.1326 0 -2.0 1e-06 
0.0 -0.1325 0 -2.0 1e-06 
0.0 -0.1324 0 -2.0 1e-06 
0.0 -0.1323 0 -2.0 1e-06 
0.0 -0.1322 0 -2.0 1e-06 
0.0 -0.1321 0 -2.0 1e-06 
0.0 -0.132 0 -2.0 1e-06 
0.0 -0.1319 0 -2.0 1e-06 
0.0 -0.1318 0 -2.0 1e-06 
0.0 -0.1317 0 -2.0 1e-06 
0.0 -0.1316 0 -2.0 1e-06 
0.0 -0.1315 0 -2.0 1e-06 
0.0 -0.1314 0 -2.0 1e-06 
0.0 -0.1313 0 -2.0 1e-06 
0.0 -0.1312 0 -2.0 1e-06 
0.0 -0.1311 0 -2.0 1e-06 
0.0 -0.131 0 -2.0 1e-06 
0.0 -0.1309 0 -2.0 1e-06 
0.0 -0.1308 0 -2.0 1e-06 
0.0 -0.1307 0 -2.0 1e-06 
0.0 -0.1306 0 -2.0 1e-06 
0.0 -0.1305 0 -2.0 1e-06 
0.0 -0.1304 0 -2.0 1e-06 
0.0 -0.1303 0 -2.0 1e-06 
0.0 -0.1302 0 -2.0 1e-06 
0.0 -0.1301 0 -2.0 1e-06 
0.0 -0.13 0 -2.0 1e-06 
0.0 -0.1299 0 -2.0 1e-06 
0.0 -0.1298 0 -2.0 1e-06 
0.0 -0.1297 0 -2.0 1e-06 
0.0 -0.1296 0 -2.0 1e-06 
0.0 -0.1295 0 -2.0 1e-06 
0.0 -0.1294 0 -2.0 1e-06 
0.0 -0.1293 0 -2.0 1e-06 
0.0 -0.1292 0 -2.0 1e-06 
0.0 -0.1291 0 -2.0 1e-06 
0.0 -0.129 0 -2.0 1e-06 
0.0 -0.1289 0 -2.0 1e-06 
0.0 -0.1288 0 -2.0 1e-06 
0.0 -0.1287 0 -2.0 1e-06 
0.0 -0.1286 0 -2.0 1e-06 
0.0 -0.1285 0 -2.0 1e-06 
0.0 -0.1284 0 -2.0 1e-06 
0.0 -0.1283 0 -2.0 1e-06 
0.0 -0.1282 0 -2.0 1e-06 
0.0 -0.1281 0 -2.0 1e-06 
0.0 -0.128 0 -2.0 1e-06 
0.0 -0.1279 0 -2.0 1e-06 
0.0 -0.1278 0 -2.0 1e-06 
0.0 -0.1277 0 -2.0 1e-06 
0.0 -0.1276 0 -2.0 1e-06 
0.0 -0.1275 0 -2.0 1e-06 
0.0 -0.1274 0 -2.0 1e-06 
0.0 -0.1273 0 -2.0 1e-06 
0.0 -0.1272 0 -2.0 1e-06 
0.0 -0.1271 0 -2.0 1e-06 
0.0 -0.127 0 -2.0 1e-06 
0.0 -0.1269 0 -2.0 1e-06 
0.0 -0.1268 0 -2.0 1e-06 
0.0 -0.1267 0 -2.0 1e-06 
0.0 -0.1266 0 -2.0 1e-06 
0.0 -0.1265 0 -2.0 1e-06 
0.0 -0.1264 0 -2.0 1e-06 
0.0 -0.1263 0 -2.0 1e-06 
0.0 -0.1262 0 -2.0 1e-06 
0.0 -0.1261 0 -2.0 1e-06 
0.0 -0.126 0 -2.0 1e-06 
0.0 -0.1259 0 -2.0 1e-06 
0.0 -0.1258 0 -2.0 1e-06 
0.0 -0.1257 0 -2.0 1e-06 
0.0 -0.1256 0 -2.0 1e-06 
0.0 -0.1255 0 -2.0 1e-06 
0.0 -0.1254 0 -2.0 1e-06 
0.0 -0.1253 0 -2.0 1e-06 
0.0 -0.1252 0 -2.0 1e-06 
0.0 -0.1251 0 -2.0 1e-06 
0.0 -0.125 0 -2.0 1e-06 
0.0 -0.1249 0 -2.0 1e-06 
0.0 -0.1248 0 -2.0 1e-06 
0.0 -0.1247 0 -2.0 1e-06 
0.0 -0.1246 0 -2.0 1e-06 
0.0 -0.1245 0 -2.0 1e-06 
0.0 -0.1244 0 -2.0 1e-06 
0.0 -0.1243 0 -2.0 1e-06 
0.0 -0.1242 0 -2.0 1e-06 
0.0 -0.1241 0 -2.0 1e-06 
0.0 -0.124 0 -2.0 1e-06 
0.0 -0.1239 0 -2.0 1e-06 
0.0 -0.1238 0 -2.0 1e-06 
0.0 -0.1237 0 -2.0 1e-06 
0.0 -0.1236 0 -2.0 1e-06 
0.0 -0.1235 0 -2.0 1e-06 
0.0 -0.1234 0 -2.0 1e-06 
0.0 -0.1233 0 -2.0 1e-06 
0.0 -0.1232 0 -2.0 1e-06 
0.0 -0.1231 0 -2.0 1e-06 
0.0 -0.123 0 -2.0 1e-06 
0.0 -0.1229 0 -2.0 1e-06 
0.0 -0.1228 0 -2.0 1e-06 
0.0 -0.1227 0 -2.0 1e-06 
0.0 -0.1226 0 -2.0 1e-06 
0.0 -0.1225 0 -2.0 1e-06 
0.0 -0.1224 0 -2.0 1e-06 
0.0 -0.1223 0 -2.0 1e-06 
0.0 -0.1222 0 -2.0 1e-06 
0.0 -0.1221 0 -2.0 1e-06 
0.0 -0.122 0 -2.0 1e-06 
0.0 -0.1219 0 -2.0 1e-06 
0.0 -0.1218 0 -2.0 1e-06 
0.0 -0.1217 0 -2.0 1e-06 
0.0 -0.1216 0 -2.0 1e-06 
0.0 -0.1215 0 -2.0 1e-06 
0.0 -0.1214 0 -2.0 1e-06 
0.0 -0.1213 0 -2.0 1e-06 
0.0 -0.1212 0 -2.0 1e-06 
0.0 -0.1211 0 -2.0 1e-06 
0.0 -0.121 0 -2.0 1e-06 
0.0 -0.1209 0 -2.0 1e-06 
0.0 -0.1208 0 -2.0 1e-06 
0.0 -0.1207 0 -2.0 1e-06 
0.0 -0.1206 0 -2.0 1e-06 
0.0 -0.1205 0 -2.0 1e-06 
0.0 -0.1204 0 -2.0 1e-06 
0.0 -0.1203 0 -2.0 1e-06 
0.0 -0.1202 0 -2.0 1e-06 
0.0 -0.1201 0 -2.0 1e-06 
0.0 -0.12 0 -2.0 1e-06 
0.0 -0.1199 0 -2.0 1e-06 
0.0 -0.1198 0 -2.0 1e-06 
0.0 -0.1197 0 -2.0 1e-06 
0.0 -0.1196 0 -2.0 1e-06 
0.0 -0.1195 0 -2.0 1e-06 
0.0 -0.1194 0 -2.0 1e-06 
0.0 -0.1193 0 -2.0 1e-06 
0.0 -0.1192 0 -2.0 1e-06 
0.0 -0.1191 0 -2.0 1e-06 
0.0 -0.119 0 -2.0 1e-06 
0.0 -0.1189 0 -2.0 1e-06 
0.0 -0.1188 0 -2.0 1e-06 
0.0 -0.1187 0 -2.0 1e-06 
0.0 -0.1186 0 -2.0 1e-06 
0.0 -0.1185 0 -2.0 1e-06 
0.0 -0.1184 0 -2.0 1e-06 
0.0 -0.1183 0 -2.0 1e-06 
0.0 -0.1182 0 -2.0 1e-06 
0.0 -0.1181 0 -2.0 1e-06 
0.0 -0.118 0 -2.0 1e-06 
0.0 -0.1179 0 -2.0 1e-06 
0.0 -0.1178 0 -2.0 1e-06 
0.0 -0.1177 0 -2.0 1e-06 
0.0 -0.1176 0 -2.0 1e-06 
0.0 -0.1175 0 -2.0 1e-06 
0.0 -0.1174 0 -2.0 1e-06 
0.0 -0.1173 0 -2.0 1e-06 
0.0 -0.1172 0 -2.0 1e-06 
0.0 -0.1171 0 -2.0 1e-06 
0.0 -0.117 0 -2.0 1e-06 
0.0 -0.1169 0 -2.0 1e-06 
0.0 -0.1168 0 -2.0 1e-06 
0.0 -0.1167 0 -2.0 1e-06 
0.0 -0.1166 0 -2.0 1e-06 
0.0 -0.1165 0 -2.0 1e-06 
0.0 -0.1164 0 -2.0 1e-06 
0.0 -0.1163 0 -2.0 1e-06 
0.0 -0.1162 0 -2.0 1e-06 
0.0 -0.1161 0 -2.0 1e-06 
0.0 -0.116 0 -2.0 1e-06 
0.0 -0.1159 0 -2.0 1e-06 
0.0 -0.1158 0 -2.0 1e-06 
0.0 -0.1157 0 -2.0 1e-06 
0.0 -0.1156 0 -2.0 1e-06 
0.0 -0.1155 0 -2.0 1e-06 
0.0 -0.1154 0 -2.0 1e-06 
0.0 -0.1153 0 -2.0 1e-06 
0.0 -0.1152 0 -2.0 1e-06 
0.0 -0.1151 0 -2.0 1e-06 
0.0 -0.115 0 -2.0 1e-06 
0.0 -0.1149 0 -2.0 1e-06 
0.0 -0.1148 0 -2.0 1e-06 
0.0 -0.1147 0 -2.0 1e-06 
0.0 -0.1146 0 -2.0 1e-06 
0.0 -0.1145 0 -2.0 1e-06 
0.0 -0.1144 0 -2.0 1e-06 
0.0 -0.1143 0 -2.0 1e-06 
0.0 -0.1142 0 -2.0 1e-06 
0.0 -0.1141 0 -2.0 1e-06 
0.0 -0.114 0 -2.0 1e-06 
0.0 -0.1139 0 -2.0 1e-06 
0.0 -0.1138 0 -2.0 1e-06 
0.0 -0.1137 0 -2.0 1e-06 
0.0 -0.1136 0 -2.0 1e-06 
0.0 -0.1135 0 -2.0 1e-06 
0.0 -0.1134 0 -2.0 1e-06 
0.0 -0.1133 0 -2.0 1e-06 
0.0 -0.1132 0 -2.0 1e-06 
0.0 -0.1131 0 -2.0 1e-06 
0.0 -0.113 0 -2.0 1e-06 
0.0 -0.1129 0 -2.0 1e-06 
0.0 -0.1128 0 -2.0 1e-06 
0.0 -0.1127 0 -2.0 1e-06 
0.0 -0.1126 0 -2.0 1e-06 
0.0 -0.1125 0 -2.0 1e-06 
0.0 -0.1124 0 -2.0 1e-06 
0.0 -0.1123 0 -2.0 1e-06 
0.0 -0.1122 0 -2.0 1e-06 
0.0 -0.1121 0 -2.0 1e-06 
0.0 -0.112 0 -2.0 1e-06 
0.0 -0.1119 0 -2.0 1e-06 
0.0 -0.1118 0 -2.0 1e-06 
0.0 -0.1117 0 -2.0 1e-06 
0.0 -0.1116 0 -2.0 1e-06 
0.0 -0.1115 0 -2.0 1e-06 
0.0 -0.1114 0 -2.0 1e-06 
0.0 -0.1113 0 -2.0 1e-06 
0.0 -0.1112 0 -2.0 1e-06 
0.0 -0.1111 0 -2.0 1e-06 
0.0 -0.111 0 -2.0 1e-06 
0.0 -0.1109 0 -2.0 1e-06 
0.0 -0.1108 0 -2.0 1e-06 
0.0 -0.1107 0 -2.0 1e-06 
0.0 -0.1106 0 -2.0 1e-06 
0.0 -0.1105 0 -2.0 1e-06 
0.0 -0.1104 0 -2.0 1e-06 
0.0 -0.1103 0 -2.0 1e-06 
0.0 -0.1102 0 -2.0 1e-06 
0.0 -0.1101 0 -2.0 1e-06 
0.0 -0.11 0 -2.0 1e-06 
0.0 -0.1099 0 -2.0 1e-06 
0.0 -0.1098 0 -2.0 1e-06 
0.0 -0.1097 0 -2.0 1e-06 
0.0 -0.1096 0 -2.0 1e-06 
0.0 -0.1095 0 -2.0 1e-06 
0.0 -0.1094 0 -2.0 1e-06 
0.0 -0.1093 0 -2.0 1e-06 
0.0 -0.1092 0 -2.0 1e-06 
0.0 -0.1091 0 -2.0 1e-06 
0.0 -0.109 0 -2.0 1e-06 
0.0 -0.1089 0 -2.0 1e-06 
0.0 -0.1088 0 -2.0 1e-06 
0.0 -0.1087 0 -2.0 1e-06 
0.0 -0.1086 0 -2.0 1e-06 
0.0 -0.1085 0 -2.0 1e-06 
0.0 -0.1084 0 -2.0 1e-06 
0.0 -0.1083 0 -2.0 1e-06 
0.0 -0.1082 0 -2.0 1e-06 
0.0 -0.1081 0 -2.0 1e-06 
0.0 -0.108 0 -2.0 1e-06 
0.0 -0.1079 0 -2.0 1e-06 
0.0 -0.1078 0 -2.0 1e-06 
0.0 -0.1077 0 -2.0 1e-06 
0.0 -0.1076 0 -2.0 1e-06 
0.0 -0.1075 0 -2.0 1e-06 
0.0 -0.1074 0 -2.0 1e-06 
0.0 -0.1073 0 -2.0 1e-06 
0.0 -0.1072 0 -2.0 1e-06 
0.0 -0.1071 0 -2.0 1e-06 
0.0 -0.107 0 -2.0 1e-06 
0.0 -0.1069 0 -2.0 1e-06 
0.0 -0.1068 0 -2.0 1e-06 
0.0 -0.1067 0 -2.0 1e-06 
0.0 -0.1066 0 -2.0 1e-06 
0.0 -0.1065 0 -2.0 1e-06 
0.0 -0.1064 0 -2.0 1e-06 
0.0 -0.1063 0 -2.0 1e-06 
0.0 -0.1062 0 -2.0 1e-06 
0.0 -0.1061 0 -2.0 1e-06 
0.0 -0.106 0 -2.0 1e-06 
0.0 -0.1059 0 -2.0 1e-06 
0.0 -0.1058 0 -2.0 1e-06 
0.0 -0.1057 0 -2.0 1e-06 
0.0 -0.1056 0 -2.0 1e-06 
0.0 -0.1055 0 -2.0 1e-06 
0.0 -0.1054 0 -2.0 1e-06 
0.0 -0.1053 0 -2.0 1e-06 
0.0 -0.1052 0 -2.0 1e-06 
0.0 -0.1051 0 -2.0 1e-06 
0.0 -0.105 0 -2.0 1e-06 
0.0 -0.1049 0 -2.0 1e-06 
0.0 -0.1048 0 -2.0 1e-06 
0.0 -0.1047 0 -2.0 1e-06 
0.0 -0.1046 0 -2.0 1e-06 
0.0 -0.1045 0 -2.0 1e-06 
0.0 -0.1044 0 -2.0 1e-06 
0.0 -0.1043 0 -2.0 1e-06 
0.0 -0.1042 0 -2.0 1e-06 
0.0 -0.1041 0 -2.0 1e-06 
0.0 -0.104 0 -2.0 1e-06 
0.0 -0.1039 0 -2.0 1e-06 
0.0 -0.1038 0 -2.0 1e-06 
0.0 -0.1037 0 -2.0 1e-06 
0.0 -0.1036 0 -2.0 1e-06 
0.0 -0.1035 0 -2.0 1e-06 
0.0 -0.1034 0 -2.0 1e-06 
0.0 -0.1033 0 -2.0 1e-06 
0.0 -0.1032 0 -2.0 1e-06 
0.0 -0.1031 0 -2.0 1e-06 
0.0 -0.103 0 -2.0 1e-06 
0.0 -0.1029 0 -2.0 1e-06 
0.0 -0.1028 0 -2.0 1e-06 
0.0 -0.1027 0 -2.0 1e-06 
0.0 -0.1026 0 -2.0 1e-06 
0.0 -0.1025 0 -2.0 1e-06 
0.0 -0.1024 0 -2.0 1e-06 
0.0 -0.1023 0 -2.0 1e-06 
0.0 -0.1022 0 -2.0 1e-06 
0.0 -0.1021 0 -2.0 1e-06 
0.0 -0.102 0 -2.0 1e-06 
0.0 -0.1019 0 -2.0 1e-06 
0.0 -0.1018 0 -2.0 1e-06 
0.0 -0.1017 0 -2.0 1e-06 
0.0 -0.1016 0 -2.0 1e-06 
0.0 -0.1015 0 -2.0 1e-06 
0.0 -0.1014 0 -2.0 1e-06 
0.0 -0.1013 0 -2.0 1e-06 
0.0 -0.1012 0 -2.0 1e-06 
0.0 -0.1011 0 -2.0 1e-06 
0.0 -0.101 0 -2.0 1e-06 
0.0 -0.1009 0 -2.0 1e-06 
0.0 -0.1008 0 -2.0 1e-06 
0.0 -0.1007 0 -2.0 1e-06 
0.0 -0.1006 0 -2.0 1e-06 
0.0 -0.1005 0 -2.0 1e-06 
0.0 -0.1004 0 -2.0 1e-06 
0.0 -0.1003 0 -2.0 1e-06 
0.0 -0.1002 0 -2.0 1e-06 
0.0 -0.1001 0 -2.0 1e-06 
0.0 -0.1 0 -2.0 1e-06 
0.0 -0.0999000000002 0 -2.0 1e-06 
0.0 -0.0998000000002 0 -2.0 1e-06 
0.0 -0.0997000000002 0 -2.0 1e-06 
0.0 -0.0996000000002 0 -2.0 1e-06 
0.0 -0.0995000000002 0 -2.0 1e-06 
0.0 -0.0994000000002 0 -2.0 1e-06 
0.0 -0.0993000000002 0 -2.0 1e-06 
0.0 -0.0992000000002 0 -2.0 1e-06 
0.0 -0.0991000000002 0 -2.0 1e-06 
0.0 -0.0990000000002 0 -2.0 1e-06 
0.0 -0.0989000000002 0 -2.0 1e-06 
0.0 -0.0988000000002 0 -2.0 1e-06 
0.0 -0.0987000000002 0 -2.0 1e-06 
0.0 -0.0986000000002 0 -2.0 1e-06 
0.0 -0.0985000000002 0 -2.0 1e-06 
0.0 -0.0984000000002 0 -2.0 1e-06 
0.0 -0.0983000000002 0 -2.0 1e-06 
0.0 -0.0982000000002 0 -2.0 1e-06 
0.0 -0.0981000000002 0 -2.0 1e-06 
0.0 -0.0980000000002 0 -2.0 1e-06 
0.0 -0.0979000000002 0 -2.0 1e-06 
0.0 -0.0978000000002 0 -2.0 1e-06 
0.0 -0.0977000000002 0 -2.0 1e-06 
0.0 -0.0976000000002 0 -2.0 1e-06 
0.0 -0.0975000000002 0 -2.0 1e-06 
0.0 -0.0974000000002 0 -2.0 1e-06 
0.0 -0.0973000000002 0 -2.0 1e-06 
0.0 -0.0972000000002 0 -2.0 1e-06 
0.0 -0.0971000000002 0 -2.0 1e-06 
0.0 -0.0970000000002 0 -2.0 1e-06 
0.0 -0.0969000000002 0 -2.0 1e-06 
0.0 -0.0968000000002 0 -2.0 1e-06 
0.0 -0.0967000000002 0 -2.0 1e-06 
0.0 -0.0966000000002 0 -2.0 1e-06 
0.0 -0.0965000000002 0 -2.0 1e-06 
0.0 -0.0964000000002 0 -2.0 1e-06 
0.0 -0.0963000000002 0 -2.0 1e-06 
0.0 -0.0962000000002 0 -2.0 1e-06 
0.0 -0.0961000000002 0 -2.0 1e-06 
0.0 -0.0960000000002 0 -2.0 1e-06 
0.0 -0.0959000000002 0 -2.0 1e-06 
0.0 -0.0958000000002 0 -2.0 1e-06 
0.0 -0.0957000000002 0 -2.0 1e-06 
0.0 -0.0956000000002 0 -2.0 1e-06 
0.0 -0.0955000000002 0 -2.0 1e-06 
0.0 -0.0954000000002 0 -2.0 1e-06 
0.0 -0.0953000000002 0 -2.0 1e-06 
0.0 -0.0952000000002 0 -2.0 1e-06 
0.0 -0.0951000000002 0 -2.0 1e-06 
0.0 -0.0950000000002 0 -2.0 1e-06 
0.0 -0.0949000000002 0 -2.0 1e-06 
0.0 -0.0948000000002 0 -2.0 1e-06 
0.0 -0.0947000000002 0 -2.0 1e-06 
0.0 -0.0946000000002 0 -2.0 1e-06 
0.0 -0.0945000000002 0 -2.0 1e-06 
0.0 -0.0944000000002 0 -2.0 1e-06 
0.0 -0.0943000000002 0 -2.0 1e-06 
0.0 -0.0942000000002 0 -2.0 1e-06 
0.0 -0.0941000000002 0 -2.0 1e-06 
0.0 -0.0940000000002 0 -2.0 1e-06 
0.0 -0.0939000000002 0 -2.0 1e-06 
0.0 -0.0938000000002 0 -2.0 1e-06 
0.0 -0.0937000000002 0 -2.0 1e-06 
0.0 -0.0936000000002 0 -2.0 1e-06 
0.0 -0.0935000000002 0 -2.0 1e-06 
0.0 -0.0934000000002 0 -2.0 1e-06 
0.0 -0.0933000000002 0 -2.0 1e-06 
0.0 -0.0932000000002 0 -2.0 1e-06 
0.0 -0.0931000000002 0 -2.0 1e-06 
0.0 -0.0930000000002 0 -2.0 1e-06 
0.0 -0.0929000000002 0 -2.0 1e-06 
0.0 -0.0928000000002 0 -2.0 1e-06 
0.0 -0.0927000000002 0 -2.0 1e-06 
0.0 -0.0926000000002 0 -2.0 1e-06 
0.0 -0.0925000000002 0 -2.0 1e-06 
0.0 -0.0924000000002 0 -2.0 1e-06 
0.0 -0.0923000000002 0 -2.0 1e-06 
0.0 -0.0922000000002 0 -2.0 1e-06 
0.0 -0.0921000000002 0 -2.0 1e-06 
0.0 -0.0920000000002 0 -2.0 1e-06 
0.0 -0.0919000000002 0 -2.0 1e-06 
0.0 -0.0918000000002 0 -2.0 1e-06 
0.0 -0.0917000000002 0 -2.0 1e-06 
0.0 -0.0916000000002 0 -2.0 1e-06 
0.0 -0.0915000000002 0 -2.0 1e-06 
0.0 -0.0914000000002 0 -2.0 1e-06 
0.0 -0.0913000000002 0 -2.0 1e-06 
0.0 -0.0912000000002 0 -2.0 1e-06 
0.0 -0.0911000000002 0 -2.0 1e-06 
0.0 -0.0910000000002 0 -2.0 1e-06 
0.0 -0.0909000000002 0 -2.0 1e-06 
0.0 -0.0908000000002 0 -2.0 1e-06 
0.0 -0.0907000000002 0 -2.0 1e-06 
0.0 -0.0906000000002 0 -2.0 1e-06 
0.0 -0.0905000000002 0 -2.0 1e-06 
0.0 -0.0904000000002 0 -2.0 1e-06 
0.0 -0.0903000000002 0 -2.0 1e-06 
0.0 -0.0902000000002 0 -2.0 1e-06 
0.0 -0.0901000000002 0 -2.0 1e-06 
0.0 -0.0900000000002 0 -2.0 1e-06 
0.0 -0.0899000000002 0 -2.0 1e-06 
0.0 -0.0898000000002 0 -2.0 1e-06 
0.0 -0.0897000000002 0 -2.0 1e-06 
0.0 -0.0896000000002 0 -2.0 1e-06 
0.0 -0.0895000000002 0 -2.0 1e-06 
0.0 -0.0894000000002 0 -2.0 1e-06 
0.0 -0.0893000000002 0 -2.0 1e-06 
0.0 -0.0892000000002 0 -2.0 1e-06 
0.0 -0.0891000000002 0 -2.0 1e-06 
0.0 -0.0890000000002 0 -2.0 1e-06 
0.0 -0.0889000000002 0 -2.0 1e-06 
0.0 -0.0888000000002 0 -2.0 1e-06 
0.0 -0.0887000000002 0 -2.0 1e-06 
0.0 -0.0886000000002 0 -2.0 1e-06 
0.0 -0.0885000000002 0 -2.0 1e-06 
0.0 -0.0884000000002 0 -2.0 1e-06 
0.0 -0.0883000000002 0 -2.0 1e-06 
0.0 -0.0882000000002 0 -2.0 1e-06 
0.0 -0.0881000000002 0 -2.0 1e-06 
0.0 -0.0880000000002 0 -2.0 1e-06 
0.0 -0.0879000000002 0 -2.0 1e-06 
0.0 -0.0878000000002 0 -2.0 1e-06 
0.0 -0.0877000000002 0 -2.0 1e-06 
0.0 -0.0876000000002 0 -2.0 1e-06 
0.0 -0.0875000000002 0 -2.0 1e-06 
0.0 -0.0874000000002 0 -2.0 1e-06 
0.0 -0.0873000000002 0 -2.0 1e-06 
0.0 -0.0872000000002 0 -2.0 1e-06 
0.0 -0.0871000000002 0 -2.0 1e-06 
0.0 -0.0870000000002 0 -2.0 1e-06 
0.0 -0.0869000000002 0 -2.0 1e-06 
0.0 -0.0868000000002 0 -2.0 1e-06 
0.0 -0.0867000000002 0 -2.0 1e-06 
0.0 -0.0866000000002 0 -2.0 1e-06 
0.0 -0.0865000000002 0 -2.0 1e-06 
0.0 -0.0864000000002 0 -2.0 1e-06 
0.0 -0.0863000000002 0 -2.0 1e-06 
0.0 -0.0862000000002 0 -2.0 1e-06 
0.0 -0.0861000000002 0 -2.0 1e-06 
0.0 -0.0860000000002 0 -2.0 1e-06 
0.0 -0.0859000000002 0 -2.0 1e-06 
0.0 -0.0858000000002 0 -2.0 1e-06 
0.0 -0.0857000000002 0 -2.0 1e-06 
0.0 -0.0856000000002 0 -2.0 1e-06 
0.0 -0.0855000000002 0 -2.0 1e-06 
0.0 -0.0854000000002 0 -2.0 1e-06 
0.0 -0.0853000000002 0 -2.0 1e-06 
0.0 -0.0852000000002 0 -2.0 1e-06 
0.0 -0.0851000000002 0 -2.0 1e-06 
0.0 -0.0850000000002 0 -2.0 1e-06 
0.0 -0.0849000000002 0 -2.0 1e-06 
0.0 -0.0848000000002 0 -2.0 1e-06 
0.0 -0.0847000000002 0 -2.0 1e-06 
0.0 -0.0846000000002 0 -2.0 1e-06 
0.0 -0.0845000000002 0 -2.0 1e-06 
0.0 -0.0844000000002 0 -2.0 1e-06 
0.0 -0.0843000000002 0 -2.0 1e-06 
0.0 -0.0842000000002 0 -2.0 1e-06 
0.0 -0.0841000000002 0 -2.0 1e-06 
0.0 -0.0840000000002 0 -2.0 1e-06 
0.0 -0.0839000000002 0 -2.0 1e-06 
0.0 -0.0838000000002 0 -2.0 1e-06 
0.0 -0.0837000000002 0 -2.0 1e-06 
0.0 -0.0836000000002 0 -2.0 1e-06 
0.0 -0.0835000000002 0 -2.0 1e-06 
0.0 -0.0834000000002 0 -2.0 1e-06 
0.0 -0.0833000000002 0 -2.0 1e-06 
0.0 -0.0832000000002 0 -2.0 1e-06 
0.0 -0.0831000000002 0 -2.0 1e-06 
0.0 -0.0830000000002 0 -2.0 1e-06 
0.0 -0.0829000000002 0 -2.0 1e-06 
0.0 -0.0828000000002 0 -2.0 1e-06 
0.0 -0.0827000000002 0 -2.0 1e-06 
0.0 -0.0826000000002 0 -2.0 1e-06 
0.0 -0.0825000000002 0 -2.0 1e-06 
0.0 -0.0824000000002 0 -2.0 1e-06 
0.0 -0.0823000000002 0 -2.0 1e-06 
0.0 -0.0822000000002 0 -2.0 1e-06 
0.0 -0.0821000000002 0 -2.0 1e-06 
0.0 -0.0820000000002 0 -2.0 1e-06 
0.0 -0.0819000000002 0 -2.0 1e-06 
0.0 -0.0818000000002 0 -2.0 1e-06 
0.0 -0.0817000000002 0 -2.0 1e-06 
0.0 -0.0816000000002 0 -2.0 1e-06 
0.0 -0.0815000000002 0 -2.0 1e-06 
0.0 -0.0814000000002 0 -2.0 1e-06 
0.0 -0.0813000000002 0 -2.0 1e-06 
0.0 -0.0812000000002 0 -2.0 1e-06 
0.0 -0.0811000000002 0 -2.0 1e-06 
0.0 -0.0810000000002 0 -2.0 1e-06 
0.0 -0.0809000000002 0 -2.0 1e-06 
0.0 -0.0808000000002 0 -2.0 1e-06 
0.0 -0.0807000000002 0 -2.0 1e-06 
0.0 -0.0806000000002 0 -2.0 1e-06 
0.0 -0.0805000000002 0 -2.0 1e-06 
0.0 -0.0804000000002 0 -2.0 1e-06 
0.0 -0.0803000000002 0 -2.0 1e-06 
0.0 -0.0802000000002 0 -2.0 1e-06 
0.0 -0.0801000000002 0 -2.0 1e-06 
0.0 -0.0800000000002 0 -2.0 1e-06 
0.0 -0.0799000000002 0 -2.0 1e-06 
0.0 -0.0798000000002 0 -2.0 1e-06 
0.0 -0.0797000000002 0 -2.0 1e-06 
0.0 -0.0796000000002 0 -2.0 1e-06 
0.0 -0.0795000000002 0 -2.0 1e-06 
0.0 -0.0794000000002 0 -2.0 1e-06 
0.0 -0.0793000000002 0 -2.0 1e-06 
0.0 -0.0792000000002 0 -2.0 1e-06 
0.0 -0.0791000000002 0 -2.0 1e-06 
0.0 -0.0790000000002 0 -2.0 1e-06 
0.0 -0.0789000000002 0 -2.0 1e-06 
0.0 -0.0788000000002 0 -2.0 1e-06 
0.0 -0.0787000000002 0 -2.0 1e-06 
0.0 -0.0786000000002 0 -2.0 1e-06 
0.0 -0.0785000000002 0 -2.0 1e-06 
0.0 -0.0784000000002 0 -2.0 1e-06 
0.0 -0.0783000000002 0 -2.0 1e-06 
0.0 -0.0782000000002 0 -2.0 1e-06 
0.0 -0.0781000000002 0 -2.0 1e-06 
0.0 -0.0780000000002 0 -2.0 1e-06 
0.0 -0.0779000000002 0 -2.0 1e-06 
0.0 -0.0778000000002 0 -2.0 1e-06 
0.0 -0.0777000000002 0 -2.0 1e-06 
0.0 -0.0776000000002 0 -2.0 1e-06 
0.0 -0.0775000000002 0 -2.0 1e-06 
0.0 -0.0774000000002 0 -2.0 1e-06 
0.0 -0.0773000000002 0 -2.0 1e-06 
0.0 -0.0772000000002 0 -2.0 1e-06 
0.0 -0.0771000000002 0 -2.0 1e-06 
0.0 -0.0770000000002 0 -2.0 1e-06 
0.0 -0.0769000000002 0 -2.0 1e-06 
0.0 -0.0768000000002 0 -2.0 1e-06 
0.0 -0.0767000000002 0 -2.0 1e-06 
0.0 -0.0766000000002 0 -2.0 1e-06 
0.0 -0.0765000000002 0 -2.0 1e-06 
0.0 -0.0764000000002 0 -2.0 1e-06 
0.0 -0.0763000000002 0 -2.0 1e-06 
0.0 -0.0762000000002 0 -2.0 1e-06 
0.0 -0.0761000000002 0 -2.0 1e-06 
0.0 -0.0760000000002 0 -2.0 1e-06 
0.0 -0.0759000000002 0 -2.0 1e-06 
0.0 -0.0758000000002 0 -2.0 1e-06 
0.0 -0.0757000000002 0 -2.0 1e-06 
0.0 -0.0756000000002 0 -2.0 1e-06 
0.0 -0.0755000000002 0 -2.0 1e-06 
0.0 -0.0754000000002 0 -2.0 1e-06 
0.0 -0.0753000000002 0 -2.0 1e-06 
0.0 -0.0752000000002 0 -2.0 1e-06 
0.0 -0.0751000000002 0 -2.0 1e-06 
0.0 -0.0750000000002 0 -2.0 1e-06 
0.0 -0.0749000000002 0 -2.0 1e-06 
0.0 -0.0748000000002 0 -2.0 1e-06 
0.0 -0.0747000000002 0 -2.0 1e-06 
0.0 -0.0746000000002 0 -2.0 1e-06 
0.0 -0.0745000000002 0 -2.0 1e-06 
0.0 -0.0744000000002 0 -2.0 1e-06 
0.0 -0.0743000000002 0 -2.0 1e-06 
0.0 -0.0742000000002 0 -2.0 1e-06 
0.0 -0.0741000000002 0 -2.0 1e-06 
0.0 -0.0740000000002 0 -2.0 1e-06 
0.0 -0.0739000000002 0 -2.0 1e-06 
0.0 -0.0738000000002 0 -2.0 1e-06 
0.0 -0.0737000000002 0 -2.0 1e-06 
0.0 -0.0736000000002 0 -2.0 1e-06 
0.0 -0.0735000000002 0 -2.0 1e-06 
0.0 -0.0734000000002 0 -2.0 1e-06 
0.0 -0.0733000000002 0 -2.0 1e-06 
0.0 -0.0732000000002 0 -2.0 1e-06 
0.0 -0.0731000000002 0 -2.0 1e-06 
0.0 -0.0730000000002 0 -2.0 1e-06 
0.0 -0.0729000000002 0 -2.0 1e-06 
0.0 -0.0728000000002 0 -2.0 1e-06 
0.0 -0.0727000000002 0 -2.0 1e-06 
0.0 -0.0726000000002 0 -2.0 1e-06 
0.0 -0.0725000000002 0 -2.0 1e-06 
0.0 -0.0724000000002 0 -2.0 1e-06 
0.0 -0.0723000000002 0 -2.0 1e-06 
0.0 -0.0722000000002 0 -2.0 1e-06 
0.0 -0.0721000000002 0 -2.0 1e-06 
0.0 -0.0720000000002 0 -2.0 1e-06 
0.0 -0.0719000000002 0 -2.0 1e-06 
0.0 -0.0718000000002 0 -2.0 1e-06 
0.0 -0.0717000000002 0 -2.0 1e-06 
0.0 -0.0716000000002 0 -2.0 1e-06 
0.0 -0.0715000000002 0 -2.0 1e-06 
0.0 -0.0714000000002 0 -2.0 1e-06 
0.0 -0.0713000000002 0 -2.0 1e-06 
0.0 -0.0712000000002 0 -2.0 1e-06 
0.0 -0.0711000000002 0 -2.0 1e-06 
0.0 -0.0710000000002 0 -2.0 1e-06 
0.0 -0.0709000000002 0 -2.0 1e-06 
0.0 -0.0708000000002 0 -2.0 1e-06 
0.0 -0.0707000000002 0 -2.0 1e-06 
0.0 -0.0706000000002 0 -2.0 1e-06 
0.0 -0.0705000000002 0 -2.0 1e-06 
0.0 -0.0704000000002 0 -2.0 1e-06 
0.0 -0.0703000000002 0 -2.0 1e-06 
0.0 -0.0702000000002 0 -2.0 1e-06 
0.0 -0.0701000000002 0 -2.0 1e-06 
0.0 -0.0700000000002 0 -2.0 1e-06 
0.0 -0.0699000000002 0 -2.0 1e-06 
0.0 -0.0698000000002 0 -2.0 1e-06 
0.0 -0.0697000000002 0 -2.0 1e-06 
0.0 -0.0696000000002 0 -2.0 1e-06 
0.0 -0.0695000000002 0 -2.0 1e-06 
0.0 -0.0694000000002 0 -2.0 1e-06 
0.0 -0.0693000000002 0 -2.0 1e-06 
0.0 -0.0692000000002 0 -2.0 1e-06 
0.0 -0.0691000000002 0 -2.0 1e-06 
0.0 -0.0690000000002 0 -2.0 1e-06 
0.0 -0.0689000000002 0 -2.0 1e-06 
0.0 -0.0688000000002 0 -2.0 1e-06 
0.0 -0.0687000000002 0 -2.0 1e-06 
0.0 -0.0686000000002 0 -2.0 1e-06 
0.0 -0.0685000000002 0 -2.0 1e-06 
0.0 -0.0684000000002 0 -2.0 1e-06 
0.0 -0.0683000000002 0 -2.0 1e-06 
0.0 -0.0682000000002 0 -2.0 1e-06 
0.0 -0.0681000000002 0 -2.0 1e-06 
0.0 -0.0680000000002 0 -2.0 1e-06 
0.0 -0.0679000000002 0 -2.0 1e-06 
0.0 -0.0678000000002 0 -2.0 1e-06 
0.0 -0.0677000000002 0 -2.0 1e-06 
0.0 -0.0676000000002 0 -2.0 1e-06 
0.0 -0.0675000000002 0 -2.0 1e-06 
0.0 -0.0674000000002 0 -2.0 1e-06 
0.0 -0.0673000000002 0 -2.0 1e-06 
0.0 -0.0672000000002 0 -2.0 1e-06 
0.0 -0.0671000000002 0 -2.0 1e-06 
0.0 -0.0670000000002 0 -2.0 1e-06 
0.0 -0.0669000000002 0 -2.0 1e-06 
0.0 -0.0668000000002 0 -2.0 1e-06 
0.0 -0.0667000000002 0 -2.0 1e-06 
0.0 -0.0666000000002 0 -2.0 1e-06 
0.0 -0.0665000000002 0 -2.0 1e-06 
0.0 -0.0664000000002 0 -2.0 1e-06 
0.0 -0.0663000000002 0 -2.0 1e-06 
0.0 -0.0662000000002 0 -2.0 1e-06 
0.0 -0.0661000000002 0 -2.0 1e-06 
0.0 -0.0660000000002 0 -2.0 1e-06 
0.0 -0.0659000000002 0 -2.0 1e-06 
0.0 -0.0658000000002 0 -2.0 1e-06 
0.0 -0.0657000000002 0 -2.0 1e-06 
0.0 -0.0656000000002 0 -2.0 1e-06 
0.0 -0.0655000000002 0 -2.0 1e-06 
0.0 -0.0654000000002 0 -2.0 1e-06 
0.0 -0.0653000000002 0 -2.0 1e-06 
0.0 -0.0652000000002 0 -2.0 1e-06 
0.0 -0.0651000000002 0 -2.0 1e-06 
0.0 -0.0650000000002 0 -2.0 1e-06 
0.0 -0.0649000000002 0 -2.0 1e-06 
0.0 -0.0648000000002 0 -2.0 1e-06 
0.0 -0.0647000000002 0 -2.0 1e-06 
0.0 -0.0646000000002 0 -2.0 1e-06 
0.0 -0.0645000000002 0 -2.0 1e-06 
0.0 -0.0644000000002 0 -2.0 1e-06 
0.0 -0.0643000000002 0 -2.0 1e-06 
0.0 -0.0642000000002 0 -2.0 1e-06 
0.0 -0.0641000000002 0 -2.0 1e-06 
0.0 -0.0640000000002 0 -2.0 1e-06 
0.0 -0.0639000000002 0 -2.0 1e-06 
0.0 -0.0638000000002 0 -2.0 1e-06 
0.0 -0.0637000000002 0 -2.0 1e-06 
0.0 -0.0636000000002 0 -2.0 1e-06 
0.0 -0.0635000000002 0 -2.0 1e-06 
0.0 -0.0634000000002 0 -2.0 1e-06 
0.0 -0.0633000000002 0 -2.0 1e-06 
0.0 -0.0632000000002 0 -2.0 1e-06 
0.0 -0.0631000000002 0 -2.0 1e-06 
0.0 -0.0630000000002 0 -2.0 1e-06 
0.0 -0.0629000000002 0 -2.0 1e-06 
0.0 -0.0628000000002 0 -2.0 1e-06 
0.0 -0.0627000000002 0 -2.0 1e-06 
0.0 -0.0626000000002 0 -2.0 1e-06 
0.0 -0.0625000000002 0 -2.0 1e-06 
0.0 -0.0624000000002 0 -2.0 1e-06 
0.0 -0.0623000000002 0 -2.0 1e-06 
0.0 -0.0622000000002 0 -2.0 1e-06 
0.0 -0.0621000000002 0 -2.0 1e-06 
0.0 -0.0620000000002 0 -2.0 1e-06 
0.0 -0.0619000000002 0 -2.0 1e-06 
0.0 -0.0618000000002 0 -2.0 1e-06 
0.0 -0.0617000000002 0 -2.0 1e-06 
0.0 -0.0616000000002 0 -2.0 1e-06 
0.0 -0.0615000000002 0 -2.0 1e-06 
0.0 -0.0614000000002 0 -2.0 1e-06 
0.0 -0.0613000000002 0 -2.0 1e-06 
0.0 -0.0612000000002 0 -2.0 1e-06 
0.0 -0.0611000000002 0 -2.0 1e-06 
0.0 -0.0610000000002 0 -2.0 1e-06 
0.0 -0.0609000000002 0 -2.0 1e-06 
0.0 -0.0608000000002 0 -2.0 1e-06 
0.0 -0.0607000000002 0 -2.0 1e-06 
0.0 -0.0606000000002 0 -2.0 1e-06 
0.0 -0.0605000000002 0 -2.0 1e-06 
0.0 -0.0604000000002 0 -2.0 1e-06 
0.0 -0.0603000000002 0 -2.0 1e-06 
0.0 -0.0602000000002 0 -2.0 1e-06 
0.0 -0.0601000000002 0 -2.0 1e-06 
0.0 -0.0600000000002 0 -2.0 1e-06 
0.0 -0.0599000000002 0 -2.0 1e-06 
0.0 -0.0598000000002 0 -2.0 1e-06 
0.0 -0.0597000000002 0 -2.0 1e-06 
0.0 -0.0596000000002 0 -2.0 1e-06 
0.0 -0.0595000000002 0 -2.0 1e-06 
0.0 -0.0594000000002 0 -2.0 1e-06 
0.0 -0.0593000000002 0 -2.0 1e-06 
0.0 -0.0592000000002 0 -2.0 1e-06 
0.0 -0.0591000000002 0 -2.0 1e-06 
0.0 -0.0590000000002 0 -2.0 1e-06 
0.0 -0.0589000000002 0 -2.0 1e-06 
0.0 -0.0588000000002 0 -2.0 1e-06 
0.0 -0.0587000000002 0 -2.0 1e-06 
0.0 -0.0586000000002 0 -2.0 1e-06 
0.0 -0.0585000000002 0 -2.0 1e-06 
0.0 -0.0584000000002 0 -2.0 1e-06 
0.0 -0.0583000000002 0 -2.0 1e-06 
0.0 -0.0582000000002 0 -2.0 1e-06 
0.0 -0.0581000000002 0 -2.0 1e-06 
0.0 -0.0580000000002 0 -2.0 1e-06 
0.0 -0.0579000000002 0 -2.0 1e-06 
0.0 -0.0578000000002 0 -2.0 1e-06 
0.0 -0.0577000000002 0 -2.0 1e-06 
0.0 -0.0576000000002 0 -2.0 1e-06 
0.0 -0.0575000000002 0 -2.0 1e-06 
0.0 -0.0574000000002 0 -2.0 1e-06 
0.0 -0.0573000000002 0 -2.0 1e-06 
0.0 -0.0572000000002 0 -2.0 1e-06 
0.0 -0.0571000000002 0 -2.0 1e-06 
0.0 -0.0570000000002 0 -2.0 1e-06 
0.0 -0.0569000000002 0 -2.0 1e-06 
0.0 -0.0568000000002 0 -2.0 1e-06 
0.0 -0.0567000000002 0 -2.0 1e-06 
0.0 -0.0566000000002 0 -2.0 1e-06 
0.0 -0.0565000000002 0 -2.0 1e-06 
0.0 -0.0564000000002 0 -2.0 1e-06 
0.0 -0.0563000000002 0 -2.0 1e-06 
0.0 -0.0562000000002 0 -2.0 1e-06 
0.0 -0.0561000000002 0 -2.0 1e-06 
0.0 -0.0560000000002 0 -2.0 1e-06 
0.0 -0.0559000000002 0 -2.0 1e-06 
0.0 -0.0558000000002 0 -2.0 1e-06 
0.0 -0.0557000000002 0 -2.0 1e-06 
0.0 -0.0556000000002 0 -2.0 1e-06 
0.0 -0.0555000000002 0 -2.0 1e-06 
0.0 -0.0554000000002 0 -2.0 1e-06 
0.0 -0.0553000000002 0 -2.0 1e-06 
0.0 -0.0552000000002 0 -2.0 1e-06 
0.0 -0.0551000000002 0 -2.0 1e-06 
0.0 -0.0550000000002 0 -2.0 1e-06 
0.0 -0.0549000000002 0 -2.0 1e-06 
0.0 -0.0548000000002 0 -2.0 1e-06 
0.0 -0.0547000000002 0 -2.0 1e-06 
0.0 -0.0546000000002 0 -2.0 1e-06 
0.0 -0.0545000000002 0 -2.0 1e-06 
0.0 -0.0544000000002 0 -2.0 1e-06 
0.0 -0.0543000000002 0 -2.0 1e-06 
0.0 -0.0542000000002 0 -2.0 1e-06 
0.0 -0.0541000000002 0 -2.0 1e-06 
0.0 -0.0540000000002 0 -2.0 1e-06 
0.0 -0.0539000000002 0 -2.0 1e-06 
0.0 -0.0538000000002 0 -2.0 1e-06 
0.0 -0.0537000000002 0 -2.0 1e-06 
0.0 -0.0536000000002 0 -2.0 1e-06 
0.0 -0.0535000000002 0 -2.0 1e-06 
0.0 -0.0534000000002 0 -2.0 1e-06 
0.0 -0.0533000000002 0 -2.0 1e-06 
0.0 -0.0532000000002 0 -2.0 1e-06 
0.0 -0.0531000000002 0 -2.0 1e-06 
0.0 -0.0530000000002 0 -2.0 1e-06 
0.0 -0.0529000000002 0 -2.0 1e-06 
0.0 -0.0528000000002 0 -2.0 1e-06 
0.0 -0.0527000000002 0 -2.0 1e-06 
0.0 -0.0526000000002 0 -2.0 1e-06 
0.0 -0.0525000000002 0 -2.0 1e-06 
0.0 -0.0524000000002 0 -2.0 1e-06 
0.0 -0.0523000000002 0 -2.0 1e-06 
0.0 -0.0522000000002 0 -2.0 1e-06 
0.0 -0.0521000000002 0 -2.0 1e-06 
0.0 -0.0520000000002 0 -2.0 1e-06 
0.0 -0.0519000000002 0 -2.0 1e-06 
0.0 -0.0518000000002 0 -2.0 1e-06 
0.0 -0.0517000000002 0 -2.0 1e-06 
0.0 -0.0516000000002 0 -2.0 1e-06 
0.0 -0.0515000000002 0 -2.0 1e-06 
0.0 -0.0514000000002 0 -2.0 1e-06 
0.0 -0.0513000000002 0 -2.0 1e-06 
0.0 -0.0512000000002 0 -2.0 1e-06 
0.0 -0.0511000000002 0 -2.0 1e-06 
0.0 -0.0510000000002 0 -2.0 1e-06 
0.0 -0.0509000000002 0 -2.0 1e-06 
0.0 -0.0508000000002 0 -2.0 1e-06 
0.0 -0.0507000000002 0 -2.0 1e-06 
0.0 -0.0506000000002 0 -2.0 1e-06 
0.0 -0.0505000000002 0 -2.0 1e-06 
0.0 -0.0504000000002 0 -2.0 1e-06 
0.0 -0.0503000000002 0 -2.0 1e-06 
0.0 -0.0502000000002 0 -2.0 1e-06 
0.0 -0.0501000000002 0 -2.0 1e-06 
0.0 -0.0500000000002 0 -2.0 1e-06 
0.0 -0.0499000000002 0 -2.0 1e-06 
0.0 -0.0498000000002 0 -2.0 1e-06 
0.0 -0.0497000000002 0 -2.0 1e-06 
0.0 -0.0496000000002 0 -2.0 1e-06 
0.0 -0.0495000000002 0 -2.0 1e-06 
0.0 -0.0494000000002 0 -2.0 1e-06 
0.0 -0.0493000000002 0 -2.0 1e-06 
0.0 -0.0492000000002 0 -2.0 1e-06 
0.0 -0.0491000000002 0 -2.0 1e-06 
0.0 -0.0490000000002 0 -2.0 1e-06 
0.0 -0.0489000000002 0 -2.0 1e-06 
0.0 -0.0488000000002 0 -2.0 1e-06 
0.0 -0.0487000000002 0 -2.0 1e-06 
0.0 -0.0486000000002 0 -2.0 1e-06 
0.0 -0.0485000000002 0 -2.0 1e-06 
0.0 -0.0484000000002 0 -2.0 1e-06 
0.0 -0.0483000000002 0 -2.0 1e-06 
0.0 -0.0482000000002 0 -2.0 1e-06 
0.0 -0.0481000000002 0 -2.0 1e-06 
0.0 -0.0480000000002 0 -2.0 1e-06 
0.0 -0.0479000000002 0 -2.0 1e-06 
0.0 -0.0478000000002 0 -2.0 1e-06 
0.0 -0.0477000000002 0 -2.0 1e-06 
0.0 -0.0476000000002 0 -2.0 1e-06 
0.0 -0.0475000000002 0 -2.0 1e-06 
0.0 -0.0474000000002 0 -2.0 1e-06 
0.0 -0.0473000000002 0 -2.0 1e-06 
0.0 -0.0472000000002 0 -2.0 1e-06 
0.0 -0.0471000000002 0 -2.0 1e-06 
0.0 -0.0470000000002 0 -2.0 1e-06 
0.0 -0.0469000000002 0 -2.0 1e-06 
0.0 -0.0468000000002 0 -2.0 1e-06 
0.0 -0.0467000000002 0 -2.0 1e-06 
0.0 -0.0466000000002 0 -2.0 1e-06 
0.0 -0.0465000000002 0 -2.0 1e-06 
0.0 -0.0464000000002 0 -2.0 1e-06 
0.0 -0.0463000000002 0 -2.0 1e-06 
0.0 -0.0462000000002 0 -2.0 1e-06 
0.0 -0.0461000000002 0 -2.0 1e-06 
0.0 -0.0460000000002 0 -2.0 1e-06 
0.0 -0.0459000000002 0 -2.0 1e-06 
0.0 -0.0458000000002 0 -2.0 1e-06 
0.0 -0.0457000000002 0 -2.0 1e-06 
0.0 -0.0456000000002 0 -2.0 1e-06 
0.0 -0.0455000000002 0 -2.0 1e-06 
0.0 -0.0454000000002 0 -2.0 1e-06 
0.0 -0.0453000000002 0 -2.0 1e-06 
0.0 -0.0452000000002 0 -2.0 1e-06 
0.0 -0.0451000000002 0 -2.0 1e-06 
0.0 -0.0450000000002 0 -2.0 1e-06 
0.0 -0.0449000000002 0 -2.0 1e-06 
0.0 -0.0448000000002 0 -2.0 1e-06 
0.0 -0.0447000000002 0 -2.0 1e-06 
0.0 -0.0446000000002 0 -2.0 1e-06 
0.0 -0.0445000000002 0 -2.0 1e-06 
0.0 -0.0444000000002 0 -2.0 1e-06 
0.0 -0.0443000000002 0 -2.0 1e-06 
0.0 -0.0442000000002 0 -2.0 1e-06 
0.0 -0.0441000000002 0 -2.0 1e-06 
0.0 -0.0440000000002 0 -2.0 1e-06 
0.0 -0.0439000000002 0 -2.0 1e-06 
0.0 -0.0438000000002 0 -2.0 1e-06 
0.0 -0.0437000000002 0 -2.0 1e-06 
0.0 -0.0436000000002 0 -2.0 1e-06 
0.0 -0.0435000000002 0 -2.0 1e-06 
0.0 -0.0434000000002 0 -2.0 1e-06 
0.0 -0.0433000000002 0 -2.0 1e-06 
0.0 -0.0432000000002 0 -2.0 1e-06 
0.0 -0.0431000000002 0 -2.0 1e-06 
0.0 -0.0430000000002 0 -2.0 1e-06 
0.0 -0.0429000000002 0 -2.0 1e-06 
0.0 -0.0428000000002 0 -2.0 1e-06 
0.0 -0.0427000000002 0 -2.0 1e-06 
0.0 -0.0426000000002 0 -2.0 1e-06 
0.0 -0.0425000000002 0 -2.0 1e-06 
0.0 -0.0424000000002 0 -2.0 1e-06 
0.0 -0.0423000000002 0 -2.0 1e-06 
0.0 -0.0422000000002 0 -2.0 1e-06 
0.0 -0.0421000000002 0 -2.0 1e-06 
0.0 -0.0420000000002 0 -2.0 1e-06 
0.0 -0.0419000000002 0 -2.0 1e-06 
0.0 -0.0418000000002 0 -2.0 1e-06 
0.0 -0.0417000000002 0 -2.0 1e-06 
0.0 -0.0416000000002 0 -2.0 1e-06 
0.0 -0.0415000000002 0 -2.0 1e-06 
0.0 -0.0414000000002 0 -2.0 1e-06 
0.0 -0.0413000000002 0 -2.0 1e-06 
0.0 -0.0412000000002 0 -2.0 1e-06 
0.0 -0.0411000000002 0 -2.0 1e-06 
0.0 -0.0410000000002 0 -2.0 1e-06 
0.0 -0.0409000000002 0 -2.0 1e-06 
0.0 -0.0408000000002 0 -2.0 1e-06 
0.0 -0.0407000000002 0 -2.0 1e-06 
0.0 -0.0406000000002 0 -2.0 1e-06 
0.0 -0.0405000000002 0 -2.0 1e-06 
0.0 -0.0404000000002 0 -2.0 1e-06 
0.0 -0.0403000000002 0 -2.0 1e-06 
0.0 -0.0402000000002 0 -2.0 1e-06 
0.0 -0.0401000000002 0 -2.0 1e-06 
0.0 -0.0400000000002 0 -2.0 1e-06 
0.0 -0.0399000000002 0 -2.0 1e-06 
0.0 -0.0398000000002 0 -2.0 1e-06 
0.0 -0.0397000000002 0 -2.0 1e-06 
0.0 -0.0396000000002 0 -2.0 1e-06 
0.0 -0.0395000000002 0 -2.0 1e-06 
0.0 -0.0394000000002 0 -2.0 1e-06 
0.0 -0.0393000000002 0 -2.0 1e-06 
0.0 -0.0392000000002 0 -2.0 1e-06 
0.0 -0.0391000000002 0 -2.0 1e-06 
0.0 -0.0390000000002 0 -2.0 1e-06 
0.0 -0.0389000000002 0 -2.0 1e-06 
0.0 -0.0388000000002 0 -2.0 1e-06 
0.0 -0.0387000000002 0 -2.0 1e-06 
0.0 -0.0386000000002 0 -2.0 1e-06 
0.0 -0.0385000000002 0 -2.0 1e-06 
0.0 -0.0384000000002 0 -2.0 1e-06 
0.0 -0.0383000000002 0 -2.0 1e-06 
0.0 -0.0382000000002 0 -2.0 1e-06 
0.0 -0.0381000000002 0 -2.0 1e-06 
0.0 -0.0380000000002 0 -2.0 1e-06 
0.0 -0.0379000000002 0 -2.0 1e-06 
0.0 -0.0378000000002 0 -2.0 1e-06 
0.0 -0.0377000000002 0 -2.0 1e-06 
0.0 -0.0376000000002 0 -2.0 1e-06 
0.0 -0.0375000000002 0 -2.0 1e-06 
0.0 -0.0374000000002 0 -2.0 1e-06 
0.0 -0.0373000000002 0 -2.0 1e-06 
0.0 -0.0372000000002 0 -2.0 1e-06 
0.0 -0.0371000000002 0 -2.0 1e-06 
0.0 -0.0370000000002 0 -2.0 1e-06 
0.0 -0.0369000000002 0 -2.0 1e-06 
0.0 -0.0368000000002 0 -2.0 1e-06 
0.0 -0.0367000000002 0 -2.0 1e-06 
0.0 -0.0366000000002 0 -2.0 1e-06 
0.0 -0.0365000000002 0 -2.0 1e-06 
0.0 -0.0364000000002 0 -2.0 1e-06 
0.0 -0.0363000000002 0 -2.0 1e-06 
0.0 -0.0362000000002 0 -2.0 1e-06 
0.0 -0.0361000000002 0 -2.0 1e-06 
0.0 -0.0360000000002 0 -2.0 1e-06 
0.0 -0.0359000000002 0 -2.0 1e-06 
0.0 -0.0358000000002 0 -2.0 1e-06 
0.0 -0.0357000000002 0 -2.0 1e-06 
0.0 -0.0356000000002 0 -2.0 1e-06 
0.0 -0.0355000000002 0 -2.0 1e-06 
0.0 -0.0354000000002 0 -2.0 1e-06 
0.0 -0.0353000000002 0 -2.0 1e-06 
0.0 -0.0352000000002 0 -2.0 1e-06 
0.0 -0.0351000000002 0 -2.0 1e-06 
0.0 -0.0350000000002 0 -2.0 1e-06 
0.0 -0.0349000000002 0 -2.0 1e-06 
0.0 -0.0348000000002 0 -2.0 1e-06 
0.0 -0.0347000000002 0 -2.0 1e-06 
0.0 -0.0346000000002 0 -2.0 1e-06 
0.0 -0.0345000000002 0 -2.0 1e-06 
0.0 -0.0344000000002 0 -2.0 1e-06 
0.0 -0.0343000000002 0 -2.0 1e-06 
0.0 -0.0342000000002 0 -2.0 1e-06 
0.0 -0.0341000000002 0 -2.0 1e-06 
0.0 -0.0340000000002 0 -2.0 1e-06 
0.0 -0.0339000000002 0 -2.0 1e-06 
0.0 -0.0338000000002 0 -2.0 1e-06 
0.0 -0.0337000000002 0 -2.0 1e-06 
0.0 -0.0336000000002 0 -2.0 1e-06 
0.0 -0.0335000000002 0 -2.0 1e-06 
0.0 -0.0334000000002 0 -2.0 1e-06 
0.0 -0.0333000000002 0 -2.0 1e-06 
0.0 -0.0332000000002 0 -2.0 1e-06 
0.0 -0.0331000000002 0 -2.0 1e-06 
0.0 -0.0330000000002 0 -2.0 1e-06 
0.0 -0.0329000000002 0 -2.0 1e-06 
0.0 -0.0328000000002 0 -2.0 1e-06 
0.0 -0.0327000000002 0 -2.0 1e-06 
0.0 -0.0326000000002 0 -2.0 1e-06 
0.0 -0.0325000000002 0 -2.0 1e-06 
0.0 -0.0324000000002 0 -2.0 1e-06 
0.0 -0.0323000000002 0 -2.0 1e-06 
0.0 -0.0322000000002 0 -2.0 1e-06 
0.0 -0.0321000000002 0 -2.0 1e-06 
0.0 -0.0320000000002 0 -2.0 1e-06 
0.0 -0.0319000000002 0 -2.0 1e-06 
0.0 -0.0318000000002 0 -2.0 1e-06 
0.0 -0.0317000000002 0 -2.0 1e-06 
0.0 -0.0316000000002 0 -2.0 1e-06 
0.0 -0.0315000000002 0 -2.0 1e-06 
0.0 -0.0314000000002 0 -2.0 1e-06 
0.0 -0.0313000000002 0 -2.0 1e-06 
0.0 -0.0312000000002 0 -2.0 1e-06 
0.0 -0.0311000000002 0 -2.0 1e-06 
0.0 -0.0310000000002 0 -2.0 1e-06 
0.0 -0.0309000000002 0 -2.0 1e-06 
0.0 -0.0308000000002 0 -2.0 1e-06 
0.0 -0.0307000000002 0 -2.0 1e-06 
0.0 -0.0306000000002 0 -2.0 1e-06 
0.0 -0.0305000000002 0 -2.0 1e-06 
0.0 -0.0304000000002 0 -2.0 1e-06 
0.0 -0.0303000000002 0 -2.0 1e-06 
0.0 -0.0302000000002 0 -2.0 1e-06 
0.0 -0.0301000000002 0 -2.0 1e-06 
0.0 -0.0300000000002 0 -2.0 1e-06 
0.0 -0.0299000000002 0 -2.0 1e-06 
0.0 -0.0298000000002 0 -2.0 1e-06 
0.0 -0.0297000000002 0 -2.0 1e-06 
0.0 -0.0296000000002 0 -2.0 1e-06 
0.0 -0.0295000000002 0 -2.0 1e-06 
0.0 -0.0294000000002 0 -2.0 1e-06 
0.0 -0.0293000000002 0 -2.0 1e-06 
0.0 -0.0292000000002 0 -2.0 1e-06 
0.0 -0.0291000000002 0 -2.0 1e-06 
0.0 -0.0290000000002 0 -2.0 1e-06 
0.0 -0.0289000000002 0 -2.0 1e-06 
0.0 -0.0288000000002 0 -2.0 1e-06 
0.0 -0.0287000000002 0 -2.0 1e-06 
0.0 -0.0286000000002 0 -2.0 1e-06 
0.0 -0.0285000000002 0 -2.0 1e-06 
0.0 -0.0284000000002 0 -2.0 1e-06 
0.0 -0.0283000000002 0 -2.0 1e-06 
0.0 -0.0282000000002 0 -2.0 1e-06 
0.0 -0.0281000000002 0 -2.0 1e-06 
0.0 -0.0280000000002 0 -2.0 1e-06 
0.0 -0.0279000000002 0 -2.0 1e-06 
0.0 -0.0278000000002 0 -2.0 1e-06 
0.0 -0.0277000000002 0 -2.0 1e-06 
0.0 -0.0276000000002 0 -2.0 1e-06 
0.0 -0.0275000000002 0 -2.0 1e-06 
0.0 -0.0274000000002 0 -2.0 1e-06 
0.0 -0.0273000000002 0 -2.0 1e-06 
0.0 -0.0272000000002 0 -2.0 1e-06 
0.0 -0.0271000000002 0 -2.0 1e-06 
0.0 -0.0270000000002 0 -2.0 1e-06 
0.0 -0.0269000000002 0 -2.0 1e-06 
0.0 -0.0268000000002 0 -2.0 1e-06 
0.0 -0.0267000000002 0 -2.0 1e-06 
0.0 -0.0266000000002 0 -2.0 1e-06 
0.0 -0.0265000000002 0 -2.0 1e-06 
0.0 -0.0264000000002 0 -2.0 1e-06 
0.0 -0.0263000000002 0 -2.0 1e-06 
0.0 -0.0262000000002 0 -2.0 1e-06 
0.0 -0.0261000000002 0 -2.0 1e-06 
0.0 -0.0260000000002 0 -2.0 1e-06 
0.0 -0.0259000000002 0 -2.0 1e-06 
0.0 -0.0258000000002 0 -2.0 1e-06 
0.0 -0.0257000000002 0 -2.0 1e-06 
0.0 -0.0256000000002 0 -2.0 1e-06 
0.0 -0.0255000000002 0 -2.0 1e-06 
0.0 -0.0254000000002 0 -2.0 1e-06 
0.0 -0.0253000000002 0 -2.0 1e-06 
0.0 -0.0252000000002 0 -2.0 1e-06 
0.0 -0.0251000000002 0 -2.0 1e-06 
0.0 -0.0250000000002 0 -2.0 1e-06 
0.0 -0.0249000000002 0 -2.0 1e-06 
0.0 -0.0248000000002 0 -2.0 1e-06 
0.0 -0.0247000000002 0 -2.0 1e-06 
0.0 -0.0246000000002 0 -2.0 1e-06 
0.0 -0.0245000000002 0 -2.0 1e-06 
0.0 -0.0244000000002 0 -2.0 1e-06 
0.0 -0.0243000000002 0 -2.0 1e-06 
0.0 -0.0242000000002 0 -2.0 1e-06 
0.0 -0.0241000000002 0 -2.0 1e-06 
0.0 -0.0240000000002 0 -2.0 1e-06 
0.0 -0.0239000000002 0 -2.0 1e-06 
0.0 -0.0238000000002 0 -2.0 1e-06 
0.0 -0.0237000000002 0 -2.0 1e-06 
0.0 -0.0236000000002 0 -2.0 1e-06 
0.0 -0.0235000000002 0 -2.0 1e-06 
0.0 -0.0234000000002 0 -2.0 1e-06 
0.0 -0.0233000000002 0 -2.0 1e-06 
0.0 -0.0232000000002 0 -2.0 1e-06 
0.0 -0.0231000000002 0 -2.0 1e-06 
0.0 -0.0230000000002 0 -2.0 1e-06 
0.0 -0.0229000000002 0 -2.0 1e-06 
0.0 -0.0228000000002 0 -2.0 1e-06 
0.0 -0.0227000000002 0 -2.0 1e-06 
0.0 -0.0226000000002 0 -2.0 1e-06 
0.0 -0.0225000000002 0 -2.0 1e-06 
0.0 -0.0224000000002 0 -2.0 1e-06 
0.0 -0.0223000000002 0 -2.0 1e-06 
0.0 -0.0222000000002 0 -2.0 1e-06 
0.0 -0.0221000000002 0 -2.0 1e-06 
0.0 -0.0220000000002 0 -2.0 1e-06 
0.0 -0.0219000000002 0 -2.0 1e-06 
0.0 -0.0218000000002 0 -2.0 1e-06 
0.0 -0.0217000000002 0 -2.0 1e-06 
0.0 -0.0216000000002 0 -2.0 1e-06 
0.0 -0.0215000000002 0 -2.0 1e-06 
0.0 -0.0214000000002 0 -2.0 1e-06 
0.0 -0.0213000000002 0 -2.0 1e-06 
0.0 -0.0212000000002 0 -2.0 1e-06 
0.0 -0.0211000000002 0 -2.0 1e-06 
0.0 -0.0210000000002 0 -2.0 1e-06 
0.0 -0.0209000000002 0 -2.0 1e-06 
0.0 -0.0208000000002 0 -2.0 1e-06 
0.0 -0.0207000000002 0 -2.0 1e-06 
0.0 -0.0206000000002 0 -2.0 1e-06 
0.0 -0.0205000000002 0 -2.0 1e-06 
0.0 -0.0204000000002 0 -2.0 1e-06 
0.0 -0.0203000000002 0 -2.0 1e-06 
0.0 -0.0202000000002 0 -2.0 1e-06 
0.0 -0.0201000000002 0 -2.0 1e-06 
0.0 -0.0200000000002 0 -2.0 1e-06 
0.0 -0.0199000000002 0 -2.0 1e-06 
0.0 -0.0198000000002 0 -2.0 1e-06 
0.0 -0.0197000000002 0 -2.0 1e-06 
0.0 -0.0196000000002 0 -2.0 1e-06 
0.0 -0.0195000000002 0 -2.0 1e-06 
0.0 -0.0194000000002 0 -2.0 1e-06 
0.0 -0.0193000000002 0 -2.0 1e-06 
0.0 -0.0192000000002 0 -2.0 1e-06 
0.0 -0.0191000000002 0 -2.0 1e-06 
0.0 -0.0190000000002 0 -2.0 1e-06 
0.0 -0.0189000000002 0 -2.0 1e-06 
0.0 -0.0188000000002 0 -2.0 1e-06 
0.0 -0.0187000000002 0 -2.0 1e-06 
0.0 -0.0186000000002 0 -2.0 1e-06 
0.0 -0.0185000000002 0 -2.0 1e-06 
0.0 -0.0184000000002 0 -2.0 1e-06 
0.0 -0.0183000000002 0 -2.0 1e-06 
0.0 -0.0182000000002 0 -2.0 1e-06 
0.0 -0.0181000000002 0 -2.0 1e-06 
0.0 -0.0180000000002 0 -2.0 1e-06 
0.0 -0.0179000000002 0 -2.0 1e-06 
0.0 -0.0178000000002 0 -2.0 1e-06 
0.0 -0.0177000000002 0 -2.0 1e-06 
0.0 -0.0176000000002 0 -2.0 1e-06 
0.0 -0.0175000000002 0 -2.0 1e-06 
0.0 -0.0174000000002 0 -2.0 1e-06 
0.0 -0.0173000000002 0 -2.0 1e-06 
0.0 -0.0172000000002 0 -2.0 1e-06 
0.0 -0.0171000000002 0 -2.0 1e-06 
0.0 -0.0170000000002 0 -2.0 1e-06 
0.0 -0.0169000000002 0 -2.0 1e-06 
0.0 -0.0168000000002 0 -2.0 1e-06 
0.0 -0.0167000000002 0 -2.0 1e-06 
0.0 -0.0166000000002 0 -2.0 1e-06 
0.0 -0.0165000000002 0 -2.0 1e-06 
0.0 -0.0164000000002 0 -2.0 1e-06 
0.0 -0.0163000000002 0 -2.0 1e-06 
0.0 -0.0162000000002 0 -2.0 1e-06 
0.0 -0.0161000000002 0 -2.0 1e-06 
0.0 -0.0160000000002 0 -2.0 1e-06 
0.0 -0.0159000000002 0 -2.0 1e-06 
0.0 -0.0158000000002 0 -2.0 1e-06 
0.0 -0.0157000000002 0 -2.0 1e-06 
0.0 -0.0156000000002 0 -2.0 1e-06 
0.0 -0.0155000000002 0 -2.0 1e-06 
0.0 -0.0154000000002 0 -2.0 1e-06 
0.0 -0.0153000000002 0 -2.0 1e-06 
0.0 -0.0152000000002 0 -2.0 1e-06 
0.0 -0.0151000000002 0 -2.0 1e-06 
0.0 -0.0150000000002 0 -2.0 1e-06 
0.0 -0.0149000000002 0 -2.0 1e-06 
0.0 -0.0148000000002 0 -2.0 1e-06 
0.0 -0.0147000000002 0 -2.0 1e-06 
0.0 -0.0146000000002 0 -2.0 1e-06 
0.0 -0.0145000000002 0 -2.0 1e-06 
0.0 -0.0144000000002 0 -2.0 1e-06 
0.0 -0.0143000000002 0 -2.0 1e-06 
0.0 -0.0142000000002 0 -2.0 1e-06 
0.0 -0.0141000000002 0 -2.0 1e-06 
0.0 -0.0140000000002 0 -2.0 1e-06 
0.0 -0.0139000000002 0 -2.0 1e-06 
0.0 -0.0138000000002 0 -2.0 1e-06 
0.0 -0.0137000000002 0 -2.0 1e-06 
0.0 -0.0136000000002 0 -2.0 1e-06 
0.0 -0.0135000000002 0 -2.0 1e-06 
0.0 -0.0134000000002 0 -2.0 1e-06 
0.0 -0.0133000000002 0 -2.0 1e-06 
0.0 -0.0132000000002 0 -2.0 1e-06 
0.0 -0.0131000000002 0 -2.0 1e-06 
0.0 -0.0130000000002 0 -2.0 1e-06 
0.0 -0.0129000000002 0 -2.0 1e-06 
0.0 -0.0128000000002 0 -2.0 1e-06 
0.0 -0.0127000000002 0 -2.0 1e-06 
0.0 -0.0126000000002 0 -2.0 1e-06 
0.0 -0.0125000000002 0 -2.0 1e-06 
0.0 -0.0124000000002 0 -2.0 1e-06 
0.0 -0.0123000000002 0 -2.0 1e-06 
0.0 -0.0122000000002 0 -2.0 1e-06 
0.0 -0.0121000000002 0 -2.0 1e-06 
0.0 -0.0120000000002 0 -2.0 1e-06 
0.0 -0.0119000000002 0 -2.0 1e-06 
0.0 -0.0118000000002 0 -2.0 1e-06 
0.0 -0.0117000000002 0 -2.0 1e-06 
0.0 -0.0116000000002 0 -2.0 1e-06 
0.0 -0.0115000000002 0 -2.0 1e-06 
0.0 -0.0114000000002 0 -2.0 1e-06 
0.0 -0.0113000000002 0 -2.0 1e-06 
0.0 -0.0112000000002 0 -2.0 1e-06 
0.0 -0.0111000000002 0 -2.0 1e-06 
0.0 -0.0110000000002 0 -2.0 1e-06 
0.0 -0.0109000000002 0 -2.0 1e-06 
0.0 -0.0108000000002 0 -2.0 1e-06 
0.0 -0.0107000000002 0 -2.0 1e-06 
0.0 -0.0106000000002 0 -2.0 1e-06 
0.0 -0.0105000000002 0 -2.0 1e-06 
0.0 -0.0104000000002 0 -2.0 1e-06 
0.0 -0.0103000000002 0 -2.0 1e-06 
0.0 -0.0102000000002 0 -2.0 1e-06 
0.0 -0.0101000000002 0 -2.0 1e-06 
0.0 -0.0100000000002 0 -2.0 1e-06 
0.0 -0.00990000000016 0 -2.0 1e-06 
0.0 -0.00980000000016 0 -2.0 1e-06 
0.0 -0.00970000000016 0 -2.0 1e-06 
0.0 -0.00960000000016 0 -2.0 1e-06 
0.0 -0.00950000000016 0 -2.0 1e-06 
0.0 -0.00940000000016 0 -2.0 1e-06 
0.0 -0.00930000000016 0 -2.0 1e-06 
0.0 -0.00920000000016 0 -2.0 1e-06 
0.0 -0.00910000000016 0 -2.0 1e-06 
0.0 -0.00900000000016 0 -2.0 1e-06 
0.0 -0.00890000000016 0 -2.0 1e-06 
0.0 -0.00880000000016 0 -2.0 1e-06 
0.0 -0.00870000000016 0 -2.0 1e-06 
0.0 -0.00860000000016 0 -2.0 1e-06 
0.0 -0.00850000000016 0 -2.0 1e-06 
0.0 -0.00840000000016 0 -2.0 1e-06 
0.0 -0.00830000000016 0 -2.0 1e-06 
0.0 -0.00820000000016 0 -2.0 1e-06 
0.0 -0.00810000000016 0 -2.0 1e-06 
0.0 -0.00800000000016 0 -2.0 1e-06 
0.0 -0.00790000000016 0 -2.0 1e-06 
0.0 -0.00780000000016 0 -2.0 1e-06 
0.0 -0.00770000000016 0 -2.0 1e-06 
0.0 -0.00760000000016 0 -2.0 1e-06 
0.0 -0.00750000000016 0 -2.0 1e-06 
0.0 -0.00740000000016 0 -2.0 1e-06 
0.0 -0.00730000000016 0 -2.0 1e-06 
0.0 -0.00720000000016 0 -2.0 1e-06 
0.0 -0.00710000000016 0 -2.0 1e-06 
0.0 -0.00700000000016 0 -2.0 1e-06 
0.0 -0.00690000000016 0 -2.0 1e-06 
0.0 -0.00680000000016 0 -2.0 1e-06 
0.0 -0.00670000000016 0 -2.0 1e-06 
0.0 -0.00660000000016 0 -2.0 1e-06 
0.0 -0.00650000000016 0 -2.0 1e-06 
0.0 -0.00640000000016 0 -2.0 1e-06 
0.0 -0.00630000000016 0 -2.0 1e-06 
0.0 -0.00620000000016 0 -2.0 1e-06 
0.0 -0.00610000000016 0 -2.0 1e-06 
0.0 -0.00600000000016 0 -2.0 1e-06 
0.0 -0.00590000000016 0 -2.0 1e-06 
0.0 -0.00580000000016 0 -2.0 1e-06 
0.0 -0.00570000000016 0 -2.0 1e-06 
0.0 -0.00560000000016 0 -2.0 1e-06 
0.0 -0.00550000000016 0 -2.0 1e-06 
0.0 -0.00540000000016 0 -2.0 1e-06 
0.0 -0.00530000000016 0 -2.0 1e-06 
0.0 -0.00520000000016 0 -2.0 1e-06 
0.0 -0.00510000000016 0 -2.0 1e-06 
0.0 -0.00500000000016 0 -2.0 1e-06 
0.0 -0.00490000000016 0 -2.0 1e-06 
0.0 -0.00480000000016 0 -2.0 1e-06 
0.0 -0.00470000000016 0 -2.0 1e-06 
0.0 -0.00460000000016 0 -2.0 1e-06 
0.0 -0.00450000000016 0 -2.0 1e-06 
0.0 -0.00440000000016 0 -2.0 1e-06 
0.0 -0.00430000000016 0 -2.0 1e-06 
0.0 -0.00420000000016 0 -2.0 1e-06 
0.0 -0.00410000000016 0 -2.0 1e-06 
0.0 -0.00400000000016 0 -2.0 1e-06 
0.0 -0.00390000000016 0 -2.0 1e-06 
0.0 -0.00380000000016 0 -2.0 1e-06 
0.0 -0.00370000000016 0 -2.0 1e-06 
0.0 -0.00360000000016 0 -2.0 1e-06 
0.0 -0.00350000000016 0 -2.0 1e-06 
0.0 -0.00340000000016 0 -2.0 1e-06 
0.0 -0.00330000000016 0 -2.0 1e-06 
0.0 -0.00320000000016 0 -2.0 1e-06 
0.0 -0.00310000000016 0 -2.0 1e-06 
0.0 -0.00300000000016 0 -2.0 1e-06 
0.0 -0.00290000000016 0 -2.0 1e-06 
0.0 -0.00280000000016 0 -2.0 1e-06 
0.0 -0.00270000000016 0 -2.0 1e-06 
0.0 -0.00260000000016 0 -2.0 1e-06 
0.0 -0.00250000000016 0 -2.0 1e-06 
0.0 -0.00240000000016 0 -2.0 1e-06 
0.0 -0.00230000000016 0 -2.0 1e-06 
0.0 -0.00220000000016 0 -2.0 1e-06 
0.0 -0.00210000000016 0 -2.0 1e-06 
0.0 -0.00200000000016 0 -2.0 1e-06 
0.0 -0.00190000000016 0 -2.0 1e-06 
0.0 -0.00180000000017 0 -2.0 1e-06 
0.0 -0.00170000000017 0 -2.0 1e-06 
0.0 -0.00160000000017 0 -2.0 1e-06 
0.0 -0.00150000000017 0 -2.0 1e-06 
0.0 -0.00140000000017 0 -2.0 1e-06 
0.0 -0.00130000000017 0 -2.0 1e-06 
0.0 -0.00120000000017 0 -2.0 1e-06 
0.0 -0.00110000000017 0 -2.0 1e-06 
0.0 -0.00100000000017 0 -2.0 1e-06 
0.0 -0.000900000000165 0 -2.0 1e-06 
0.0 -0.000800000000165 0 -2.0 1e-06 
0.0 -0.000700000000165 0 -2.0 1e-06 
0.0 -0.000600000000165 0 -2.0 1e-06 
0.0 -0.000500000000165 0 -2.0 1e-06 
0.0 -0.000400000000165 0 -2.0 1e-06 
0.0 -0.000300000000165 0 -2.0 1e-06 
0.0 -0.000200000000165 0 -2.0 1e-06 
0.0 -0.000100000000165 0 -2.0 1e-06 
0.0 -1.65201186064e-13 0 -2.0 1e-06 
0.0 9.99999998348e-05 0 -2.0 1e-06 
0.0 0.000199999999835 0 -2.0 1e-06 
0.0 0.000299999999835 0 -2.0 1e-06 
0.0 0.000399999999835 0 -2.0 1e-06 
0.0 0.000499999999835 0 -2.0 1e-06 
0.0 0.000599999999835 0 -2.0 1e-06 
0.0 0.000699999999835 0 -2.0 1e-06 
0.0 0.000799999999835 0 -2.0 1e-06 
0.0 0.000899999999835 0 -2.0 1e-06 
0.0 0.000999999999835 0 -2.0 1e-06 
0.0 0.00109999999983 0 -2.0 1e-06 
0.0 0.00119999999983 0 -2.0 1e-06 
0.0 0.00129999999983 0 -2.0 1e-06 
0.0 0.00139999999983 0 -2.0 1e-06 
0.0 0.00149999999983 0 -2.0 1e-06 
0.0 0.00159999999983 0 -2.0 1e-06 
0.0 0.00169999999983 0 -2.0 1e-06 
0.0 0.00179999999983 0 -2.0 1e-06 
0.0 0.00189999999983 0 -2.0 1e-06 
0.0 0.00199999999983 0 -2.0 1e-06 
0.0 0.00209999999983 0 -2.0 1e-06 
0.0 0.00219999999983 0 -2.0 1e-06 
0.0 0.00229999999983 0 -2.0 1e-06 
0.0 0.00239999999983 0 -2.0 1e-06 
0.0 0.00249999999983 0 -2.0 1e-06 
0.0 0.00259999999983 0 -2.0 1e-06 
0.0 0.00269999999983 0 -2.0 1e-06 
0.0 0.00279999999983 0 -2.0 1e-06 
0.0 0.00289999999983 0 -2.0 1e-06 
0.0 0.00299999999983 0 -2.0 1e-06 
0.0 0.00309999999983 0 -2.0 1e-06 
0.0 0.00319999999983 0 -2.0 1e-06 
0.0 0.00329999999983 0 -2.0 1e-06 
0.0 0.00339999999983 0 -2.0 1e-06 
0.0 0.00349999999983 0 -2.0 1e-06 
0.0 0.00359999999983 0 -2.0 1e-06 
0.0 0.00369999999983 0 -2.0 1e-06 
0.0 0.00379999999983 0 -2.0 1e-06 
0.0 0.00389999999983 0 -2.0 1e-06 
0.0 0.00399999999983 0 -2.0 1e-06 
0.0 0.00409999999983 0 -2.0 1e-06 
0.0 0.00419999999983 0 -2.0 1e-06 
0.0 0.00429999999983 0 -2.0 1e-06 
0.0 0.00439999999983 0 -2.0 1e-06 
0.0 0.00449999999983 0 -2.0 1e-06 
0.0 0.00459999999983 0 -2.0 1e-06 
0.0 0.00469999999983 0 -2.0 1e-06 
0.0 0.00479999999983 0 -2.0 1e-06 
0.0 0.00489999999983 0 -2.0 1e-06 
0.0 0.00499999999983 0 -2.0 1e-06 
0.0 0.00509999999983 0 -2.0 1e-06 
0.0 0.00519999999983 0 -2.0 1e-06 
0.0 0.00529999999983 0 -2.0 1e-06 
0.0 0.00539999999983 0 -2.0 1e-06 
0.0 0.00549999999983 0 -2.0 1e-06 
0.0 0.00559999999983 0 -2.0 1e-06 
0.0 0.00569999999983 0 -2.0 1e-06 
0.0 0.00579999999983 0 -2.0 1e-06 
0.0 0.00589999999983 0 -2.0 1e-06 
0.0 0.00599999999983 0 -2.0 1e-06 
0.0 0.00609999999983 0 -2.0 1e-06 
0.0 0.00619999999983 0 -2.0 1e-06 
0.0 0.00629999999983 0 -2.0 1e-06 
0.0 0.00639999999983 0 -2.0 1e-06 
0.0 0.00649999999983 0 -2.0 1e-06 
0.0 0.00659999999983 0 -2.0 1e-06 
0.0 0.00669999999983 0 -2.0 1e-06 
0.0 0.00679999999983 0 -2.0 1e-06 
0.0 0.00689999999983 0 -2.0 1e-06 
0.0 0.00699999999983 0 -2.0 1e-06 
0.0 0.00709999999983 0 -2.0 1e-06 
0.0 0.00719999999983 0 -2.0 1e-06 
0.0 0.00729999999983 0 -2.0 1e-06 
0.0 0.00739999999983 0 -2.0 1e-06 
0.0 0.00749999999983 0 -2.0 1e-06 
0.0 0.00759999999983 0 -2.0 1e-06 
0.0 0.00769999999983 0 -2.0 1e-06 
0.0 0.00779999999983 0 -2.0 1e-06 
0.0 0.00789999999983 0 -2.0 1e-06 
0.0 0.00799999999983 0 -2.0 1e-06 
0.0 0.00809999999983 0 -2.0 1e-06 
0.0 0.00819999999983 0 -2.0 1e-06 
0.0 0.00829999999983 0 -2.0 1e-06 
0.0 0.00839999999983 0 -2.0 1e-06 
0.0 0.00849999999983 0 -2.0 1e-06 
0.0 0.00859999999983 0 -2.0 1e-06 
0.0 0.00869999999983 0 -2.0 1e-06 
0.0 0.00879999999983 0 -2.0 1e-06 
0.0 0.00889999999983 0 -2.0 1e-06 
0.0 0.00899999999983 0 -2.0 1e-06 
0.0 0.00909999999983 0 -2.0 1e-06 
0.0 0.00919999999983 0 -2.0 1e-06 
0.0 0.00929999999983 0 -2.0 1e-06 
0.0 0.00939999999983 0 -2.0 1e-06 
0.0 0.00949999999983 0 -2.0 1e-06 
0.0 0.00959999999983 0 -2.0 1e-06 
0.0 0.00969999999983 0 -2.0 1e-06 
0.0 0.00979999999983 0 -2.0 1e-06 
0.0 0.00989999999983 0 -2.0 1e-06 
0.0 0.00999999999983 0 -2.0 1e-06 
0.0 0.0100999999998 0 -2.0 1e-06 
0.0 0.0101999999998 0 -2.0 1e-06 
0.0 0.0102999999998 0 -2.0 1e-06 
0.0 0.0103999999998 0 -2.0 1e-06 
0.0 0.0104999999998 0 -2.0 1e-06 
0.0 0.0105999999998 0 -2.0 1e-06 
0.0 0.0106999999998 0 -2.0 1e-06 
0.0 0.0107999999998 0 -2.0 1e-06 
0.0 0.0108999999998 0 -2.0 1e-06 
0.0 0.0109999999998 0 -2.0 1e-06 
0.0 0.0110999999998 0 -2.0 1e-06 
0.0 0.0111999999998 0 -2.0 1e-06 
0.0 0.0112999999998 0 -2.0 1e-06 
0.0 0.0113999999998 0 -2.0 1e-06 
0.0 0.0114999999998 0 -2.0 1e-06 
0.0 0.0115999999998 0 -2.0 1e-06 
0.0 0.0116999999998 0 -2.0 1e-06 
0.0 0.0117999999998 0 -2.0 1e-06 
0.0 0.0118999999998 0 -2.0 1e-06 
0.0 0.0119999999998 0 -2.0 1e-06 
0.0 0.0120999999998 0 -2.0 1e-06 
0.0 0.0121999999998 0 -2.0 1e-06 
0.0 0.0122999999998 0 -2.0 1e-06 
0.0 0.0123999999998 0 -2.0 1e-06 
0.0 0.0124999999998 0 -2.0 1e-06 
0.0 0.0125999999998 0 -2.0 1e-06 
0.0 0.0126999999998 0 -2.0 1e-06 
0.0 0.0127999999998 0 -2.0 1e-06 
0.0 0.0128999999998 0 -2.0 1e-06 
0.0 0.0129999999998 0 -2.0 1e-06 
0.0 0.0130999999998 0 -2.0 1e-06 
0.0 0.0131999999998 0 -2.0 1e-06 
0.0 0.0132999999998 0 -2.0 1e-06 
0.0 0.0133999999998 0 -2.0 1e-06 
0.0 0.0134999999998 0 -2.0 1e-06 
0.0 0.0135999999998 0 -2.0 1e-06 
0.0 0.0136999999998 0 -2.0 1e-06 
0.0 0.0137999999998 0 -2.0 1e-06 
0.0 0.0138999999998 0 -2.0 1e-06 
0.0 0.0139999999998 0 -2.0 1e-06 
0.0 0.0140999999998 0 -2.0 1e-06 
0.0 0.0141999999998 0 -2.0 1e-06 
0.0 0.0142999999998 0 -2.0 1e-06 
0.0 0.0143999999998 0 -2.0 1e-06 
0.0 0.0144999999998 0 -2.0 1e-06 
0.0 0.0145999999998 0 -2.0 1e-06 
0.0 0.0146999999998 0 -2.0 1e-06 
0.0 0.0147999999998 0 -2.0 1e-06 
0.0 0.0148999999998 0 -2.0 1e-06 
0.0 0.0149999999998 0 -2.0 1e-06 
0.0 0.0150999999998 0 -2.0 1e-06 
0.0 0.0151999999998 0 -2.0 1e-06 
0.0 0.0152999999998 0 -2.0 1e-06 
0.0 0.0153999999998 0 -2.0 1e-06 
0.0 0.0154999999998 0 -2.0 1e-06 
0.0 0.0155999999998 0 -2.0 1e-06 
0.0 0.0156999999998 0 -2.0 1e-06 
0.0 0.0157999999998 0 -2.0 1e-06 
0.0 0.0158999999998 0 -2.0 1e-06 
0.0 0.0159999999998 0 -2.0 1e-06 
0.0 0.0160999999998 0 -2.0 1e-06 
0.0 0.0161999999998 0 -2.0 1e-06 
0.0 0.0162999999998 0 -2.0 1e-06 
0.0 0.0163999999998 0 -2.0 1e-06 
0.0 0.0164999999998 0 -2.0 1e-06 
0.0 0.0165999999998 0 -2.0 1e-06 
0.0 0.0166999999998 0 -2.0 1e-06 
0.0 0.0167999999998 0 -2.0 1e-06 
0.0 0.0168999999998 0 -2.0 1e-06 
0.0 0.0169999999998 0 -2.0 1e-06 
0.0 0.0170999999998 0 -2.0 1e-06 
0.0 0.0171999999998 0 -2.0 1e-06 
0.0 0.0172999999998 0 -2.0 1e-06 
0.0 0.0173999999998 0 -2.0 1e-06 
0.0 0.0174999999998 0 -2.0 1e-06 
0.0 0.0175999999998 0 -2.0 1e-06 
0.0 0.0176999999998 0 -2.0 1e-06 
0.0 0.0177999999998 0 -2.0 1e-06 
0.0 0.0178999999998 0 -2.0 1e-06 
0.0 0.0179999999998 0 -2.0 1e-06 
0.0 0.0180999999998 0 -2.0 1e-06 
0.0 0.0181999999998 0 -2.0 1e-06 
0.0 0.0182999999998 0 -2.0 1e-06 
0.0 0.0183999999998 0 -2.0 1e-06 
0.0 0.0184999999998 0 -2.0 1e-06 
0.0 0.0185999999998 0 -2.0 1e-06 
0.0 0.0186999999998 0 -2.0 1e-06 
0.0 0.0187999999998 0 -2.0 1e-06 
0.0 0.0188999999998 0 -2.0 1e-06 
0.0 0.0189999999998 0 -2.0 1e-06 
0.0 0.0190999999998 0 -2.0 1e-06 
0.0 0.0191999999998 0 -2.0 1e-06 
0.0 0.0192999999998 0 -2.0 1e-06 
0.0 0.0193999999998 0 -2.0 1e-06 
0.0 0.0194999999998 0 -2.0 1e-06 
0.0 0.0195999999998 0 -2.0 1e-06 
0.0 0.0196999999998 0 -2.0 1e-06 
0.0 0.0197999999998 0 -2.0 1e-06 
0.0 0.0198999999998 0 -2.0 1e-06 
0.0 0.0199999999998 0 -2.0 1e-06 
0.0 0.0200999999998 0 -2.0 1e-06 
0.0 0.0201999999998 0 -2.0 1e-06 
0.0 0.0202999999998 0 -2.0 1e-06 
0.0 0.0203999999998 0 -2.0 1e-06 
0.0 0.0204999999998 0 -2.0 1e-06 
0.0 0.0205999999998 0 -2.0 1e-06 
0.0 0.0206999999998 0 -2.0 1e-06 
0.0 0.0207999999998 0 -2.0 1e-06 
0.0 0.0208999999998 0 -2.0 1e-06 
0.0 0.0209999999998 0 -2.0 1e-06 
0.0 0.0210999999998 0 -2.0 1e-06 
0.0 0.0211999999998 0 -2.0 1e-06 
0.0 0.0212999999998 0 -2.0 1e-06 
0.0 0.0213999999998 0 -2.0 1e-06 
0.0 0.0214999999998 0 -2.0 1e-06 
0.0 0.0215999999998 0 -2.0 1e-06 
0.0 0.0216999999998 0 -2.0 1e-06 
0.0 0.0217999999998 0 -2.0 1e-06 
0.0 0.0218999999998 0 -2.0 1e-06 
0.0 0.0219999999998 0 -2.0 1e-06 
0.0 0.0220999999998 0 -2.0 1e-06 
0.0 0.0221999999998 0 -2.0 1e-06 
0.0 0.0222999999998 0 -2.0 1e-06 
0.0 0.0223999999998 0 -2.0 1e-06 
0.0 0.0224999999998 0 -2.0 1e-06 
0.0 0.0225999999998 0 -2.0 1e-06 
0.0 0.0226999999998 0 -2.0 1e-06 
0.0 0.0227999999998 0 -2.0 1e-06 
0.0 0.0228999999998 0 -2.0 1e-06 
0.0 0.0229999999998 0 -2.0 1e-06 
0.0 0.0230999999998 0 -2.0 1e-06 
0.0 0.0231999999998 0 -2.0 1e-06 
0.0 0.0232999999998 0 -2.0 1e-06 
0.0 0.0233999999998 0 -2.0 1e-06 
0.0 0.0234999999998 0 -2.0 1e-06 
0.0 0.0235999999998 0 -2.0 1e-06 
0.0 0.0236999999998 0 -2.0 1e-06 
0.0 0.0237999999998 0 -2.0 1e-06 
0.0 0.0238999999998 0 -2.0 1e-06 
0.0 0.0239999999998 0 -2.0 1e-06 
0.0 0.0240999999998 0 -2.0 1e-06 
0.0 0.0241999999998 0 -2.0 1e-06 
0.0 0.0242999999998 0 -2.0 1e-06 
0.0 0.0243999999998 0 -2.0 1e-06 
0.0 0.0244999999998 0 -2.0 1e-06 
0.0 0.0245999999998 0 -2.0 1e-06 
0.0 0.0246999999998 0 -2.0 1e-06 
0.0 0.0247999999998 0 -2.0 1e-06 
0.0 0.0248999999998 0 -2.0 1e-06 
0.0 0.0249999999998 0 -2.0 1e-06 
0.0 0.0250999999998 0 -2.0 1e-06 
0.0 0.0251999999998 0 -2.0 1e-06 
0.0 0.0252999999998 0 -2.0 1e-06 
0.0 0.0253999999998 0 -2.0 1e-06 
0.0 0.0254999999998 0 -2.0 1e-06 
0.0 0.0255999999998 0 -2.0 1e-06 
0.0 0.0256999999998 0 -2.0 1e-06 
0.0 0.0257999999998 0 -2.0 1e-06 
0.0 0.0258999999998 0 -2.0 1e-06 
0.0 0.0259999999998 0 -2.0 1e-06 
0.0 0.0260999999998 0 -2.0 1e-06 
0.0 0.0261999999998 0 -2.0 1e-06 
0.0 0.0262999999998 0 -2.0 1e-06 
0.0 0.0263999999998 0 -2.0 1e-06 
0.0 0.0264999999998 0 -2.0 1e-06 
0.0 0.0265999999998 0 -2.0 1e-06 
0.0 0.0266999999998 0 -2.0 1e-06 
0.0 0.0267999999998 0 -2.0 1e-06 
0.0 0.0268999999998 0 -2.0 1e-06 
0.0 0.0269999999998 0 -2.0 1e-06 
0.0 0.0270999999998 0 -2.0 1e-06 
0.0 0.0271999999998 0 -2.0 1e-06 
0.0 0.0272999999998 0 -2.0 1e-06 
0.0 0.0273999999998 0 -2.0 1e-06 
0.0 0.0274999999998 0 -2.0 1e-06 
0.0 0.0275999999998 0 -2.0 1e-06 
0.0 0.0276999999998 0 -2.0 1e-06 
0.0 0.0277999999998 0 -2.0 1e-06 
0.0 0.0278999999998 0 -2.0 1e-06 
0.0 0.0279999999998 0 -2.0 1e-06 
0.0 0.0280999999998 0 -2.0 1e-06 
0.0 0.0281999999998 0 -2.0 1e-06 
0.0 0.0282999999998 0 -2.0 1e-06 
0.0 0.0283999999998 0 -2.0 1e-06 
0.0 0.0284999999998 0 -2.0 1e-06 
0.0 0.0285999999998 0 -2.0 1e-06 
0.0 0.0286999999998 0 -2.0 1e-06 
0.0 0.0287999999998 0 -2.0 1e-06 
0.0 0.0288999999998 0 -2.0 1e-06 
0.0 0.0289999999998 0 -2.0 1e-06 
0.0 0.0290999999998 0 -2.0 1e-06 
0.0 0.0291999999998 0 -2.0 1e-06 
0.0 0.0292999999998 0 -2.0 1e-06 
0.0 0.0293999999998 0 -2.0 1e-06 
0.0 0.0294999999998 0 -2.0 1e-06 
0.0 0.0295999999998 0 -2.0 1e-06 
0.0 0.0296999999998 0 -2.0 1e-06 
0.0 0.0297999999998 0 -2.0 1e-06 
0.0 0.0298999999998 0 -2.0 1e-06 
0.0 0.0299999999998 0 -2.0 1e-06 
0.0 0.0300999999998 0 -2.0 1e-06 
0.0 0.0301999999998 0 -2.0 1e-06 
0.0 0.0302999999998 0 -2.0 1e-06 
0.0 0.0303999999998 0 -2.0 1e-06 
0.0 0.0304999999998 0 -2.0 1e-06 
0.0 0.0305999999998 0 -2.0 1e-06 
0.0 0.0306999999998 0 -2.0 1e-06 
0.0 0.0307999999998 0 -2.0 1e-06 
0.0 0.0308999999998 0 -2.0 1e-06 
0.0 0.0309999999998 0 -2.0 1e-06 
0.0 0.0310999999998 0 -2.0 1e-06 
0.0 0.0311999999998 0 -2.0 1e-06 
0.0 0.0312999999998 0 -2.0 1e-06 
0.0 0.0313999999998 0 -2.0 1e-06 
0.0 0.0314999999998 0 -2.0 1e-06 
0.0 0.0315999999998 0 -2.0 1e-06 
0.0 0.0316999999998 0 -2.0 1e-06 
0.0 0.0317999999998 0 -2.0 1e-06 
0.0 0.0318999999998 0 -2.0 1e-06 
0.0 0.0319999999998 0 -2.0 1e-06 
0.0 0.0320999999998 0 -2.0 1e-06 
0.0 0.0321999999998 0 -2.0 1e-06 
0.0 0.0322999999998 0 -2.0 1e-06 
0.0 0.0323999999998 0 -2.0 1e-06 
0.0 0.0324999999998 0 -2.0 1e-06 
0.0 0.0325999999998 0 -2.0 1e-06 
0.0 0.0326999999998 0 -2.0 1e-06 
0.0 0.0327999999998 0 -2.0 1e-06 
0.0 0.0328999999998 0 -2.0 1e-06 
0.0 0.0329999999998 0 -2.0 1e-06 
0.0 0.0330999999998 0 -2.0 1e-06 
0.0 0.0331999999998 0 -2.0 1e-06 
0.0 0.0332999999998 0 -2.0 1e-06 
0.0 0.0333999999998 0 -2.0 1e-06 
0.0 0.0334999999998 0 -2.0 1e-06 
0.0 0.0335999999998 0 -2.0 1e-06 
0.0 0.0336999999998 0 -2.0 1e-06 
0.0 0.0337999999998 0 -2.0 1e-06 
0.0 0.0338999999998 0 -2.0 1e-06 
0.0 0.0339999999998 0 -2.0 1e-06 
0.0 0.0340999999998 0 -2.0 1e-06 
0.0 0.0341999999998 0 -2.0 1e-06 
0.0 0.0342999999998 0 -2.0 1e-06 
0.0 0.0343999999998 0 -2.0 1e-06 
0.0 0.0344999999998 0 -2.0 1e-06 
0.0 0.0345999999998 0 -2.0 1e-06 
0.0 0.0346999999998 0 -2.0 1e-06 
0.0 0.0347999999998 0 -2.0 1e-06 
0.0 0.0348999999998 0 -2.0 1e-06 
0.0 0.0349999999998 0 -2.0 1e-06 
0.0 0.0350999999998 0 -2.0 1e-06 
0.0 0.0351999999998 0 -2.0 1e-06 
0.0 0.0352999999998 0 -2.0 1e-06 
0.0 0.0353999999998 0 -2.0 1e-06 
0.0 0.0354999999998 0 -2.0 1e-06 
0.0 0.0355999999998 0 -2.0 1e-06 
0.0 0.0356999999998 0 -2.0 1e-06 
0.0 0.0357999999998 0 -2.0 1e-06 
0.0 0.0358999999998 0 -2.0 1e-06 
0.0 0.0359999999998 0 -2.0 1e-06 
0.0 0.0360999999998 0 -2.0 1e-06 
0.0 0.0361999999998 0 -2.0 1e-06 
0.0 0.0362999999998 0 -2.0 1e-06 
0.0 0.0363999999998 0 -2.0 1e-06 
0.0 0.0364999999998 0 -2.0 1e-06 
0.0 0.0365999999998 0 -2.0 1e-06 
0.0 0.0366999999998 0 -2.0 1e-06 
0.0 0.0367999999998 0 -2.0 1e-06 
0.0 0.0368999999998 0 -2.0 1e-06 
0.0 0.0369999999998 0 -2.0 1e-06 
0.0 0.0370999999998 0 -2.0 1e-06 
0.0 0.0371999999998 0 -2.0 1e-06 
0.0 0.0372999999998 0 -2.0 1e-06 
0.0 0.0373999999998 0 -2.0 1e-06 
0.0 0.0374999999998 0 -2.0 1e-06 
0.0 0.0375999999998 0 -2.0 1e-06 
0.0 0.0376999999998 0 -2.0 1e-06 
0.0 0.0377999999998 0 -2.0 1e-06 
0.0 0.0378999999998 0 -2.0 1e-06 
0.0 0.0379999999998 0 -2.0 1e-06 
0.0 0.0380999999998 0 -2.0 1e-06 
0.0 0.0381999999998 0 -2.0 1e-06 
0.0 0.0382999999998 0 -2.0 1e-06 
0.0 0.0383999999998 0 -2.0 1e-06 
0.0 0.0384999999998 0 -2.0 1e-06 
0.0 0.0385999999998 0 -2.0 1e-06 
0.0 0.0386999999998 0 -2.0 1e-06 
0.0 0.0387999999998 0 -2.0 1e-06 
0.0 0.0388999999998 0 -2.0 1e-06 
0.0 0.0389999999998 0 -2.0 1e-06 
0.0 0.0390999999998 0 -2.0 1e-06 
0.0 0.0391999999998 0 -2.0 1e-06 
0.0 0.0392999999998 0 -2.0 1e-06 
0.0 0.0393999999998 0 -2.0 1e-06 
0.0 0.0394999999998 0 -2.0 1e-06 
0.0 0.0395999999998 0 -2.0 1e-06 
0.0 0.0396999999998 0 -2.0 1e-06 
0.0 0.0397999999998 0 -2.0 1e-06 
0.0 0.0398999999998 0 -2.0 1e-06 
0.0 0.0399999999998 0 -2.0 1e-06 
0.0 0.0400999999998 0 -2.0 1e-06 
0.0 0.0401999999998 0 -2.0 1e-06 
0.0 0.0402999999998 0 -2.0 1e-06 
0.0 0.0403999999998 0 -2.0 1e-06 
0.0 0.0404999999998 0 -2.0 1e-06 
0.0 0.0405999999998 0 -2.0 1e-06 
0.0 0.0406999999998 0 -2.0 1e-06 
0.0 0.0407999999998 0 -2.0 1e-06 
0.0 0.0408999999998 0 -2.0 1e-06 
0.0 0.0409999999998 0 -2.0 1e-06 
0.0 0.0410999999998 0 -2.0 1e-06 
0.0 0.0411999999998 0 -2.0 1e-06 
0.0 0.0412999999998 0 -2.0 1e-06 
0.0 0.0413999999998 0 -2.0 1e-06 
0.0 0.0414999999998 0 -2.0 1e-06 
0.0 0.0415999999998 0 -2.0 1e-06 
0.0 0.0416999999998 0 -2.0 1e-06 
0.0 0.0417999999998 0 -2.0 1e-06 
0.0 0.0418999999998 0 -2.0 1e-06 
0.0 0.0419999999998 0 -2.0 1e-06 
0.0 0.0420999999998 0 -2.0 1e-06 
0.0 0.0421999999998 0 -2.0 1e-06 
0.0 0.0422999999998 0 -2.0 1e-06 
0.0 0.0423999999998 0 -2.0 1e-06 
0.0 0.0424999999998 0 -2.0 1e-06 
0.0 0.0425999999998 0 -2.0 1e-06 
0.0 0.0426999999998 0 -2.0 1e-06 
0.0 0.0427999999998 0 -2.0 1e-06 
0.0 0.0428999999998 0 -2.0 1e-06 
0.0 0.0429999999998 0 -2.0 1e-06 
0.0 0.0430999999998 0 -2.0 1e-06 
0.0 0.0431999999998 0 -2.0 1e-06 
0.0 0.0432999999998 0 -2.0 1e-06 
0.0 0.0433999999998 0 -2.0 1e-06 
0.0 0.0434999999998 0 -2.0 1e-06 
0.0 0.0435999999998 0 -2.0 1e-06 
0.0 0.0436999999998 0 -2.0 1e-06 
0.0 0.0437999999998 0 -2.0 1e-06 
0.0 0.0438999999998 0 -2.0 1e-06 
0.0 0.0439999999998 0 -2.0 1e-06 
0.0 0.0440999999998 0 -2.0 1e-06 
0.0 0.0441999999998 0 -2.0 1e-06 
0.0 0.0442999999998 0 -2.0 1e-06 
0.0 0.0443999999998 0 -2.0 1e-06 
0.0 0.0444999999998 0 -2.0 1e-06 
0.0 0.0445999999998 0 -2.0 1e-06 
0.0 0.0446999999998 0 -2.0 1e-06 
0.0 0.0447999999998 0 -2.0 1e-06 
0.0 0.0448999999998 0 -2.0 1e-06 
0.0 0.0449999999998 0 -2.0 1e-06 
0.0 0.0450999999998 0 -2.0 1e-06 
0.0 0.0451999999998 0 -2.0 1e-06 
0.0 0.0452999999998 0 -2.0 1e-06 
0.0 0.0453999999998 0 -2.0 1e-06 
0.0 0.0454999999998 0 -2.0 1e-06 
0.0 0.0455999999998 0 -2.0 1e-06 
0.0 0.0456999999998 0 -2.0 1e-06 
0.0 0.0457999999998 0 -2.0 1e-06 
0.0 0.0458999999998 0 -2.0 1e-06 
0.0 0.0459999999998 0 -2.0 1e-06 
0.0 0.0460999999998 0 -2.0 1e-06 
0.0 0.0461999999998 0 -2.0 1e-06 
0.0 0.0462999999998 0 -2.0 1e-06 
0.0 0.0463999999998 0 -2.0 1e-06 
0.0 0.0464999999998 0 -2.0 1e-06 
0.0 0.0465999999998 0 -2.0 1e-06 
0.0 0.0466999999998 0 -2.0 1e-06 
0.0 0.0467999999998 0 -2.0 1e-06 
0.0 0.0468999999998 0 -2.0 1e-06 
0.0 0.0469999999998 0 -2.0 1e-06 
0.0 0.0470999999998 0 -2.0 1e-06 
0.0 0.0471999999998 0 -2.0 1e-06 
0.0 0.0472999999998 0 -2.0 1e-06 
0.0 0.0473999999998 0 -2.0 1e-06 
0.0 0.0474999999998 0 -2.0 1e-06 
0.0 0.0475999999998 0 -2.0 1e-06 
0.0 0.0476999999998 0 -2.0 1e-06 
0.0 0.0477999999998 0 -2.0 1e-06 
0.0 0.0478999999998 0 -2.0 1e-06 
0.0 0.0479999999998 0 -2.0 1e-06 
0.0 0.0480999999998 0 -2.0 1e-06 
0.0 0.0481999999998 0 -2.0 1e-06 
0.0 0.0482999999998 0 -2.0 1e-06 
0.0 0.0483999999998 0 -2.0 1e-06 
0.0 0.0484999999998 0 -2.0 1e-06 
0.0 0.0485999999998 0 -2.0 1e-06 
0.0 0.0486999999998 0 -2.0 1e-06 
0.0 0.0487999999998 0 -2.0 1e-06 
0.0 0.0488999999998 0 -2.0 1e-06 
0.0 0.0489999999998 0 -2.0 1e-06 
0.0 0.0490999999998 0 -2.0 1e-06 
0.0 0.0491999999998 0 -2.0 1e-06 
0.0 0.0492999999998 0 -2.0 1e-06 
0.0 0.0493999999998 0 -2.0 1e-06 
0.0 0.0494999999998 0 -2.0 1e-06 
0.0 0.0495999999998 0 -2.0 1e-06 
0.0 0.0496999999998 0 -2.0 1e-06 
0.0 0.0497999999998 0 -2.0 1e-06 
0.0 0.0498999999998 0 -2.0 1e-06 
0.0 0.0499999999998 0 -2.0 1e-06 
0.0 0.0500999999998 0 -2.0 1e-06 
0.0 0.0501999999998 0 -2.0 1e-06 
0.0 0.0502999999998 0 -2.0 1e-06 
0.0 0.0503999999998 0 -2.0 1e-06 
0.0 0.0504999999998 0 -2.0 1e-06 
0.0 0.0505999999998 0 -2.0 1e-06 
0.0 0.0506999999998 0 -2.0 1e-06 
0.0 0.0507999999998 0 -2.0 1e-06 
0.0 0.0508999999998 0 -2.0 1e-06 
0.0 0.0509999999998 0 -2.0 1e-06 
0.0 0.0510999999998 0 -2.0 1e-06 
0.0 0.0511999999998 0 -2.0 1e-06 
0.0 0.0512999999998 0 -2.0 1e-06 
0.0 0.0513999999998 0 -2.0 1e-06 
0.0 0.0514999999998 0 -2.0 1e-06 
0.0 0.0515999999998 0 -2.0 1e-06 
0.0 0.0516999999998 0 -2.0 1e-06 
0.0 0.0517999999998 0 -2.0 1e-06 
0.0 0.0518999999998 0 -2.0 1e-06 
0.0 0.0519999999998 0 -2.0 1e-06 
0.0 0.0520999999998 0 -2.0 1e-06 
0.0 0.0521999999998 0 -2.0 1e-06 
0.0 0.0522999999998 0 -2.0 1e-06 
0.0 0.0523999999998 0 -2.0 1e-06 
0.0 0.0524999999998 0 -2.0 1e-06 
0.0 0.0525999999998 0 -2.0 1e-06 
0.0 0.0526999999998 0 -2.0 1e-06 
0.0 0.0527999999998 0 -2.0 1e-06 
0.0 0.0528999999998 0 -2.0 1e-06 
0.0 0.0529999999998 0 -2.0 1e-06 
0.0 0.0530999999998 0 -2.0 1e-06 
0.0 0.0531999999998 0 -2.0 1e-06 
0.0 0.0532999999998 0 -2.0 1e-06 
0.0 0.0533999999998 0 -2.0 1e-06 
0.0 0.0534999999998 0 -2.0 1e-06 
0.0 0.0535999999998 0 -2.0 1e-06 
0.0 0.0536999999998 0 -2.0 1e-06 
0.0 0.0537999999998 0 -2.0 1e-06 
0.0 0.0538999999998 0 -2.0 1e-06 
0.0 0.0539999999998 0 -2.0 1e-06 
0.0 0.0540999999998 0 -2.0 1e-06 
0.0 0.0541999999998 0 -2.0 1e-06 
0.0 0.0542999999998 0 -2.0 1e-06 
0.0 0.0543999999998 0 -2.0 1e-06 
0.0 0.0544999999998 0 -2.0 1e-06 
0.0 0.0545999999998 0 -2.0 1e-06 
0.0 0.0546999999998 0 -2.0 1e-06 
0.0 0.0547999999998 0 -2.0 1e-06 
0.0 0.0548999999998 0 -2.0 1e-06 
0.0 0.0549999999998 0 -2.0 1e-06 
0.0 0.0550999999998 0 -2.0 1e-06 
0.0 0.0551999999998 0 -2.0 1e-06 
0.0 0.0552999999998 0 -2.0 1e-06 
0.0 0.0553999999998 0 -2.0 1e-06 
0.0 0.0554999999998 0 -2.0 1e-06 
0.0 0.0555999999998 0 -2.0 1e-06 
0.0 0.0556999999998 0 -2.0 1e-06 
0.0 0.0557999999998 0 -2.0 1e-06 
0.0 0.0558999999998 0 -2.0 1e-06 
0.0 0.0559999999998 0 -2.0 1e-06 
0.0 0.0560999999998 0 -2.0 1e-06 
0.0 0.0561999999998 0 -2.0 1e-06 
0.0 0.0562999999998 0 -2.0 1e-06 
0.0 0.0563999999998 0 -2.0 1e-06 
0.0 0.0564999999998 0 -2.0 1e-06 
0.0 0.0565999999998 0 -2.0 1e-06 
0.0 0.0566999999998 0 -2.0 1e-06 
0.0 0.0567999999998 0 -2.0 1e-06 
0.0 0.0568999999998 0 -2.0 1e-06 
0.0 0.0569999999998 0 -2.0 1e-06 
0.0 0.0570999999998 0 -2.0 1e-06 
0.0 0.0571999999998 0 -2.0 1e-06 
0.0 0.0572999999998 0 -2.0 1e-06 
0.0 0.0573999999998 0 -2.0 1e-06 
0.0 0.0574999999998 0 -2.0 1e-06 
0.0 0.0575999999998 0 -2.0 1e-06 
0.0 0.0576999999998 0 -2.0 1e-06 
0.0 0.0577999999998 0 -2.0 1e-06 
0.0 0.0578999999998 0 -2.0 1e-06 
0.0 0.0579999999998 0 -2.0 1e-06 
0.0 0.0580999999998 0 -2.0 1e-06 
0.0 0.0581999999998 0 -2.0 1e-06 
0.0 0.0582999999998 0 -2.0 1e-06 
0.0 0.0583999999998 0 -2.0 1e-06 
0.0 0.0584999999998 0 -2.0 1e-06 
0.0 0.0585999999998 0 -2.0 1e-06 
0.0 0.0586999999998 0 -2.0 1e-06 
0.0 0.0587999999998 0 -2.0 1e-06 
0.0 0.0588999999998 0 -2.0 1e-06 
0.0 0.0589999999998 0 -2.0 1e-06 
0.0 0.0590999999998 0 -2.0 1e-06 
0.0 0.0591999999998 0 -2.0 1e-06 
0.0 0.0592999999998 0 -2.0 1e-06 
0.0 0.0593999999998 0 -2.0 1e-06 
0.0 0.0594999999998 0 -2.0 1e-06 
0.0 0.0595999999998 0 -2.0 1e-06 
0.0 0.0596999999998 0 -2.0 1e-06 
0.0 0.0597999999998 0 -2.0 1e-06 
0.0 0.0598999999998 0 -2.0 1e-06 
0.0 0.0599999999998 0 -2.0 1e-06 
0.0 0.0600999999998 0 -2.0 1e-06 
0.0 0.0601999999998 0 -2.0 1e-06 
0.0 0.0602999999998 0 -2.0 1e-06 
0.0 0.0603999999998 0 -2.0 1e-06 
0.0 0.0604999999998 0 -2.0 1e-06 
0.0 0.0605999999998 0 -2.0 1e-06 
0.0 0.0606999999998 0 -2.0 1e-06 
0.0 0.0607999999998 0 -2.0 1e-06 
0.0 0.0608999999998 0 -2.0 1e-06 
0.0 0.0609999999998 0 -2.0 1e-06 
0.0 0.0610999999998 0 -2.0 1e-06 
0.0 0.0611999999998 0 -2.0 1e-06 
0.0 0.0612999999998 0 -2.0 1e-06 
0.0 0.0613999999998 0 -2.0 1e-06 
0.0 0.0614999999998 0 -2.0 1e-06 
0.0 0.0615999999998 0 -2.0 1e-06 
0.0 0.0616999999998 0 -2.0 1e-06 
0.0 0.0617999999998 0 -2.0 1e-06 
0.0 0.0618999999998 0 -2.0 1e-06 
0.0 0.0619999999998 0 -2.0 1e-06 
0.0 0.0620999999998 0 -2.0 1e-06 
0.0 0.0621999999998 0 -2.0 1e-06 
0.0 0.0622999999998 0 -2.0 1e-06 
0.0 0.0623999999998 0 -2.0 1e-06 
0.0 0.0624999999998 0 -2.0 1e-06 
0.0 0.0625999999998 0 -2.0 1e-06 
0.0 0.0626999999998 0 -2.0 1e-06 
0.0 0.0627999999998 0 -2.0 1e-06 
0.0 0.0628999999998 0 -2.0 1e-06 
0.0 0.0629999999998 0 -2.0 1e-06 
0.0 0.0630999999998 0 -2.0 1e-06 
0.0 0.0631999999998 0 -2.0 1e-06 
0.0 0.0632999999998 0 -2.0 1e-06 
0.0 0.0633999999998 0 -2.0 1e-06 
0.0 0.0634999999998 0 -2.0 1e-06 
0.0 0.0635999999998 0 -2.0 1e-06 
0.0 0.0636999999998 0 -2.0 1e-06 
0.0 0.0637999999998 0 -2.0 1e-06 
0.0 0.0638999999998 0 -2.0 1e-06 
0.0 0.0639999999998 0 -2.0 1e-06 
0.0 0.0640999999998 0 -2.0 1e-06 
0.0 0.0641999999998 0 -2.0 1e-06 
0.0 0.0642999999998 0 -2.0 1e-06 
0.0 0.0643999999998 0 -2.0 1e-06 
0.0 0.0644999999998 0 -2.0 1e-06 
0.0 0.0645999999998 0 -2.0 1e-06 
0.0 0.0646999999998 0 -2.0 1e-06 
0.0 0.0647999999998 0 -2.0 1e-06 
0.0 0.0648999999998 0 -2.0 1e-06 
0.0 0.0649999999998 0 -2.0 1e-06 
0.0 0.0650999999998 0 -2.0 1e-06 
0.0 0.0651999999998 0 -2.0 1e-06 
0.0 0.0652999999998 0 -2.0 1e-06 
0.0 0.0653999999998 0 -2.0 1e-06 
0.0 0.0654999999998 0 -2.0 1e-06 
0.0 0.0655999999998 0 -2.0 1e-06 
0.0 0.0656999999998 0 -2.0 1e-06 
0.0 0.0657999999998 0 -2.0 1e-06 
0.0 0.0658999999998 0 -2.0 1e-06 
0.0 0.0659999999998 0 -2.0 1e-06 
0.0 0.0660999999998 0 -2.0 1e-06 
0.0 0.0661999999998 0 -2.0 1e-06 
0.0 0.0662999999998 0 -2.0 1e-06 
0.0 0.0663999999998 0 -2.0 1e-06 
0.0 0.0664999999998 0 -2.0 1e-06 
0.0 0.0665999999998 0 -2.0 1e-06 
0.0 0.0666999999998 0 -2.0 1e-06 
0.0 0.0667999999998 0 -2.0 1e-06 
0.0 0.0668999999998 0 -2.0 1e-06 
0.0 0.0669999999998 0 -2.0 1e-06 
0.0 0.0670999999998 0 -2.0 1e-06 
0.0 0.0671999999998 0 -2.0 1e-06 
0.0 0.0672999999998 0 -2.0 1e-06 
0.0 0.0673999999998 0 -2.0 1e-06 
0.0 0.0674999999998 0 -2.0 1e-06 
0.0 0.0675999999998 0 -2.0 1e-06 
0.0 0.0676999999998 0 -2.0 1e-06 
0.0 0.0677999999998 0 -2.0 1e-06 
0.0 0.0678999999998 0 -2.0 1e-06 
0.0 0.0679999999998 0 -2.0 1e-06 
0.0 0.0680999999998 0 -2.0 1e-06 
0.0 0.0681999999998 0 -2.0 1e-06 
0.0 0.0682999999998 0 -2.0 1e-06 
0.0 0.0683999999998 0 -2.0 1e-06 
0.0 0.0684999999998 0 -2.0 1e-06 
0.0 0.0685999999998 0 -2.0 1e-06 
0.0 0.0686999999998 0 -2.0 1e-06 
0.0 0.0687999999998 0 -2.0 1e-06 
0.0 0.0688999999998 0 -2.0 1e-06 
0.0 0.0689999999998 0 -2.0 1e-06 
0.0 0.0690999999998 0 -2.0 1e-06 
0.0 0.0691999999998 0 -2.0 1e-06 
0.0 0.0692999999998 0 -2.0 1e-06 
0.0 0.0693999999998 0 -2.0 1e-06 
0.0 0.0694999999998 0 -2.0 1e-06 
0.0 0.0695999999998 0 -2.0 1e-06 
0.0 0.0696999999998 0 -2.0 1e-06 
0.0 0.0697999999998 0 -2.0 1e-06 
0.0 0.0698999999998 0 -2.0 1e-06 
0.0 0.0699999999998 0 -2.0 1e-06 
0.0 0.0700999999998 0 -2.0 1e-06 
0.0 0.0701999999998 0 -2.0 1e-06 
0.0 0.0702999999998 0 -2.0 1e-06 
0.0 0.0703999999998 0 -2.0 1e-06 
0.0 0.0704999999998 0 -2.0 1e-06 
0.0 0.0705999999998 0 -2.0 1e-06 
0.0 0.0706999999998 0 -2.0 1e-06 
0.0 0.0707999999998 0 -2.0 1e-06 
0.0 0.0708999999998 0 -2.0 1e-06 
0.0 0.0709999999998 0 -2.0 1e-06 
0.0 0.0710999999998 0 -2.0 1e-06 
0.0 0.0711999999998 0 -2.0 1e-06 
0.0 0.0712999999998 0 -2.0 1e-06 
0.0 0.0713999999998 0 -2.0 1e-06 
0.0 0.0714999999998 0 -2.0 1e-06 
0.0 0.0715999999998 0 -2.0 1e-06 
0.0 0.0716999999998 0 -2.0 1e-06 
0.0 0.0717999999998 0 -2.0 1e-06 
0.0 0.0718999999998 0 -2.0 1e-06 
0.0 0.0719999999998 0 -2.0 1e-06 
0.0 0.0720999999998 0 -2.0 1e-06 
0.0 0.0721999999998 0 -2.0 1e-06 
0.0 0.0722999999998 0 -2.0 1e-06 
0.0 0.0723999999998 0 -2.0 1e-06 
0.0 0.0724999999998 0 -2.0 1e-06 
0.0 0.0725999999998 0 -2.0 1e-06 
0.0 0.0726999999998 0 -2.0 1e-06 
0.0 0.0727999999998 0 -2.0 1e-06 
0.0 0.0728999999998 0 -2.0 1e-06 
0.0 0.0729999999998 0 -2.0 1e-06 
0.0 0.0730999999998 0 -2.0 1e-06 
0.0 0.0731999999998 0 -2.0 1e-06 
0.0 0.0732999999998 0 -2.0 1e-06 
0.0 0.0733999999998 0 -2.0 1e-06 
0.0 0.0734999999998 0 -2.0 1e-06 
0.0 0.0735999999998 0 -2.0 1e-06 
0.0 0.0736999999998 0 -2.0 1e-06 
0.0 0.0737999999998 0 -2.0 1e-06 
0.0 0.0738999999998 0 -2.0 1e-06 
0.0 0.0739999999998 0 -2.0 1e-06 
0.0 0.0740999999998 0 -2.0 1e-06 
0.0 0.0741999999998 0 -2.0 1e-06 
0.0 0.0742999999998 0 -2.0 1e-06 
0.0 0.0743999999998 0 -2.0 1e-06 
0.0 0.0744999999998 0 -2.0 1e-06 
0.0 0.0745999999998 0 -2.0 1e-06 
0.0 0.0746999999998 0 -2.0 1e-06 
0.0 0.0747999999998 0 -2.0 1e-06 
0.0 0.0748999999998 0 -2.0 1e-06 
0.0 0.0749999999998 0 -2.0 1e-06 
0.0 0.0750999999998 0 -2.0 1e-06 
0.0 0.0751999999998 0 -2.0 1e-06 
0.0 0.0752999999998 0 -2.0 1e-06 
0.0 0.0753999999998 0 -2.0 1e-06 
0.0 0.0754999999998 0 -2.0 1e-06 
0.0 0.0755999999998 0 -2.0 1e-06 
0.0 0.0756999999998 0 -2.0 1e-06 
0.0 0.0757999999998 0 -2.0 1e-06 
0.0 0.0758999999998 0 -2.0 1e-06 
0.0 0.0759999999998 0 -2.0 1e-06 
0.0 0.0760999999998 0 -2.0 1e-06 
0.0 0.0761999999998 0 -2.0 1e-06 
0.0 0.0762999999998 0 -2.0 1e-06 
0.0 0.0763999999998 0 -2.0 1e-06 
0.0 0.0764999999998 0 -2.0 1e-06 
0.0 0.0765999999998 0 -2.0 1e-06 
0.0 0.0766999999998 0 -2.0 1e-06 
0.0 0.0767999999998 0 -2.0 1e-06 
0.0 0.0768999999998 0 -2.0 1e-06 
0.0 0.0769999999998 0 -2.0 1e-06 
0.0 0.0770999999998 0 -2.0 1e-06 
0.0 0.0771999999998 0 -2.0 1e-06 
0.0 0.0772999999998 0 -2.0 1e-06 
0.0 0.0773999999998 0 -2.0 1e-06 
0.0 0.0774999999998 0 -2.0 1e-06 
0.0 0.0775999999998 0 -2.0 1e-06 
0.0 0.0776999999998 0 -2.0 1e-06 
0.0 0.0777999999998 0 -2.0 1e-06 
0.0 0.0778999999998 0 -2.0 1e-06 
0.0 0.0779999999998 0 -2.0 1e-06 
0.0 0.0780999999998 0 -2.0 1e-06 
0.0 0.0781999999998 0 -2.0 1e-06 
0.0 0.0782999999998 0 -2.0 1e-06 
0.0 0.0783999999998 0 -2.0 1e-06 
0.0 0.0784999999998 0 -2.0 1e-06 
0.0 0.0785999999998 0 -2.0 1e-06 
0.0 0.0786999999998 0 -2.0 1e-06 
0.0 0.0787999999998 0 -2.0 1e-06 
0.0 0.0788999999998 0 -2.0 1e-06 
0.0 0.0789999999998 0 -2.0 1e-06 
0.0 0.0790999999998 0 -2.0 1e-06 
0.0 0.0791999999998 0 -2.0 1e-06 
0.0 0.0792999999998 0 -2.0 1e-06 
0.0 0.0793999999998 0 -2.0 1e-06 
0.0 0.0794999999998 0 -2.0 1e-06 
0.0 0.0795999999998 0 -2.0 1e-06 
0.0 0.0796999999998 0 -2.0 1e-06 
0.0 0.0797999999998 0 -2.0 1e-06 
0.0 0.0798999999998 0 -2.0 1e-06 
0.0 0.0799999999998 0 -2.0 1e-06 
0.0 0.0800999999998 0 -2.0 1e-06 
0.0 0.0801999999998 0 -2.0 1e-06 
0.0 0.0802999999998 0 -2.0 1e-06 
0.0 0.0803999999998 0 -2.0 1e-06 
0.0 0.0804999999998 0 -2.0 1e-06 
0.0 0.0805999999998 0 -2.0 1e-06 
0.0 0.0806999999998 0 -2.0 1e-06 
0.0 0.0807999999998 0 -2.0 1e-06 
0.0 0.0808999999998 0 -2.0 1e-06 
0.0 0.0809999999998 0 -2.0 1e-06 
0.0 0.0810999999998 0 -2.0 1e-06 
0.0 0.0811999999998 0 -2.0 1e-06 
0.0 0.0812999999998 0 -2.0 1e-06 
0.0 0.0813999999998 0 -2.0 1e-06 
0.0 0.0814999999998 0 -2.0 1e-06 
0.0 0.0815999999998 0 -2.0 1e-06 
0.0 0.0816999999998 0 -2.0 1e-06 
0.0 0.0817999999998 0 -2.0 1e-06 
0.0 0.0818999999998 0 -2.0 1e-06 
0.0 0.0819999999998 0 -2.0 1e-06 
0.0 0.0820999999998 0 -2.0 1e-06 
0.0 0.0821999999998 0 -2.0 1e-06 
0.0 0.0822999999998 0 -2.0 1e-06 
0.0 0.0823999999998 0 -2.0 1e-06 
0.0 0.0824999999998 0 -2.0 1e-06 
0.0 0.0825999999998 0 -2.0 1e-06 
0.0 0.0826999999998 0 -2.0 1e-06 
0.0 0.0827999999998 0 -2.0 1e-06 
0.0 0.0828999999998 0 -2.0 1e-06 
0.0 0.0829999999998 0 -2.0 1e-06 
0.0 0.0830999999998 0 -2.0 1e-06 
0.0 0.0831999999998 0 -2.0 1e-06 
0.0 0.0832999999998 0 -2.0 1e-06 
0.0 0.0833999999998 0 -2.0 1e-06 
0.0 0.0834999999998 0 -2.0 1e-06 
0.0 0.0835999999998 0 -2.0 1e-06 
0.0 0.0836999999998 0 -2.0 1e-06 
0.0 0.0837999999998 0 -2.0 1e-06 
0.0 0.0838999999998 0 -2.0 1e-06 
0.0 0.0839999999998 0 -2.0 1e-06 
0.0 0.0840999999998 0 -2.0 1e-06 
0.0 0.0841999999998 0 -2.0 1e-06 
0.0 0.0842999999998 0 -2.0 1e-06 
0.0 0.0843999999998 0 -2.0 1e-06 
0.0 0.0844999999998 0 -2.0 1e-06 
0.0 0.0845999999998 0 -2.0 1e-06 
0.0 0.0846999999998 0 -2.0 1e-06 
0.0 0.0847999999998 0 -2.0 1e-06 
0.0 0.0848999999998 0 -2.0 1e-06 
0.0 0.0849999999998 0 -2.0 1e-06 
0.0 0.0850999999998 0 -2.0 1e-06 
0.0 0.0851999999998 0 -2.0 1e-06 
0.0 0.0852999999998 0 -2.0 1e-06 
0.0 0.0853999999998 0 -2.0 1e-06 
0.0 0.0854999999998 0 -2.0 1e-06 
0.0 0.0855999999998 0 -2.0 1e-06 
0.0 0.0856999999998 0 -2.0 1e-06 
0.0 0.0857999999998 0 -2.0 1e-06 
0.0 0.0858999999998 0 -2.0 1e-06 
0.0 0.0859999999998 0 -2.0 1e-06 
0.0 0.0860999999998 0 -2.0 1e-06 
0.0 0.0861999999998 0 -2.0 1e-06 
0.0 0.0862999999998 0 -2.0 1e-06 
0.0 0.0863999999998 0 -2.0 1e-06 
0.0 0.0864999999998 0 -2.0 1e-06 
0.0 0.0865999999998 0 -2.0 1e-06 
0.0 0.0866999999998 0 -2.0 1e-06 
0.0 0.0867999999998 0 -2.0 1e-06 
0.0 0.0868999999998 0 -2.0 1e-06 
0.0 0.0869999999998 0 -2.0 1e-06 
0.0 0.0870999999998 0 -2.0 1e-06 
0.0 0.0871999999998 0 -2.0 1e-06 
0.0 0.0872999999998 0 -2.0 1e-06 
0.0 0.0873999999998 0 -2.0 1e-06 
0.0 0.0874999999998 0 -2.0 1e-06 
0.0 0.0875999999998 0 -2.0 1e-06 
0.0 0.0876999999998 0 -2.0 1e-06 
0.0 0.0877999999998 0 -2.0 1e-06 
0.0 0.0878999999998 0 -2.0 1e-06 
0.0 0.0879999999998 0 -2.0 1e-06 
0.0 0.0880999999998 0 -2.0 1e-06 
0.0 0.0881999999998 0 -2.0 1e-06 
0.0 0.0882999999998 0 -2.0 1e-06 
0.0 0.0883999999998 0 -2.0 1e-06 
0.0 0.0884999999998 0 -2.0 1e-06 
0.0 0.0885999999998 0 -2.0 1e-06 
0.0 0.0886999999998 0 -2.0 1e-06 
0.0 0.0887999999998 0 -2.0 1e-06 
0.0 0.0888999999998 0 -2.0 1e-06 
0.0 0.0889999999998 0 -2.0 1e-06 
0.0 0.0890999999998 0 -2.0 1e-06 
0.0 0.0891999999998 0 -2.0 1e-06 
0.0 0.0892999999998 0 -2.0 1e-06 
0.0 0.0893999999998 0 -2.0 1e-06 
0.0 0.0894999999998 0 -2.0 1e-06 
0.0 0.0895999999998 0 -2.0 1e-06 
0.0 0.0896999999998 0 -2.0 1e-06 
0.0 0.0897999999998 0 -2.0 1e-06 
0.0 0.0898999999998 0 -2.0 1e-06 
0.0 0.0899999999998 0 -2.0 1e-06 
0.0 0.0900999999998 0 -2.0 1e-06 
0.0 0.0901999999998 0 -2.0 1e-06 
0.0 0.0902999999998 0 -2.0 1e-06 
0.0 0.0903999999998 0 -2.0 1e-06 
0.0 0.0904999999998 0 -2.0 1e-06 
0.0 0.0905999999998 0 -2.0 1e-06 
0.0 0.0906999999998 0 -2.0 1e-06 
0.0 0.0907999999998 0 -2.0 1e-06 
0.0 0.0908999999998 0 -2.0 1e-06 
0.0 0.0909999999998 0 -2.0 1e-06 
0.0 0.0910999999998 0 -2.0 1e-06 
0.0 0.0911999999998 0 -2.0 1e-06 
0.0 0.0912999999998 0 -2.0 1e-06 
0.0 0.0913999999998 0 -2.0 1e-06 
0.0 0.0914999999998 0 -2.0 1e-06 
0.0 0.0915999999998 0 -2.0 1e-06 
0.0 0.0916999999998 0 -2.0 1e-06 
0.0 0.0917999999998 0 -2.0 1e-06 
0.0 0.0918999999998 0 -2.0 1e-06 
0.0 0.0919999999998 0 -2.0 1e-06 
0.0 0.0920999999998 0 -2.0 1e-06 
0.0 0.0921999999998 0 -2.0 1e-06 
0.0 0.0922999999998 0 -2.0 1e-06 
0.0 0.0923999999998 0 -2.0 1e-06 
0.0 0.0924999999998 0 -2.0 1e-06 
0.0 0.0925999999998 0 -2.0 1e-06 
0.0 0.0926999999998 0 -2.0 1e-06 
0.0 0.0927999999998 0 -2.0 1e-06 
0.0 0.0928999999998 0 -2.0 1e-06 
0.0 0.0929999999998 0 -2.0 1e-06 
0.0 0.0930999999998 0 -2.0 1e-06 
0.0 0.0931999999998 0 -2.0 1e-06 
0.0 0.0932999999998 0 -2.0 1e-06 
0.0 0.0933999999998 0 -2.0 1e-06 
0.0 0.0934999999998 0 -2.0 1e-06 
0.0 0.0935999999998 0 -2.0 1e-06 
0.0 0.0936999999998 0 -2.0 1e-06 
0.0 0.0937999999998 0 -2.0 1e-06 
0.0 0.0938999999998 0 -2.0 1e-06 
0.0 0.0939999999998 0 -2.0 1e-06 
0.0 0.0940999999998 0 -2.0 1e-06 
0.0 0.0941999999998 0 -2.0 1e-06 
0.0 0.0942999999998 0 -2.0 1e-06 
0.0 0.0943999999998 0 -2.0 1e-06 
0.0 0.0944999999998 0 -2.0 1e-06 
0.0 0.0945999999998 0 -2.0 1e-06 
0.0 0.0946999999998 0 -2.0 1e-06 
0.0 0.0947999999998 0 -2.0 1e-06 
0.0 0.0948999999998 0 -2.0 1e-06 
0.0 0.0949999999998 0 -2.0 1e-06 
0.0 0.0950999999998 0 -2.0 1e-06 
0.0 0.0951999999998 0 -2.0 1e-06 
0.0 0.0952999999998 0 -2.0 1e-06 
0.0 0.0953999999998 0 -2.0 1e-06 
0.0 0.0954999999998 0 -2.0 1e-06 
0.0 0.0955999999998 0 -2.0 1e-06 
0.0 0.0956999999998 0 -2.0 1e-06 
0.0 0.0957999999998 0 -2.0 1e-06 
0.0 0.0958999999998 0 -2.0 1e-06 
0.0 0.0959999999998 0 -2.0 1e-06 
0.0 0.0960999999998 0 -2.0 1e-06 
0.0 0.0961999999998 0 -2.0 1e-06 
0.0 0.0962999999998 0 -2.0 1e-06 
0.0 0.0963999999998 0 -2.0 1e-06 
0.0 0.0964999999998 0 -2.0 1e-06 
0.0 0.0965999999998 0 -2.0 1e-06 
0.0 0.0966999999998 0 -2.0 1e-06 
0.0 0.0967999999998 0 -2.0 1e-06 
0.0 0.0968999999998 0 -2.0 1e-06 
0.0 0.0969999999998 0 -2.0 1e-06 
0.0 0.0970999999998 0 -2.0 1e-06 
0.0 0.0971999999998 0 -2.0 1e-06 
0.0 0.0972999999998 0 -2.0 1e-06 
0.0 0.0973999999998 0 -2.0 1e-06 
0.0 0.0974999999998 0 -2.0 1e-06 
0.0 0.0975999999998 0 -2.0 1e-06 
0.0 0.0976999999998 0 -2.0 1e-06 
0.0 0.0977999999998 0 -2.0 1e-06 
0.0 0.0978999999998 0 -2.0 1e-06 
0.0 0.0979999999998 0 -2.0 1e-06 
0.0 0.0980999999998 0 -2.0 1e-06 
0.0 0.0981999999998 0 -2.0 1e-06 
0.0 0.0982999999998 0 -2.0 1e-06 
0.0 0.0983999999998 0 -2.0 1e-06 
0.0 0.0984999999998 0 -2.0 1e-06 
0.0 0.0985999999998 0 -2.0 1e-06 
0.0 0.0986999999998 0 -2.0 1e-06 
0.0 0.0987999999998 0 -2.0 1e-06 
0.0 0.0988999999998 0 -2.0 1e-06 
0.0 0.0989999999998 0 -2.0 1e-06 
0.0 0.0990999999998 0 -2.0 1e-06 
0.0 0.0991999999998 0 -2.0 1e-06 
0.0 0.0992999999998 0 -2.0 1e-06 
0.0 0.0993999999998 0 -2.0 1e-06 
0.0 0.0994999999998 0 -2.0 1e-06 
0.0 0.0995999999998 0 -2.0 1e-06 
0.0 0.0996999999998 0 -2.0 1e-06 
0.0 0.0997999999998 0 -2.0 1e-06 
0.0 0.0998999999998 0 -2.0 1e-06 
0.0 0.0999999999998 0 -2.0 1e-06 
0.0 0.1001 0 -2.0 1e-06 
0.0 0.1002 0 -2.0 1e-06 
0.0 0.1003 0 -2.0 1e-06 
0.0 0.1004 0 -2.0 1e-06 
0.0 0.1005 0 -2.0 1e-06 
0.0 0.1006 0 -2.0 1e-06 
0.0 0.1007 0 -2.0 1e-06 
0.0 0.1008 0 -2.0 1e-06 
0.0 0.1009 0 -2.0 1e-06 
0.0 0.101 0 -2.0 1e-06 
0.0 0.1011 0 -2.0 1e-06 
0.0 0.1012 0 -2.0 1e-06 
0.0 0.1013 0 -2.0 1e-06 
0.0 0.1014 0 -2.0 1e-06 
0.0 0.1015 0 -2.0 1e-06 
0.0 0.1016 0 -2.0 1e-06 
0.0 0.1017 0 -2.0 1e-06 
0.0 0.1018 0 -2.0 1e-06 
0.0 0.1019 0 -2.0 1e-06 
0.0 0.102 0 -2.0 1e-06 
0.0 0.1021 0 -2.0 1e-06 
0.0 0.1022 0 -2.0 1e-06 
0.0 0.1023 0 -2.0 1e-06 
0.0 0.1024 0 -2.0 1e-06 
0.0 0.1025 0 -2.0 1e-06 
0.0 0.1026 0 -2.0 1e-06 
0.0 0.1027 0 -2.0 1e-06 
0.0 0.1028 0 -2.0 1e-06 
0.0 0.1029 0 -2.0 1e-06 
0.0 0.103 0 -2.0 1e-06 
0.0 0.1031 0 -2.0 1e-06 
0.0 0.1032 0 -2.0 1e-06 
0.0 0.1033 0 -2.0 1e-06 
0.0 0.1034 0 -2.0 1e-06 
0.0 0.1035 0 -2.0 1e-06 
0.0 0.1036 0 -2.0 1e-06 
0.0 0.1037 0 -2.0 1e-06 
0.0 0.1038 0 -2.0 1e-06 
0.0 0.1039 0 -2.0 1e-06 
0.0 0.104 0 -2.0 1e-06 
0.0 0.1041 0 -2.0 1e-06 
0.0 0.1042 0 -2.0 1e-06 
0.0 0.1043 0 -2.0 1e-06 
0.0 0.1044 0 -2.0 1e-06 
0.0 0.1045 0 -2.0 1e-06 
0.0 0.1046 0 -2.0 1e-06 
0.0 0.1047 0 -2.0 1e-06 
0.0 0.1048 0 -2.0 1e-06 
0.0 0.1049 0 -2.0 1e-06 
0.0 0.105 0 -2.0 1e-06 
0.0 0.1051 0 -2.0 1e-06 
0.0 0.1052 0 -2.0 1e-06 
0.0 0.1053 0 -2.0 1e-06 
0.0 0.1054 0 -2.0 1e-06 
0.0 0.1055 0 -2.0 1e-06 
0.0 0.1056 0 -2.0 1e-06 
0.0 0.1057 0 -2.0 1e-06 
0.0 0.1058 0 -2.0 1e-06 
0.0 0.1059 0 -2.0 1e-06 
0.0 0.106 0 -2.0 1e-06 
0.0 0.1061 0 -2.0 1e-06 
0.0 0.1062 0 -2.0 1e-06 
0.0 0.1063 0 -2.0 1e-06 
0.0 0.1064 0 -2.0 1e-06 
0.0 0.1065 0 -2.0 1e-06 
0.0 0.1066 0 -2.0 1e-06 
0.0 0.1067 0 -2.0 1e-06 
0.0 0.1068 0 -2.0 1e-06 
0.0 0.1069 0 -2.0 1e-06 
0.0 0.107 0 -2.0 1e-06 
0.0 0.1071 0 -2.0 1e-06 
0.0 0.1072 0 -2.0 1e-06 
0.0 0.1073 0 -2.0 1e-06 
0.0 0.1074 0 -2.0 1e-06 
0.0 0.1075 0 -2.0 1e-06 
0.0 0.1076 0 -2.0 1e-06 
0.0 0.1077 0 -2.0 1e-06 
0.0 0.1078 0 -2.0 1e-06 
0.0 0.1079 0 -2.0 1e-06 
0.0 0.108 0 -2.0 1e-06 
0.0 0.1081 0 -2.0 1e-06 
0.0 0.1082 0 -2.0 1e-06 
0.0 0.1083 0 -2.0 1e-06 
0.0 0.1084 0 -2.0 1e-06 
0.0 0.1085 0 -2.0 1e-06 
0.0 0.1086 0 -2.0 1e-06 
0.0 0.1087 0 -2.0 1e-06 
0.0 0.1088 0 -2.0 1e-06 
0.0 0.1089 0 -2.0 1e-06 
0.0 0.109 0 -2.0 1e-06 
0.0 0.1091 0 -2.0 1e-06 
0.0 0.1092 0 -2.0 1e-06 
0.0 0.1093 0 -2.0 1e-06 
0.0 0.1094 0 -2.0 1e-06 
0.0 0.1095 0 -2.0 1e-06 
0.0 0.1096 0 -2.0 1e-06 
0.0 0.1097 0 -2.0 1e-06 
0.0 0.1098 0 -2.0 1e-06 
0.0 0.1099 0 -2.0 1e-06 
0.0 0.11 0 -2.0 1e-06 
0.0 0.1101 0 -2.0 1e-06 
0.0 0.1102 0 -2.0 1e-06 
0.0 0.1103 0 -2.0 1e-06 
0.0 0.1104 0 -2.0 1e-06 
0.0 0.1105 0 -2.0 1e-06 
0.0 0.1106 0 -2.0 1e-06 
0.0 0.1107 0 -2.0 1e-06 
0.0 0.1108 0 -2.0 1e-06 
0.0 0.1109 0 -2.0 1e-06 
0.0 0.111 0 -2.0 1e-06 
0.0 0.1111 0 -2.0 1e-06 
0.0 0.1112 0 -2.0 1e-06 
0.0 0.1113 0 -2.0 1e-06 
0.0 0.1114 0 -2.0 1e-06 
0.0 0.1115 0 -2.0 1e-06 
0.0 0.1116 0 -2.0 1e-06 
0.0 0.1117 0 -2.0 1e-06 
0.0 0.1118 0 -2.0 1e-06 
0.0 0.1119 0 -2.0 1e-06 
0.0 0.112 0 -2.0 1e-06 
0.0 0.1121 0 -2.0 1e-06 
0.0 0.1122 0 -2.0 1e-06 
0.0 0.1123 0 -2.0 1e-06 
0.0 0.1124 0 -2.0 1e-06 
0.0 0.1125 0 -2.0 1e-06 
0.0 0.1126 0 -2.0 1e-06 
0.0 0.1127 0 -2.0 1e-06 
0.0 0.1128 0 -2.0 1e-06 
0.0 0.1129 0 -2.0 1e-06 
0.0 0.113 0 -2.0 1e-06 
0.0 0.1131 0 -2.0 1e-06 
0.0 0.1132 0 -2.0 1e-06 
0.0 0.1133 0 -2.0 1e-06 
0.0 0.1134 0 -2.0 1e-06 
0.0 0.1135 0 -2.0 1e-06 
0.0 0.1136 0 -2.0 1e-06 
0.0 0.1137 0 -2.0 1e-06 
0.0 0.1138 0 -2.0 1e-06 
0.0 0.1139 0 -2.0 1e-06 
0.0 0.114 0 -2.0 1e-06 
0.0 0.1141 0 -2.0 1e-06 
0.0 0.1142 0 -2.0 1e-06 
0.0 0.1143 0 -2.0 1e-06 
0.0 0.1144 0 -2.0 1e-06 
0.0 0.1145 0 -2.0 1e-06 
0.0 0.1146 0 -2.0 1e-06 
0.0 0.1147 0 -2.0 1e-06 
0.0 0.1148 0 -2.0 1e-06 
0.0 0.1149 0 -2.0 1e-06 
0.0 0.115 0 -2.0 1e-06 
0.0 0.1151 0 -2.0 1e-06 
0.0 0.1152 0 -2.0 1e-06 
0.0 0.1153 0 -2.0 1e-06 
0.0 0.1154 0 -2.0 1e-06 
0.0 0.1155 0 -2.0 1e-06 
0.0 0.1156 0 -2.0 1e-06 
0.0 0.1157 0 -2.0 1e-06 
0.0 0.1158 0 -2.0 1e-06 
0.0 0.1159 0 -2.0 1e-06 
0.0 0.116 0 -2.0 1e-06 
0.0 0.1161 0 -2.0 1e-06 
0.0 0.1162 0 -2.0 1e-06 
0.0 0.1163 0 -2.0 1e-06 
0.0 0.1164 0 -2.0 1e-06 
0.0 0.1165 0 -2.0 1e-06 
0.0 0.1166 0 -2.0 1e-06 
0.0 0.1167 0 -2.0 1e-06 
0.0 0.1168 0 -2.0 1e-06 
0.0 0.1169 0 -2.0 1e-06 
0.0 0.117 0 -2.0 1e-06 
0.0 0.1171 0 -2.0 1e-06 
0.0 0.1172 0 -2.0 1e-06 
0.0 0.1173 0 -2.0 1e-06 
0.0 0.1174 0 -2.0 1e-06 
0.0 0.1175 0 -2.0 1e-06 
0.0 0.1176 0 -2.0 1e-06 
0.0 0.1177 0 -2.0 1e-06 
0.0 0.1178 0 -2.0 1e-06 
0.0 0.1179 0 -2.0 1e-06 
0.0 0.118 0 -2.0 1e-06 
0.0 0.1181 0 -2.0 1e-06 
0.0 0.1182 0 -2.0 1e-06 
0.0 0.1183 0 -2.0 1e-06 
0.0 0.1184 0 -2.0 1e-06 
0.0 0.1185 0 -2.0 1e-06 
0.0 0.1186 0 -2.0 1e-06 
0.0 0.1187 0 -2.0 1e-06 
0.0 0.1188 0 -2.0 1e-06 
0.0 0.1189 0 -2.0 1e-06 
0.0 0.119 0 -2.0 1e-06 
0.0 0.1191 0 -2.0 1e-06 
0.0 0.1192 0 -2.0 1e-06 
0.0 0.1193 0 -2.0 1e-06 
0.0 0.1194 0 -2.0 1e-06 
0.0 0.1195 0 -2.0 1e-06 
0.0 0.1196 0 -2.0 1e-06 
0.0 0.1197 0 -2.0 1e-06 
0.0 0.1198 0 -2.0 1e-06 
0.0 0.1199 0 -2.0 1e-06 
0.0 0.12 0 -2.0 1e-06 
0.0 0.1201 0 -2.0 1e-06 
0.0 0.1202 0 -2.0 1e-06 
0.0 0.1203 0 -2.0 1e-06 
0.0 0.1204 0 -2.0 1e-06 
0.0 0.1205 0 -2.0 1e-06 
0.0 0.1206 0 -2.0 1e-06 
0.0 0.1207 0 -2.0 1e-06 
0.0 0.1208 0 -2.0 1e-06 
0.0 0.1209 0 -2.0 1e-06 
0.0 0.121 0 -2.0 1e-06 
0.0 0.1211 0 -2.0 1e-06 
0.0 0.1212 0 -2.0 1e-06 
0.0 0.1213 0 -2.0 1e-06 
0.0 0.1214 0 -2.0 1e-06 
0.0 0.1215 0 -2.0 1e-06 
0.0 0.1216 0 -2.0 1e-06 
0.0 0.1217 0 -2.0 1e-06 
0.0 0.1218 0 -2.0 1e-06 
0.0 0.1219 0 -2.0 1e-06 
0.0 0.122 0 -2.0 1e-06 
0.0 0.1221 0 -2.0 1e-06 
0.0 0.1222 0 -2.0 1e-06 
0.0 0.1223 0 -2.0 1e-06 
0.0 0.1224 0 -2.0 1e-06 
0.0 0.1225 0 -2.0 1e-06 
0.0 0.1226 0 -2.0 1e-06 
0.0 0.1227 0 -2.0 1e-06 
0.0 0.1228 0 -2.0 1e-06 
0.0 0.1229 0 -2.0 1e-06 
0.0 0.123 0 -2.0 1e-06 
0.0 0.1231 0 -2.0 1e-06 
0.0 0.1232 0 -2.0 1e-06 
0.0 0.1233 0 -2.0 1e-06 
0.0 0.1234 0 -2.0 1e-06 
0.0 0.1235 0 -2.0 1e-06 
0.0 0.1236 0 -2.0 1e-06 
0.0 0.1237 0 -2.0 1e-06 
0.0 0.1238 0 -2.0 1e-06 
0.0 0.1239 0 -2.0 1e-06 
0.0 0.124 0 -2.0 1e-06 
0.0 0.1241 0 -2.0 1e-06 
0.0 0.1242 0 -2.0 1e-06 
0.0 0.1243 0 -2.0 1e-06 
0.0 0.1244 0 -2.0 1e-06 
0.0 0.1245 0 -2.0 1e-06 
0.0 0.1246 0 -2.0 1e-06 
0.0 0.1247 0 -2.0 1e-06 
0.0 0.1248 0 -2.0 1e-06 
0.0 0.1249 0 -2.0 1e-06 
0.0 0.125 0 -2.0 1e-06 
0.0 0.1251 0 -2.0 1e-06 
0.0 0.1252 0 -2.0 1e-06 
0.0 0.1253 0 -2.0 1e-06 
0.0 0.1254 0 -2.0 1e-06 
0.0 0.1255 0 -2.0 1e-06 
0.0 0.1256 0 -2.0 1e-06 
0.0 0.1257 0 -2.0 1e-06 
0.0 0.1258 0 -2.0 1e-06 
0.0 0.1259 0 -2.0 1e-06 
0.0 0.126 0 -2.0 1e-06 
0.0 0.1261 0 -2.0 1e-06 
0.0 0.1262 0 -2.0 1e-06 
0.0 0.1263 0 -2.0 1e-06 
0.0 0.1264 0 -2.0 1e-06 
0.0 0.1265 0 -2.0 1e-06 
0.0 0.1266 0 -2.0 1e-06 
0.0 0.1267 0 -2.0 1e-06 
0.0 0.1268 0 -2.0 1e-06 
0.0 0.1269 0 -2.0 1e-06 
0.0 0.127 0 -2.0 1e-06 
0.0 0.1271 0 -2.0 1e-06 
0.0 0.1272 0 -2.0 1e-06 
0.0 0.1273 0 -2.0 1e-06 
0.0 0.1274 0 -2.0 1e-06 
0.0 0.1275 0 -2.0 1e-06 
0.0 0.1276 0 -2.0 1e-06 
0.0 0.1277 0 -2.0 1e-06 
0.0 0.1278 0 -2.0 1e-06 
0.0 0.1279 0 -2.0 1e-06 
0.0 0.128 0 -2.0 1e-06 
0.0 0.1281 0 -2.0 1e-06 
0.0 0.1282 0 -2.0 1e-06 
0.0 0.1283 0 -2.0 1e-06 
0.0 0.1284 0 -2.0 1e-06 
0.0 0.1285 0 -2.0 1e-06 
0.0 0.1286 0 -2.0 1e-06 
0.0 0.1287 0 -2.0 1e-06 
0.0 0.1288 0 -2.0 1e-06 
0.0 0.1289 0 -2.0 1e-06 
0.0 0.129 0 -2.0 1e-06 
0.0 0.1291 0 -2.0 1e-06 
0.0 0.1292 0 -2.0 1e-06 
0.0 0.1293 0 -2.0 1e-06 
0.0 0.1294 0 -2.0 1e-06 
0.0 0.1295 0 -2.0 1e-06 
0.0 0.1296 0 -2.0 1e-06 
0.0 0.1297 0 -2.0 1e-06 
0.0 0.1298 0 -2.0 1e-06 
0.0 0.1299 0 -2.0 1e-06 
0.0 0.13 0 -2.0 1e-06 
0.0 0.1301 0 -2.0 1e-06 
0.0 0.1302 0 -2.0 1e-06 
0.0 0.1303 0 -2.0 1e-06 
0.0 0.1304 0 -2.0 1e-06 
0.0 0.1305 0 -2.0 1e-06 
0.0 0.1306 0 -2.0 1e-06 
0.0 0.1307 0 -2.0 1e-06 
0.0 0.1308 0 -2.0 1e-06 
0.0 0.1309 0 -2.0 1e-06 
0.0 0.131 0 -2.0 1e-06 
0.0 0.1311 0 -2.0 1e-06 
0.0 0.1312 0 -2.0 1e-06 
0.0 0.1313 0 -2.0 1e-06 
0.0 0.1314 0 -2.0 1e-06 
0.0 0.1315 0 -2.0 1e-06 
0.0 0.1316 0 -2.0 1e-06 
0.0 0.1317 0 -2.0 1e-06 
0.0 0.1318 0 -2.0 1e-06 
0.0 0.1319 0 -2.0 1e-06 
0.0 0.132 0 -2.0 1e-06 
0.0 0.1321 0 -2.0 1e-06 
0.0 0.1322 0 -2.0 1e-06 
0.0 0.1323 0 -2.0 1e-06 
0.0 0.1324 0 -2.0 1e-06 
0.0 0.1325 0 -2.0 1e-06 
0.0 0.1326 0 -2.0 1e-06 
0.0 0.1327 0 -2.0 1e-06 
0.0 0.1328 0 -2.0 1e-06 
0.0 0.1329 0 -2.0 1e-06 
0.0 0.133 0 -2.0 1e-06 
0.0 0.1331 0 -2.0 1e-06 
0.0 0.1332 0 -2.0 1e-06 
0.0 0.1333 0 -2.0 1e-06 
0.0 0.1334 0 -2.0 1e-06 
0.0 0.1335 0 -2.0 1e-06 
0.0 0.1336 0 -2.0 1e-06 
0.0 0.1337 0 -2.0 1e-06 
0.0 0.1338 0 -2.0 1e-06 
0.0 0.1339 0 -2.0 1e-06 
0.0 0.134 0 -2.0 1e-06 
0.0 0.1341 0 -2.0 1e-06 
0.0 0.1342 0 -2.0 1e-06 
0.0 0.1343 0 -2.0 1e-06 
0.0 0.1344 0 -2.0 1e-06 
0.0 0.1345 0 -2.0 1e-06 
0.0 0.1346 0 -2.0 1e-06 
0.0 0.1347 0 -2.0 1e-06 
0.0 0.1348 0 -2.0 1e-06 
0.0 0.1349 0 -2.0 1e-06 
0.0 0.135 0 -2.0 1e-06 
0.0 0.1351 0 -2.0 1e-06 
0.0 0.1352 0 -2.0 1e-06 
0.0 0.1353 0 -2.0 1e-06 
0.0 0.1354 0 -2.0 1e-06 
0.0 0.1355 0 -2.0 1e-06 
0.0 0.1356 0 -2.0 1e-06 
0.0 0.1357 0 -2.0 1e-06 
0.0 0.1358 0 -2.0 1e-06 
0.0 0.1359 0 -2.0 1e-06 
0.0 0.136 0 -2.0 1e-06 
0.0 0.1361 0 -2.0 1e-06 
0.0 0.1362 0 -2.0 1e-06 
0.0 0.1363 0 -2.0 1e-06 
0.0 0.1364 0 -2.0 1e-06 
0.0 0.1365 0 -2.0 1e-06 
0.0 0.1366 0 -2.0 1e-06 
0.0 0.1367 0 -2.0 1e-06 
0.0 0.1368 0 -2.0 1e-06 
0.0 0.1369 0 -2.0 1e-06 
0.0 0.137 0 -2.0 1e-06 
0.0 0.1371 0 -2.0 1e-06 
0.0 0.1372 0 -2.0 1e-06 
0.0 0.1373 0 -2.0 1e-06 
0.0 0.1374 0 -2.0 1e-06 
0.0 0.1375 0 -2.0 1e-06 
0.0 0.1376 0 -2.0 1e-06 
0.0 0.1377 0 -2.0 1e-06 
0.0 0.1378 0 -2.0 1e-06 
0.0 0.1379 0 -2.0 1e-06 
0.0 0.138 0 -2.0 1e-06 
0.0 0.1381 0 -2.0 1e-06 
0.0 0.1382 0 -2.0 1e-06 
0.0 0.1383 0 -2.0 1e-06 
0.0 0.1384 0 -2.0 1e-06 
0.0 0.1385 0 -2.0 1e-06 
0.0 0.1386 0 -2.0 1e-06 
0.0 0.1387 0 -2.0 1e-06 
0.0 0.1388 0 -2.0 1e-06 
0.0 0.1389 0 -2.0 1e-06 
0.0 0.139 0 -2.0 1e-06 
0.0 0.1391 0 -2.0 1e-06 
0.0 0.1392 0 -2.0 1e-06 
0.0 0.1393 0 -2.0 1e-06 
0.0 0.1394 0 -2.0 1e-06 
0.0 0.1395 0 -2.0 1e-06 
0.0 0.1396 0 -2.0 1e-06 
0.0 0.1397 0 -2.0 1e-06 
0.0 0.1398 0 -2.0 1e-06 
0.0 0.1399 0 -2.0 1e-06 
0.0 0.14 0 -2.0 1e-06 
0.0 0.1401 0 -2.0 1e-06 
0.0 0.1402 0 -2.0 1e-06 
0.0 0.1403 0 -2.0 1e-06 
0.0 0.1404 0 -2.0 1e-06 
0.0 0.1405 0 -2.0 1e-06 
0.0 0.1406 0 -2.0 1e-06 
0.0 0.1407 0 -2.0 1e-06 
0.0 0.1408 0 -2.0 1e-06 
0.0 0.1409 0 -2.0 1e-06 
0.0 0.141 0 -2.0 1e-06 
0.0 0.1411 0 -2.0 1e-06 
0.0 0.1412 0 -2.0 1e-06 
0.0 0.1413 0 -2.0 1e-06 
0.0 0.1414 0 -2.0 1e-06 
0.0 0.1415 0 -2.0 1e-06 
0.0 0.1416 0 -2.0 1e-06 
0.0 0.1417 0 -2.0 1e-06 
0.0 0.1418 0 -2.0 1e-06 
0.0 0.1419 0 -2.0 1e-06 
0.0 0.142 0 -2.0 1e-06 
0.0 0.1421 0 -2.0 1e-06 
0.0 0.1422 0 -2.0 1e-06 
0.0 0.1423 0 -2.0 1e-06 
0.0 0.1424 0 -2.0 1e-06 
0.0 0.1425 0 -2.0 1e-06 
0.0 0.1426 0 -2.0 1e-06 
0.0 0.1427 0 -2.0 1e-06 
0.0 0.1428 0 -2.0 1e-06 
0.0 0.1429 0 -2.0 1e-06 
0.0 0.143 0 -2.0 1e-06 
0.0 0.1431 0 -2.0 1e-06 
0.0 0.1432 0 -2.0 1e-06 
0.0 0.1433 0 -2.0 1e-06 
0.0 0.1434 0 -2.0 1e-06 
0.0 0.1435 0 -2.0 1e-06 
0.0 0.1436 0 -2.0 1e-06 
0.0 0.1437 0 -2.0 1e-06 
0.0 0.1438 0 -2.0 1e-06 
0.0 0.1439 0 -2.0 1e-06 
0.0 0.144 0 -2.0 1e-06 
0.0 0.1441 0 -2.0 1e-06 
0.0 0.1442 0 -2.0 1e-06 
0.0 0.1443 0 -2.0 1e-06 
0.0 0.1444 0 -2.0 1e-06 
0.0 0.1445 0 -2.0 1e-06 
0.0 0.1446 0 -2.0 1e-06 
0.0 0.1447 0 -2.0 1e-06 
0.0 0.1448 0 -2.0 1e-06 
0.0 0.1449 0 -2.0 1e-06 
0.0 0.145 0 -2.0 1e-06 
0.0 0.1451 0 -2.0 1e-06 
0.0 0.1452 0 -2.0 1e-06 
0.0 0.1453 0 -2.0 1e-06 
0.0 0.1454 0 -2.0 1e-06 
0.0 0.1455 0 -2.0 1e-06 
0.0 0.1456 0 -2.0 1e-06 
0.0 0.1457 0 -2.0 1e-06 
0.0 0.1458 0 -2.0 1e-06 
0.0 0.1459 0 -2.0 1e-06 
0.0 0.146 0 -2.0 1e-06 
0.0 0.1461 0 -2.0 1e-06 
0.0 0.1462 0 -2.0 1e-06 
0.0 0.1463 0 -2.0 1e-06 
0.0 0.1464 0 -2.0 1e-06 
0.0 0.1465 0 -2.0 1e-06 
0.0 0.1466 0 -2.0 1e-06 
0.0 0.1467 0 -2.0 1e-06 
0.0 0.1468 0 -2.0 1e-06 
0.0 0.1469 0 -2.0 1e-06 
0.0 0.147 0 -2.0 1e-06 
0.0 0.1471 0 -2.0 1e-06 
0.0 0.1472 0 -2.0 1e-06 
0.0 0.1473 0 -2.0 1e-06 
0.0 0.1474 0 -2.0 1e-06 
0.0 0.1475 0 -2.0 1e-06 
0.0 0.1476 0 -2.0 1e-06 
0.0 0.1477 0 -2.0 1e-06 
0.0 0.1478 0 -2.0 1e-06 
0.0 0.1479 0 -2.0 1e-06 
0.0 0.148 0 -2.0 1e-06 
0.0 0.1481 0 -2.0 1e-06 
0.0 0.1482 0 -2.0 1e-06 
0.0 0.1483 0 -2.0 1e-06 
0.0 0.1484 0 -2.0 1e-06 
0.0 0.1485 0 -2.0 1e-06 
0.0 0.1486 0 -2.0 1e-06 
0.0 0.1487 0 -2.0 1e-06 
0.0 0.1488 0 -2.0 1e-06 
0.0 0.1489 0 -2.0 1e-06 
0.0 0.149 0 -2.0 1e-06 
0.0 0.1491 0 -2.0 1e-06 
0.0 0.1492 0 -2.0 1e-06 
0.0 0.1493 0 -2.0 1e-06 
0.0 0.1494 0 -2.0 1e-06 
0.0 0.1495 0 -2.0 1e-06 
0.0 0.1496 0 -2.0 1e-06 
0.0 0.1497 0 -2.0 1e-06 
0.0 0.1498 0 -2.0 1e-06 
0.0 0.1499 0 -2.0 1e-06 
0.0 0.15 0 -2.0 1e-06 
0.0 0.1501 0 -2.0 1e-06 
0.0 0.1502 0 -2.0 1e-06 
0.0 0.1503 0 -2.0 1e-06 
0.0 0.1504 0 -2.0 1e-06 
0.0 0.1505 0 -2.0 1e-06 
0.0 0.1506 0 -2.0 1e-06 
0.0 0.1507 0 -2.0 1e-06 
0.0 0.1508 0 -2.0 1e-06 
0.0 0.1509 0 -2.0 1e-06 
0.0 0.151 0 -2.0 1e-06 
0.0 0.1511 0 -2.0 1e-06 
0.0 0.1512 0 -2.0 1e-06 
0.0 0.1513 0 -2.0 1e-06 
0.0 0.1514 0 -2.0 1e-06 
0.0 0.1515 0 -2.0 1e-06 
0.0 0.1516 0 -2.0 1e-06 
0.0 0.1517 0 -2.0 1e-06 
0.0 0.1518 0 -2.0 1e-06 
0.0 0.1519 0 -2.0 1e-06 
0.0 0.152 0 -2.0 1e-06 
0.0 0.1521 0 -2.0 1e-06 
0.0 0.1522 0 -2.0 1e-06 
0.0 0.1523 0 -2.0 1e-06 
0.0 0.1524 0 -2.0 1e-06 
0.0 0.1525 0 -2.0 1e-06 
0.0 0.1526 0 -2.0 1e-06 
0.0 0.1527 0 -2.0 1e-06 
0.0 0.1528 0 -2.0 1e-06 
0.0 0.1529 0 -2.0 1e-06 
0.0 0.153 0 -2.0 1e-06 
0.0 0.1531 0 -2.0 1e-06 
0.0 0.1532 0 -2.0 1e-06 
0.0 0.1533 0 -2.0 1e-06 
0.0 0.1534 0 -2.0 1e-06 
0.0 0.1535 0 -2.0 1e-06 
0.0 0.1536 0 -2.0 1e-06 
0.0 0.1537 0 -2.0 1e-06 
0.0 0.1538 0 -2.0 1e-06 
0.0 0.1539 0 -2.0 1e-06 
0.0 0.154 0 -2.0 1e-06 
0.0 0.1541 0 -2.0 1e-06 
0.0 0.1542 0 -2.0 1e-06 
0.0 0.1543 0 -2.0 1e-06 
0.0 0.1544 0 -2.0 1e-06 
0.0 0.1545 0 -2.0 1e-06 
0.0 0.1546 0 -2.0 1e-06 
0.0 0.1547 0 -2.0 1e-06 
0.0 0.1548 0 -2.0 1e-06 
0.0 0.1549 0 -2.0 1e-06 
0.0 0.155 0 -2.0 1e-06 
0.0 0.1551 0 -2.0 1e-06 
0.0 0.1552 0 -2.0 1e-06 
0.0 0.1553 0 -2.0 1e-06 
0.0 0.1554 0 -2.0 1e-06 
0.0 0.1555 0 -2.0 1e-06 
0.0 0.1556 0 -2.0 1e-06 
0.0 0.1557 0 -2.0 1e-06 
0.0 0.1558 0 -2.0 1e-06 
0.0 0.1559 0 -2.0 1e-06 
0.0 0.156 0 -2.0 1e-06 
0.0 0.1561 0 -2.0 1e-06 
0.0 0.1562 0 -2.0 1e-06 
0.0 0.1563 0 -2.0 1e-06 
0.0 0.1564 0 -2.0 1e-06 
0.0 0.1565 0 -2.0 1e-06 
0.0 0.1566 0 -2.0 1e-06 
0.0 0.1567 0 -2.0 1e-06 
0.0 0.1568 0 -2.0 1e-06 
0.0 0.1569 0 -2.0 1e-06 
0.0 0.157 0 -2.0 1e-06 
0.0 0.1571 0 -2.0 1e-06 
0.0 0.1572 0 -2.0 1e-06 
0.0 0.1573 0 -2.0 1e-06 
0.0 0.1574 0 -2.0 1e-06 
0.0 0.1575 0 -2.0 1e-06 
0.0 0.1576 0 -2.0 1e-06 
0.0 0.1577 0 -2.0 1e-06 
0.0 0.1578 0 -2.0 1e-06 
0.0 0.1579 0 -2.0 1e-06 
0.0 0.158 0 -2.0 1e-06 
0.0 0.1581 0 -2.0 1e-06 
0.0 0.1582 0 -2.0 1e-06 
0.0 0.1583 0 -2.0 1e-06 
0.0 0.1584 0 -2.0 1e-06 
0.0 0.1585 0 -2.0 1e-06 
0.0 0.1586 0 -2.0 1e-06 
0.0 0.1587 0 -2.0 1e-06 
0.0 0.1588 0 -2.0 1e-06 
0.0 0.1589 0 -2.0 1e-06 
0.0 0.159 0 -2.0 1e-06 
0.0 0.1591 0 -2.0 1e-06 
0.0 0.1592 0 -2.0 1e-06 
0.0 0.1593 0 -2.0 1e-06 
0.0 0.1594 0 -2.0 1e-06 
0.0 0.1595 0 -2.0 1e-06 
0.0 0.1596 0 -2.0 1e-06 
0.0 0.1597 0 -2.0 1e-06 
0.0 0.1598 0 -2.0 1e-06 
0.0 0.1599 0 -2.0 1e-06 
0.0 0.16 0 -2.0 1e-06 
0.0 0.1601 0 -2.0 1e-06 
0.0 0.1602 0 -2.0 1e-06 
0.0 0.1603 0 -2.0 1e-06 
0.0 0.1604 0 -2.0 1e-06 
0.0 0.1605 0 -2.0 1e-06 
0.0 0.1606 0 -2.0 1e-06 
0.0 0.1607 0 -2.0 1e-06 
0.0 0.1608 0 -2.0 1e-06 
0.0 0.1609 0 -2.0 1e-06 
0.0 0.161 0 -2.0 1e-06 
0.0 0.1611 0 -2.0 1e-06 
0.0 0.1612 0 -2.0 1e-06 
0.0 0.1613 0 -2.0 1e-06 
0.0 0.1614 0 -2.0 1e-06 
0.0 0.1615 0 -2.0 1e-06 
0.0 0.1616 0 -2.0 1e-06 
0.0 0.1617 0 -2.0 1e-06 
0.0 0.1618 0 -2.0 1e-06 
0.0 0.1619 0 -2.0 1e-06 
0.0 0.162 0 -2.0 1e-06 
0.0 0.1621 0 -2.0 1e-06 
0.0 0.1622 0 -2.0 1e-06 
0.0 0.1623 0 -2.0 1e-06 
0.0 0.1624 0 -2.0 1e-06 
0.0 0.1625 0 -2.0 1e-06 
0.0 0.1626 0 -2.0 1e-06 
0.0 0.1627 0 -2.0 1e-06 
0.0 0.1628 0 -2.0 1e-06 
0.0 0.1629 0 -2.0 1e-06 
0.0 0.163 0 -2.0 1e-06 
0.0 0.1631 0 -2.0 1e-06 
0.0 0.1632 0 -2.0 1e-06 
0.0 0.1633 0 -2.0 1e-06 
0.0 0.1634 0 -2.0 1e-06 
0.0 0.1635 0 -2.0 1e-06 
0.0 0.1636 0 -2.0 1e-06 
0.0 0.1637 0 -2.0 1e-06 
0.0 0.1638 0 -2.0 1e-06 
0.0 0.1639 0 -2.0 1e-06 
0.0 0.164 0 -2.0 1e-06 
0.0 0.1641 0 -2.0 1e-06 
0.0 0.1642 0 -2.0 1e-06 
0.0 0.1643 0 -2.0 1e-06 
0.0 0.1644 0 -2.0 1e-06 
0.0 0.1645 0 -2.0 1e-06 
0.0 0.1646 0 -2.0 1e-06 
0.0 0.1647 0 -2.0 1e-06 
0.0 0.1648 0 -2.0 1e-06 
0.0 0.1649 0 -2.0 1e-06 
0.0 0.165 0 -2.0 1e-06 
0.0 0.1651 0 -2.0 1e-06 
0.0 0.1652 0 -2.0 1e-06 
0.0 0.1653 0 -2.0 1e-06 
0.0 0.1654 0 -2.0 1e-06 
0.0 0.1655 0 -2.0 1e-06 
0.0 0.1656 0 -2.0 1e-06 
0.0 0.1657 0 -2.0 1e-06 
0.0 0.1658 0 -2.0 1e-06 
0.0 0.1659 0 -2.0 1e-06 
0.0 0.166 0 -2.0 1e-06 
0.0 0.1661 0 -2.0 1e-06 
0.0 0.1662 0 -2.0 1e-06 
0.0 0.1663 0 -2.0 1e-06 
0.0 0.1664 0 -2.0 1e-06 
0.0 0.1665 0 -2.0 1e-06 
0.0 0.1666 0 -2.0 1e-06 
0.0 0.1667 0 -2.0 1e-06 
0.0 0.1668 0 -2.0 1e-06 
0.0 0.1669 0 -2.0 1e-06 
0.0 0.167 0 -2.0 1e-06 
0.0 0.1671 0 -2.0 1e-06 
0.0 0.1672 0 -2.0 1e-06 
0.0 0.1673 0 -2.0 1e-06 
0.0 0.1674 0 -2.0 1e-06 
0.0 0.1675 0 -2.0 1e-06 
0.0 0.1676 0 -2.0 1e-06 
0.0 0.1677 0 -2.0 1e-06 
0.0 0.1678 0 -2.0 1e-06 
0.0 0.1679 0 -2.0 1e-06 
0.0 0.168 0 -2.0 1e-06 
0.0 0.1681 0 -2.0 1e-06 
0.0 0.1682 0 -2.0 1e-06 
0.0 0.1683 0 -2.0 1e-06 
0.0 0.1684 0 -2.0 1e-06 
0.0 0.1685 0 -2.0 1e-06 
0.0 0.1686 0 -2.0 1e-06 
0.0 0.1687 0 -2.0 1e-06 
0.0 0.1688 0 -2.0 1e-06 
0.0 0.1689 0 -2.0 1e-06 
0.0 0.169 0 -2.0 1e-06 
0.0 0.1691 0 -2.0 1e-06 
0.0 0.1692 0 -2.0 1e-06 
0.0 0.1693 0 -2.0 1e-06 
0.0 0.1694 0 -2.0 1e-06 
0.0 0.1695 0 -2.0 1e-06 
0.0 0.1696 0 -2.0 1e-06 
0.0 0.1697 0 -2.0 1e-06 
0.0 0.1698 0 -2.0 1e-06 
0.0 0.1699 0 -2.0 1e-06 
0.0 0.17 0 -2.0 1e-06 
0.0 0.1701 0 -2.0 1e-06 
0.0 0.1702 0 -2.0 1e-06 
0.0 0.1703 0 -2.0 1e-06 
0.0 0.1704 0 -2.0 1e-06 
0.0 0.1705 0 -2.0 1e-06 
0.0 0.1706 0 -2.0 1e-06 
0.0 0.1707 0 -2.0 1e-06 
0.0 0.1708 0 -2.0 1e-06 
0.0 0.1709 0 -2.0 1e-06 
0.0 0.171 0 -2.0 1e-06 
0.0 0.1711 0 -2.0 1e-06 
0.0 0.1712 0 -2.0 1e-06 
0.0 0.1713 0 -2.0 1e-06 
0.0 0.1714 0 -2.0 1e-06 
0.0 0.1715 0 -2.0 1e-06 
0.0 0.1716 0 -2.0 1e-06 
0.0 0.1717 0 -2.0 1e-06 
0.0 0.1718 0 -2.0 1e-06 
0.0 0.1719 0 -2.0 1e-06 
0.0 0.172 0 -2.0 1e-06 
0.0 0.1721 0 -2.0 1e-06 
0.0 0.1722 0 -2.0 1e-06 
0.0 0.1723 0 -2.0 1e-06 
0.0 0.1724 0 -2.0 1e-06 
0.0 0.1725 0 -2.0 1e-06 
0.0 0.1726 0 -2.0 1e-06 
0.0 0.1727 0 -2.0 1e-06 
0.0 0.1728 0 -2.0 1e-06 
0.0 0.1729 0 -2.0 1e-06 
0.0 0.173 0 -2.0 1e-06 
0.0 0.1731 0 -2.0 1e-06 
0.0 0.1732 0 -2.0 1e-06 
0.0 0.1733 0 -2.0 1e-06 
0.0 0.1734 0 -2.0 1e-06 
0.0 0.1735 0 -2.0 1e-06 
0.0 0.1736 0 -2.0 1e-06 
0.0 0.1737 0 -2.0 1e-06 
0.0 0.1738 0 -2.0 1e-06 
0.0 0.1739 0 -2.0 1e-06 
0.0 0.174 0 -2.0 1e-06 
0.0 0.1741 0 -2.0 1e-06 
0.0 0.1742 0 -2.0 1e-06 
0.0 0.1743 0 -2.0 1e-06 
0.0 0.1744 0 -2.0 1e-06 
0.0 0.1745 0 -2.0 1e-06 
0.0 0.1746 0 -2.0 1e-06 
0.0 0.1747 0 -2.0 1e-06 
0.0 0.1748 0 -2.0 1e-06 
0.0 0.1749 0 -2.0 1e-06 
0.0 0.175 0 -2.0 1e-06 
0.0 0.1751 0 -2.0 1e-06 
0.0 0.1752 0 -2.0 1e-06 
0.0 0.1753 0 -2.0 1e-06 
0.0 0.1754 0 -2.0 1e-06 
0.0 0.1755 0 -2.0 1e-06 
0.0 0.1756 0 -2.0 1e-06 
0.0 0.1757 0 -2.0 1e-06 
0.0 0.1758 0 -2.0 1e-06 
0.0 0.1759 0 -2.0 1e-06 
0.0 0.176 0 -2.0 1e-06 
0.0 0.1761 0 -2.0 1e-06 
0.0 0.1762 0 -2.0 1e-06 
0.0 0.1763 0 -2.0 1e-06 
0.0 0.1764 0 -2.0 1e-06 
0.0 0.1765 0 -2.0 1e-06 
0.0 0.1766 0 -2.0 1e-06 
0.0 0.1767 0 -2.0 1e-06 
0.0 0.1768 0 -2.0 1e-06 
0.0 0.1769 0 -2.0 1e-06 
0.0 0.177 0 -2.0 1e-06 
0.0 0.1771 0 -2.0 1e-06 
0.0 0.1772 0 -2.0 1e-06 
0.0 0.1773 0 -2.0 1e-06 
0.0 0.1774 0 -2.0 1e-06 
0.0 0.1775 0 -2.0 1e-06 
0.0 0.1776 0 -2.0 1e-06 
0.0 0.1777 0 -2.0 1e-06 
0.0 0.1778 0 -2.0 1e-06 
0.0 0.1779 0 -2.0 1e-06 
0.0 0.178 0 -2.0 1e-06 
0.0 0.1781 0 -2.0 1e-06 
0.0 0.1782 0 -2.0 1e-06 
0.0 0.1783 0 -2.0 1e-06 
0.0 0.1784 0 -2.0 1e-06 
0.0 0.1785 0 -2.0 1e-06 
0.0 0.1786 0 -2.0 1e-06 
0.0 0.1787 0 -2.0 1e-06 
0.0 0.1788 0 -2.0 1e-06 
0.0 0.1789 0 -2.0 1e-06 
0.0 0.179 0 -2.0 1e-06 
0.0 0.1791 0 -2.0 1e-06 
0.0 0.1792 0 -2.0 1e-06 
0.0 0.1793 0 -2.0 1e-06 
0.0 0.1794 0 -2.0 1e-06 
0.0 0.1795 0 -2.0 1e-06 
0.0 0.1796 0 -2.0 1e-06 
0.0 0.1797 0 -2.0 1e-06 
0.0 0.1798 0 -2.0 1e-06 
0.0 0.1799 0 -2.0 1e-06 
0.0 0.18 0 -2.0 1e-06 
0.0 0.1801 0 -2.0 1e-06 
0.0 0.1802 0 -2.0 1e-06 
0.0 0.1803 0 -2.0 1e-06 
0.0 0.1804 0 -2.0 1e-06 
0.0 0.1805 0 -2.0 1e-06 
0.0 0.1806 0 -2.0 1e-06 
0.0 0.1807 0 -2.0 1e-06 
0.0 0.1808 0 -2.0 1e-06 
0.0 0.1809 0 -2.0 1e-06 
0.0 0.181 0 -2.0 1e-06 
0.0 0.1811 0 -2.0 1e-06 
0.0 0.1812 0 -2.0 1e-06 
0.0 0.1813 0 -2.0 1e-06 
0.0 0.1814 0 -2.0 1e-06 
0.0 0.1815 0 -2.0 1e-06 
0.0 0.1816 0 -2.0 1e-06 
0.0 0.1817 0 -2.0 1e-06 
0.0 0.1818 0 -2.0 1e-06 
0.0 0.1819 0 -2.0 1e-06 
0.0 0.182 0 -2.0 1e-06 
0.0 0.1821 0 -2.0 1e-06 
0.0 0.1822 0 -2.0 1e-06 
0.0 0.1823 0 -2.0 1e-06 
0.0 0.1824 0 -2.0 1e-06 
0.0 0.1825 0 -2.0 1e-06 
0.0 0.1826 0 -2.0 1e-06 
0.0 0.1827 0 -2.0 1e-06 
0.0 0.1828 0 -2.0 1e-06 
0.0 0.1829 0 -2.0 1e-06 
0.0 0.183 0 -2.0 1e-06 
0.0 0.1831 0 -2.0 1e-06 
0.0 0.1832 0 -2.0 1e-06 
0.0 0.1833 0 -2.0 1e-06 
0.0 0.1834 0 -2.0 1e-06 
0.0 0.1835 0 -2.0 1e-06 
0.0 0.1836 0 -2.0 1e-06 
0.0 0.1837 0 -2.0 1e-06 
0.0 0.1838 0 -2.0 1e-06 
0.0 0.1839 0 -2.0 1e-06 
0.0 0.184 0 -2.0 1e-06 
0.0 0.1841 0 -2.0 1e-06 
0.0 0.1842 0 -2.0 1e-06 
0.0 0.1843 0 -2.0 1e-06 
0.0 0.1844 0 -2.0 1e-06 
0.0 0.1845 0 -2.0 1e-06 
0.0 0.1846 0 -2.0 1e-06 
0.0 0.1847 0 -2.0 1e-06 
0.0 0.1848 0 -2.0 1e-06 
0.0 0.1849 0 -2.0 1e-06 
0.0 0.185 0 -2.0 1e-06 
0.0 0.1851 0 -2.0 1e-06 
0.0 0.1852 0 -2.0 1e-06 
0.0 0.1853 0 -2.0 1e-06 
0.0 0.1854 0 -2.0 1e-06 
0.0 0.1855 0 -2.0 1e-06 
0.0 0.1856 0 -2.0 1e-06 
0.0 0.1857 0 -2.0 1e-06 
0.0 0.1858 0 -2.0 1e-06 
0.0 0.1859 0 -2.0 1e-06 
0.0 0.186 0 -2.0 1e-06 
0.0 0.1861 0 -2.0 1e-06 
0.0 0.1862 0 -2.0 1e-06 
0.0 0.1863 0 -2.0 1e-06 
0.0 0.1864 0 -2.0 1e-06 
0.0 0.1865 0 -2.0 1e-06 
0.0 0.1866 0 -2.0 1e-06 
0.0 0.1867 0 -2.0 1e-06 
0.0 0.1868 0 -2.0 1e-06 
0.0 0.1869 0 -2.0 1e-06 
0.0 0.187 0 -2.0 1e-06 
0.0 0.1871 0 -2.0 1e-06 
0.0 0.1872 0 -2.0 1e-06 
0.0 0.1873 0 -2.0 1e-06 
0.0 0.1874 0 -2.0 1e-06 
0.0 0.1875 0 -2.0 1e-06 
0.0 0.1876 0 -2.0 1e-06 
0.0 0.1877 0 -2.0 1e-06 
0.0 0.1878 0 -2.0 1e-06 
0.0 0.1879 0 -2.0 1e-06 
0.0 0.188 0 -2.0 1e-06 
0.0 0.1881 0 -2.0 1e-06 
0.0 0.1882 0 -2.0 1e-06 
0.0 0.1883 0 -2.0 1e-06 
0.0 0.1884 0 -2.0 1e-06 
0.0 0.1885 0 -2.0 1e-06 
0.0 0.1886 0 -2.0 1e-06 
0.0 0.1887 0 -2.0 1e-06 
0.0 0.1888 0 -2.0 1e-06 
0.0 0.1889 0 -2.0 1e-06 
0.0 0.189 0 -2.0 1e-06 
0.0 0.1891 0 -2.0 1e-06 
0.0 0.1892 0 -2.0 1e-06 
0.0 0.1893 0 -2.0 1e-06 
0.0 0.1894 0 -2.0 1e-06 
0.0 0.1895 0 -2.0 1e-06 
0.0 0.1896 0 -2.0 1e-06 
0.0 0.1897 0 -2.0 1e-06 
0.0 0.1898 0 -2.0 1e-06 
0.0 0.1899 0 -2.0 1e-06 
0.0 0.19 0 -2.0 1e-06 
0.0 0.1901 0 -2.0 1e-06 
0.0 0.1902 0 -2.0 1e-06 
0.0 0.1903 0 -2.0 1e-06 
0.0 0.1904 0 -2.0 1e-06 
0.0 0.1905 0 -2.0 1e-06 
0.0 0.1906 0 -2.0 1e-06 
0.0 0.1907 0 -2.0 1e-06 
0.0 0.1908 0 -2.0 1e-06 
0.0 0.1909 0 -2.0 1e-06 
0.0 0.191 0 -2.0 1e-06 
0.0 0.1911 0 -2.0 1e-06 
0.0 0.1912 0 -2.0 1e-06 
0.0 0.1913 0 -2.0 1e-06 
0.0 0.1914 0 -2.0 1e-06 
0.0 0.1915 0 -2.0 1e-06 
0.0 0.1916 0 -2.0 1e-06 
0.0 0.1917 0 -2.0 1e-06 
0.0 0.1918 0 -2.0 1e-06 
0.0 0.1919 0 -2.0 1e-06 
0.0 0.192 0 -2.0 1e-06 
0.0 0.1921 0 -2.0 1e-06 
0.0 0.1922 0 -2.0 1e-06 
0.0 0.1923 0 -2.0 1e-06 
0.0 0.1924 0 -2.0 1e-06 
0.0 0.1925 0 -2.0 1e-06 
0.0 0.1926 0 -2.0 1e-06 
0.0 0.1927 0 -2.0 1e-06 
0.0 0.1928 0 -2.0 1e-06 
0.0 0.1929 0 -2.0 1e-06 
0.0 0.193 0 -2.0 1e-06 
0.0 0.1931 0 -2.0 1e-06 
0.0 0.1932 0 -2.0 1e-06 
0.0 0.1933 0 -2.0 1e-06 
0.0 0.1934 0 -2.0 1e-06 
0.0 0.1935 0 -2.0 1e-06 
0.0 0.1936 0 -2.0 1e-06 
0.0 0.1937 0 -2.0 1e-06 
0.0 0.1938 0 -2.0 1e-06 
0.0 0.1939 0 -2.0 1e-06 
0.0 0.194 0 -2.0 1e-06 
0.0 0.1941 0 -2.0 1e-06 
0.0 0.1942 0 -2.0 1e-06 
0.0 0.1943 0 -2.0 1e-06 
0.0 0.1944 0 -2.0 1e-06 
0.0 0.1945 0 -2.0 1e-06 
0.0 0.1946 0 -2.0 1e-06 
0.0 0.1947 0 -2.0 1e-06 
0.0 0.1948 0 -2.0 1e-06 
0.0 0.1949 0 -2.0 1e-06 
0.0 0.195 0 -2.0 1e-06 
0.0 0.1951 0 -2.0 1e-06 
0.0 0.1952 0 -2.0 1e-06 
0.0 0.1953 0 -2.0 1e-06 
0.0 0.1954 0 -2.0 1e-06 
0.0 0.1955 0 -2.0 1e-06 
0.0 0.1956 0 -2.0 1e-06 
0.0 0.1957 0 -2.0 1e-06 
0.0 0.1958 0 -2.0 1e-06 
0.0 0.1959 0 -2.0 1e-06 
0.0 0.196 0 -2.0 1e-06 
0.0 0.1961 0 -2.0 1e-06 
0.0 0.1962 0 -2.0 1e-06 
0.0 0.1963 0 -2.0 1e-06 
0.0 0.1964 0 -2.0 1e-06 
0.0 0.1965 0 -2.0 1e-06 
0.0 0.1966 0 -2.0 1e-06 
0.0 0.1967 0 -2.0 1e-06 
0.0 0.1968 0 -2.0 1e-06 
0.0 0.1969 0 -2.0 1e-06 
0.0 0.197 0 -2.0 1e-06 
0.0 0.1971 0 -2.0 1e-06 
0.0 0.1972 0 -2.0 1e-06 
0.0 0.1973 0 -2.0 1e-06 
0.0 0.1974 0 -2.0 1e-06 
0.0 0.1975 0 -2.0 1e-06 
0.0 0.1976 0 -2.0 1e-06 
0.0 0.1977 0 -2.0 1e-06 
0.0 0.1978 0 -2.0 1e-06 
0.0 0.1979 0 -2.0 1e-06 
0.0 0.198 0 -2.0 1e-06 
0.0 0.1981 0 -2.0 1e-06 
0.0 0.1982 0 -2.0 1e-06 
0.0 0.1983 0 -2.0 1e-06 
0.0 0.1984 0 -2.0 1e-06 
0.0 0.1985 0 -2.0 1e-06 
0.0 0.1986 0 -2.0 1e-06 
0.0 0.1987 0 -2.0 1e-06 
0.0 0.1988 0 -2.0 1e-06 
0.0 0.1989 0 -2.0 1e-06 
0.0 0.199 0 -2.0 1e-06 
0.0 0.1991 0 -2.0 1e-06 
0.0 0.1992 0 -2.0 1e-06 
0.0 0.1993 0 -2.0 1e-06 
0.0 0.1994 0 -2.0 1e-06 
0.0 0.1995 0 -2.0 1e-06 
0.0 0.1996 0 -2.0 1e-06 
0.0 0.1997 0 -2.0 1e-06 
0.0 0.1998 0 -2.0 1e-06 
0.0 0.1999 0 -2.0 1e-06 
0.0 0.2 0 -2.0 1e-06 
0.0 0.2001 0 -2.0 1e-06 
0.0 0.2002 0 -2.0 1e-06 
0.0 0.2003 0 -2.0 1e-06 
0.0 0.2004 0 -2.0 1e-06 
0.0 0.2005 0 -2.0 1e-06 
0.0 0.2006 0 -2.0 1e-06 
0.0 0.2007 0 -2.0 1e-06 
0.0 0.2008 0 -2.0 1e-06 
0.0 0.2009 0 -2.0 1e-06 
0.0 0.201 0 -2.0 1e-06 
0.0 0.2011 0 -2.0 1e-06 
0.0 0.2012 0 -2.0 1e-06 
0.0 0.2013 0 -2.0 1e-06 
0.0 0.2014 0 -2.0 1e-06 
0.0 0.2015 0 -2.0 1e-06 
0.0 0.2016 0 -2.0 1e-06 
0.0 0.2017 0 -2.0 1e-06 
0.0 0.2018 0 -2.0 1e-06 
0.0 0.2019 0 -2.0 1e-06 
0.0 0.202 0 -2.0 1e-06 
0.0 0.2021 0 -2.0 1e-06 
0.0 0.2022 0 -2.0 1e-06 
0.0 0.2023 0 -2.0 1e-06 
0.0 0.2024 0 -2.0 1e-06 
0.0 0.2025 0 -2.0 1e-06 
0.0 0.2026 0 -2.0 1e-06 
0.0 0.2027 0 -2.0 1e-06 
0.0 0.2028 0 -2.0 1e-06 
0.0 0.2029 0 -2.0 1e-06 
0.0 0.203 0 -2.0 1e-06 
0.0 0.2031 0 -2.0 1e-06 
0.0 0.2032 0 -2.0 1e-06 
0.0 0.2033 0 -2.0 1e-06 
0.0 0.2034 0 -2.0 1e-06 
0.0 0.2035 0 -2.0 1e-06 
0.0 0.2036 0 -2.0 1e-06 
0.0 0.2037 0 -2.0 1e-06 
0.0 0.2038 0 -2.0 1e-06 
0.0 0.2039 0 -2.0 1e-06 
0.0 0.204 0 -2.0 1e-06 
0.0 0.2041 0 -2.0 1e-06 
0.0 0.2042 0 -2.0 1e-06 
0.0 0.2043 0 -2.0 1e-06 
0.0 0.2044 0 -2.0 1e-06 
0.0 0.2045 0 -2.0 1e-06 
0.0 0.2046 0 -2.0 1e-06 
0.0 0.2047 0 -2.0 1e-06 
0.0 0.2048 0 -2.0 1e-06 
0.0 0.2049 0 -2.0 1e-06 
0.0 0.205 0 -2.0 1e-06 
0.0 0.2051 0 -2.0 1e-06 
0.0 0.2052 0 -2.0 1e-06 
0.0 0.2053 0 -2.0 1e-06 
0.0 0.2054 0 -2.0 1e-06 
0.0 0.2055 0 -2.0 1e-06 
0.0 0.2056 0 -2.0 1e-06 
0.0 0.2057 0 -2.0 1e-06 
0.0 0.2058 0 -2.0 1e-06 
0.0 0.2059 0 -2.0 1e-06 
0.0 0.206 0 -2.0 1e-06 
0.0 0.2061 0 -2.0 1e-06 
0.0 0.2062 0 -2.0 1e-06 
0.0 0.2063 0 -2.0 1e-06 
0.0 0.2064 0 -2.0 1e-06 
0.0 0.2065 0 -2.0 1e-06 
0.0 0.2066 0 -2.0 1e-06 
0.0 0.2067 0 -2.0 1e-06 
0.0 0.2068 0 -2.0 1e-06 
0.0 0.2069 0 -2.0 1e-06 
0.0 0.207 0 -2.0 1e-06 
0.0 0.2071 0 -2.0 1e-06 
0.0 0.2072 0 -2.0 1e-06 
0.0 0.2073 0 -2.0 1e-06 
0.0 0.2074 0 -2.0 1e-06 
0.0 0.2075 0 -2.0 1e-06 
0.0 0.2076 0 -2.0 1e-06 
0.0 0.2077 0 -2.0 1e-06 
0.0 0.2078 0 -2.0 1e-06 
0.0 0.2079 0 -2.0 1e-06 
0.0 0.208 0 -2.0 1e-06 
0.0 0.2081 0 -2.0 1e-06 
0.0 0.2082 0 -2.0 1e-06 
0.0 0.2083 0 -2.0 1e-06 
0.0 0.2084 0 -2.0 1e-06 
0.0 0.2085 0 -2.0 1e-06 
0.0 0.2086 0 -2.0 1e-06 
0.0 0.2087 0 -2.0 1e-06 
0.0 0.2088 0 -2.0 1e-06 
0.0 0.2089 0 -2.0 1e-06 
0.0 0.209 0 -2.0 1e-06 
0.0 0.2091 0 -2.0 1e-06 
0.0 0.2092 0 -2.0 1e-06 
0.0 0.2093 0 -2.0 1e-06 
0.0 0.2094 0 -2.0 1e-06 
0.0 0.2095 0 -2.0 1e-06 
0.0 0.2096 0 -2.0 1e-06 
0.0 0.2097 0 -2.0 1e-06 
0.0 0.2098 0 -2.0 1e-06 
0.0 0.2099 0 -2.0 1e-06 
0.0 0.21 0 -2.0 1e-06 
0.0 0.2101 0 -2.0 1e-06 
0.0 0.2102 0 -2.0 1e-06 
0.0 0.2103 0 -2.0 1e-06 
0.0 0.2104 0 -2.0 1e-06 
0.0 0.2105 0 -2.0 1e-06 
0.0 0.2106 0 -2.0 1e-06 
0.0 0.2107 0 -2.0 1e-06 
0.0 0.2108 0 -2.0 1e-06 
0.0 0.2109 0 -2.0 1e-06 
0.0 0.211 0 -2.0 1e-06 
0.0 0.2111 0 -2.0 1e-06 
0.0 0.2112 0 -2.0 1e-06 
0.0 0.2113 0 -2.0 1e-06 
0.0 0.2114 0 -2.0 1e-06 
0.0 0.2115 0 -2.0 1e-06 
0.0 0.2116 0 -2.0 1e-06 
0.0 0.2117 0 -2.0 1e-06 
0.0 0.2118 0 -2.0 1e-06 
0.0 0.2119 0 -2.0 1e-06 
0.0 0.212 0 -2.0 1e-06 
0.0 0.2121 0 -2.0 1e-06 
0.0 0.2122 0 -2.0 1e-06 
0.0 0.2123 0 -2.0 1e-06 
0.0 0.2124 0 -2.0 1e-06 
0.0 0.2125 0 -2.0 1e-06 
0.0 0.2126 0 -2.0 1e-06 
0.0 0.2127 0 -2.0 1e-06 
0.0 0.2128 0 -2.0 1e-06 
0.0 0.2129 0 -2.0 1e-06 
0.0 0.213 0 -2.0 1e-06 
0.0 0.2131 0 -2.0 1e-06 
0.0 0.2132 0 -2.0 1e-06 
0.0 0.2133 0 -2.0 1e-06 
0.0 0.2134 0 -2.0 1e-06 
0.0 0.2135 0 -2.0 1e-06 
0.0 0.2136 0 -2.0 1e-06 
0.0 0.2137 0 -2.0 1e-06 
0.0 0.2138 0 -2.0 1e-06 
0.0 0.2139 0 -2.0 1e-06 
0.0 0.214 0 -2.0 1e-06 
0.0 0.2141 0 -2.0 1e-06 
0.0 0.2142 0 -2.0 1e-06 
0.0 0.2143 0 -2.0 1e-06 
0.0 0.2144 0 -2.0 1e-06 
0.0 0.2145 0 -2.0 1e-06 
0.0 0.2146 0 -2.0 1e-06 
0.0 0.2147 0 -2.0 1e-06 
0.0 0.2148 0 -2.0 1e-06 
0.0 0.2149 0 -2.0 1e-06 
0.0 0.215 0 -2.0 1e-06 
0.0 0.2151 0 -2.0 1e-06 
0.0 0.2152 0 -2.0 1e-06 
0.0 0.2153 0 -2.0 1e-06 
0.0 0.2154 0 -2.0 1e-06 
0.0 0.2155 0 -2.0 1e-06 
0.0 0.2156 0 -2.0 1e-06 
0.0 0.2157 0 -2.0 1e-06 
0.0 0.2158 0 -2.0 1e-06 
0.0 0.2159 0 -2.0 1e-06 
0.0 0.216 0 -2.0 1e-06 
0.0 0.2161 0 -2.0 1e-06 
0.0 0.2162 0 -2.0 1e-06 
0.0 0.2163 0 -2.0 1e-06 
0.0 0.2164 0 -2.0 1e-06 
0.0 0.2165 0 -2.0 1e-06 
0.0 0.2166 0 -2.0 1e-06 
0.0 0.2167 0 -2.0 1e-06 
0.0 0.2168 0 -2.0 1e-06 
0.0 0.2169 0 -2.0 1e-06 
0.0 0.217 0 -2.0 1e-06 
0.0 0.2171 0 -2.0 1e-06 
0.0 0.2172 0 -2.0 1e-06 
0.0 0.2173 0 -2.0 1e-06 
0.0 0.2174 0 -2.0 1e-06 
0.0 0.2175 0 -2.0 1e-06 
0.0 0.2176 0 -2.0 1e-06 
0.0 0.2177 0 -2.0 1e-06 
0.0 0.2178 0 -2.0 1e-06 
0.0 0.2179 0 -2.0 1e-06 
0.0 0.218 0 -2.0 1e-06 
0.0 0.2181 0 -2.0 1e-06 
0.0 0.2182 0 -2.0 1e-06 
0.0 0.2183 0 -2.0 1e-06 
0.0 0.2184 0 -2.0 1e-06 
0.0 0.2185 0 -2.0 1e-06 
0.0 0.2186 0 -2.0 1e-06 
0.0 0.2187 0 -2.0 1e-06 
0.0 0.2188 0 -2.0 1e-06 
0.0 0.2189 0 -2.0 1e-06 
0.0 0.219 0 -2.0 1e-06 
0.0 0.2191 0 -2.0 1e-06 
0.0 0.2192 0 -2.0 1e-06 
0.0 0.2193 0 -2.0 1e-06 
0.0 0.2194 0 -2.0 1e-06 
0.0 0.2195 0 -2.0 1e-06 
0.0 0.2196 0 -2.0 1e-06 
0.0 0.2197 0 -2.0 1e-06 
0.0 0.2198 0 -2.0 1e-06 
0.0 0.2199 0 -2.0 1e-06 
0.0 0.22 0 -2.0 1e-06 
0.0 0.2201 0 -2.0 1e-06 
0.0 0.2202 0 -2.0 1e-06 
0.0 0.2203 0 -2.0 1e-06 
0.0 0.2204 0 -2.0 1e-06 
0.0 0.2205 0 -2.0 1e-06 
0.0 0.2206 0 -2.0 1e-06 
0.0 0.2207 0 -2.0 1e-06 
0.0 0.2208 0 -2.0 1e-06 
0.0 0.2209 0 -2.0 1e-06 
0.0 0.221 0 -2.0 1e-06 
0.0 0.2211 0 -2.0 1e-06 
0.0 0.2212 0 -2.0 1e-06 
0.0 0.2213 0 -2.0 1e-06 
0.0 0.2214 0 -2.0 1e-06 
0.0 0.2215 0 -2.0 1e-06 
0.0 0.2216 0 -2.0 1e-06 
0.0 0.2217 0 -2.0 1e-06 
0.0 0.2218 0 -2.0 1e-06 
0.0 0.2219 0 -2.0 1e-06 
0.0 0.222 0 -2.0 1e-06 
0.0 0.2221 0 -2.0 1e-06 
0.0 0.2222 0 -2.0 1e-06 
0.0 0.2223 0 -2.0 1e-06 
0.0 0.2224 0 -2.0 1e-06 
0.0 0.2225 0 -2.0 1e-06 
0.0 0.2226 0 -2.0 1e-06 
0.0 0.2227 0 -2.0 1e-06 
0.0 0.2228 0 -2.0 1e-06 
0.0 0.2229 0 -2.0 1e-06 
0.0 0.223 0 -2.0 1e-06 
0.0 0.2231 0 -2.0 1e-06 
0.0 0.2232 0 -2.0 1e-06 
0.0 0.2233 0 -2.0 1e-06 
0.0 0.2234 0 -2.0 1e-06 
0.0 0.2235 0 -2.0 1e-06 
0.0 0.2236 0 -2.0 1e-06 
0.0 0.2237 0 -2.0 1e-06 
0.0 0.2238 0 -2.0 1e-06 
0.0 0.2239 0 -2.0 1e-06 
0.0 0.224 0 -2.0 1e-06 
0.0 0.2241 0 -2.0 1e-06 
0.0 0.2242 0 -2.0 1e-06 
0.0 0.2243 0 -2.0 1e-06 
0.0 0.2244 0 -2.0 1e-06 
0.0 0.2245 0 -2.0 1e-06 
0.0 0.2246 0 -2.0 1e-06 
0.0 0.2247 0 -2.0 1e-06 
0.0 0.2248 0 -2.0 1e-06 
0.0 0.2249 0 -2.0 1e-06 
0.0 0.225 0 -2.0 1e-06 
0.0 0.2251 0 -2.0 1e-06 
0.0 0.2252 0 -2.0 1e-06 
0.0 0.2253 0 -2.0 1e-06 
0.0 0.2254 0 -2.0 1e-06 
0.0 0.2255 0 -2.0 1e-06 
0.0 0.2256 0 -2.0 1e-06 
0.0 0.2257 0 -2.0 1e-06 
0.0 0.2258 0 -2.0 1e-06 
0.0 0.2259 0 -2.0 1e-06 
0.0 0.226 0 -2.0 1e-06 
0.0 0.2261 0 -2.0 1e-06 
0.0 0.2262 0 -2.0 1e-06 
0.0 0.2263 0 -2.0 1e-06 
0.0 0.2264 0 -2.0 1e-06 
0.0 0.2265 0 -2.0 1e-06 
0.0 0.2266 0 -2.0 1e-06 
0.0 0.2267 0 -2.0 1e-06 
0.0 0.2268 0 -2.0 1e-06 
0.0 0.2269 0 -2.0 1e-06 
0.0 0.227 0 -2.0 1e-06 
0.0 0.2271 0 -2.0 1e-06 
0.0 0.2272 0 -2.0 1e-06 
0.0 0.2273 0 -2.0 1e-06 
0.0 0.2274 0 -2.0 1e-06 
0.0 0.2275 0 -2.0 1e-06 
0.0 0.2276 0 -2.0 1e-06 
0.0 0.2277 0 -2.0 1e-06 
0.0 0.2278 0 -2.0 1e-06 
0.0 0.2279 0 -2.0 1e-06 
0.0 0.228 0 -2.0 1e-06 
0.0 0.2281 0 -2.0 1e-06 
0.0 0.2282 0 -2.0 1e-06 
0.0 0.2283 0 -2.0 1e-06 
0.0 0.2284 0 -2.0 1e-06 
0.0 0.2285 0 -2.0 1e-06 
0.0 0.2286 0 -2.0 1e-06 
0.0 0.2287 0 -2.0 1e-06 
0.0 0.2288 0 -2.0 1e-06 
0.0 0.2289 0 -2.0 1e-06 
0.0 0.229 0 -2.0 1e-06 
0.0 0.2291 0 -2.0 1e-06 
0.0 0.2292 0 -2.0 1e-06 
0.0 0.2293 0 -2.0 1e-06 
0.0 0.2294 0 -2.0 1e-06 
0.0 0.2295 0 -2.0 1e-06 
0.0 0.2296 0 -2.0 1e-06 
0.0 0.2297 0 -2.0 1e-06 
0.0 0.2298 0 -2.0 1e-06 
0.0 0.2299 0 -2.0 1e-06 
0.0 0.23 0 -2.0 1e-06 
0.0 0.2301 0 -2.0 1e-06 
0.0 0.2302 0 -2.0 1e-06 
0.0 0.2303 0 -2.0 1e-06 
0.0 0.2304 0 -2.0 1e-06 
0.0 0.2305 0 -2.0 1e-06 
0.0 0.2306 0 -2.0 1e-06 
0.0 0.2307 0 -2.0 1e-06 
0.0 0.2308 0 -2.0 1e-06 
0.0 0.2309 0 -2.0 1e-06 
0.0 0.231 0 -2.0 1e-06 
0.0 0.2311 0 -2.0 1e-06 
0.0 0.2312 0 -2.0 1e-06 
0.0 0.2313 0 -2.0 1e-06 
0.0 0.2314 0 -2.0 1e-06 
0.0 0.2315 0 -2.0 1e-06 
0.0 0.2316 0 -2.0 1e-06 
0.0 0.2317 0 -2.0 1e-06 
0.0 0.2318 0 -2.0 1e-06 
0.0 0.2319 0 -2.0 1e-06 
0.0 0.232 0 -2.0 1e-06 
0.0 0.2321 0 -2.0 1e-06 
0.0 0.2322 0 -2.0 1e-06 
0.0 0.2323 0 -2.0 1e-06 
0.0 0.2324 0 -2.0 1e-06 
0.0 0.2325 0 -2.0 1e-06 
0.0 0.2326 0 -2.0 1e-06 
0.0 0.2327 0 -2.0 1e-06 
0.0 0.2328 0 -2.0 1e-06 
0.0 0.2329 0 -2.0 1e-06 
0.0 0.233 0 -2.0 1e-06 
0.0 0.2331 0 -2.0 1e-06 
0.0 0.2332 0 -2.0 1e-06 
0.0 0.2333 0 -2.0 1e-06 
0.0 0.2334 0 -2.0 1e-06 
0.0 0.2335 0 -2.0 1e-06 
0.0 0.2336 0 -2.0 1e-06 
0.0 0.2337 0 -2.0 1e-06 
0.0 0.2338 0 -2.0 1e-06 
0.0 0.2339 0 -2.0 1e-06 
0.0 0.234 0 -2.0 1e-06 
0.0 0.2341 0 -2.0 1e-06 
0.0 0.2342 0 -2.0 1e-06 
0.0 0.2343 0 -2.0 1e-06 
0.0 0.2344 0 -2.0 1e-06 
0.0 0.2345 0 -2.0 1e-06 
0.0 0.2346 0 -2.0 1e-06 
0.0 0.2347 0 -2.0 1e-06 
0.0 0.2348 0 -2.0 1e-06 
0.0 0.2349 0 -2.0 1e-06 
0.0 0.235 0 -2.0 1e-06 
0.0 0.2351 0 -2.0 1e-06 
0.0 0.2352 0 -2.0 1e-06 
0.0 0.2353 0 -2.0 1e-06 
0.0 0.2354 0 -2.0 1e-06 
0.0 0.2355 0 -2.0 1e-06 
0.0 0.2356 0 -2.0 1e-06 
0.0 0.2357 0 -2.0 1e-06 
0.0 0.2358 0 -2.0 1e-06 
0.0 0.2359 0 -2.0 1e-06 
0.0 0.236 0 -2.0 1e-06 
0.0 0.2361 0 -2.0 1e-06 
0.0 0.2362 0 -2.0 1e-06 
0.0 0.2363 0 -2.0 1e-06 
0.0 0.2364 0 -2.0 1e-06 
0.0 0.2365 0 -2.0 1e-06 
0.0 0.2366 0 -2.0 1e-06 
0.0 0.2367 0 -2.0 1e-06 
0.0 0.2368 0 -2.0 1e-06 
0.0 0.2369 0 -2.0 1e-06 
0.0 0.237 0 -2.0 1e-06 
0.0 0.2371 0 -2.0 1e-06 
0.0 0.2372 0 -2.0 1e-06 
0.0 0.2373 0 -2.0 1e-06 
0.0 0.2374 0 -2.0 1e-06 
0.0 0.2375 0 -2.0 1e-06 
0.0 0.2376 0 -2.0 1e-06 
0.0 0.2377 0 -2.0 1e-06 
0.0 0.2378 0 -2.0 1e-06 
0.0 0.2379 0 -2.0 1e-06 
0.0 0.238 0 -2.0 1e-06 
0.0 0.2381 0 -2.0 1e-06 
0.0 0.2382 0 -2.0 1e-06 
0.0 0.2383 0 -2.0 1e-06 
0.0 0.2384 0 -2.0 1e-06 
0.0 0.2385 0 -2.0 1e-06 
0.0 0.2386 0 -2.0 1e-06 
0.0 0.2387 0 -2.0 1e-06 
0.0 0.2388 0 -2.0 1e-06 
0.0 0.2389 0 -2.0 1e-06 
0.0 0.239 0 -2.0 1e-06 
0.0 0.2391 0 -2.0 1e-06 
0.0 0.2392 0 -2.0 1e-06 
0.0 0.2393 0 -2.0 1e-06 
0.0 0.2394 0 -2.0 1e-06 
0.0 0.2395 0 -2.0 1e-06 
0.0 0.2396 0 -2.0 1e-06 
0.0 0.2397 0 -2.0 1e-06 
0.0 0.2398 0 -2.0 1e-06 
0.0 0.2399 0 -2.0 1e-06 
0.0 0.24 0 -2.0 1e-06 
0.0 0.2401 0 -2.0 1e-06 
0.0 0.2402 0 -2.0 1e-06 
0.0 0.2403 0 -2.0 1e-06 
0.0 0.2404 0 -2.0 1e-06 
0.0 0.2405 0 -2.0 1e-06 
0.0 0.2406 0 -2.0 1e-06 
0.0 0.2407 0 -2.0 1e-06 
0.0 0.2408 0 -2.0 1e-06 
0.0 0.2409 0 -2.0 1e-06 
0.0 0.241 0 -2.0 1e-06 
0.0 0.2411 0 -2.0 1e-06 
0.0 0.2412 0 -2.0 1e-06 
0.0 0.2413 0 -2.0 1e-06 
0.0 0.2414 0 -2.0 1e-06 
0.0 0.2415 0 -2.0 1e-06 
0.0 0.2416 0 -2.0 1e-06 
0.0 0.2417 0 -2.0 1e-06 
0.0 0.2418 0 -2.0 1e-06 
0.0 0.2419 0 -2.0 1e-06 
0.0 0.242 0 -2.0 1e-06 
0.0 0.2421 0 -2.0 1e-06 
0.0 0.2422 0 -2.0 1e-06 
0.0 0.2423 0 -2.0 1e-06 
0.0 0.2424 0 -2.0 1e-06 
0.0 0.2425 0 -2.0 1e-06 
0.0 0.2426 0 -2.0 1e-06 
0.0 0.2427 0 -2.0 1e-06 
0.0 0.2428 0 -2.0 1e-06 
0.0 0.2429 0 -2.0 1e-06 
0.0 0.243 0 -2.0 1e-06 
0.0 0.2431 0 -2.0 1e-06 
0.0 0.2432 0 -2.0 1e-06 
0.0 0.2433 0 -2.0 1e-06 
0.0 0.2434 0 -2.0 1e-06 
0.0 0.2435 0 -2.0 1e-06 
0.0 0.2436 0 -2.0 1e-06 
0.0 0.2437 0 -2.0 1e-06 
0.0 0.2438 0 -2.0 1e-06 
0.0 0.2439 0 -2.0 1e-06 
0.0 0.244 0 -2.0 1e-06 
0.0 0.2441 0 -2.0 1e-06 
0.0 0.2442 0 -2.0 1e-06 
0.0 0.2443 0 -2.0 1e-06 
0.0 0.2444 0 -2.0 1e-06 
0.0 0.2445 0 -2.0 1e-06 
0.0 0.2446 0 -2.0 1e-06 
0.0 0.2447 0 -2.0 1e-06 
0.0 0.2448 0 -2.0 1e-06 
0.0 0.2449 0 -2.0 1e-06 
0.0 0.245 0 -2.0 1e-06 
0.0 0.2451 0 -2.0 1e-06 
0.0 0.2452 0 -2.0 1e-06 
0.0 0.2453 0 -2.0 1e-06 
0.0 0.2454 0 -2.0 1e-06 
0.0 0.2455 0 -2.0 1e-06 
0.0 0.2456 0 -2.0 1e-06 
0.0 0.2457 0 -2.0 1e-06 
0.0 0.2458 0 -2.0 1e-06 
0.0 0.2459 0 -2.0 1e-06 
0.0 0.246 0 -2.0 1e-06 
0.0 0.2461 0 -2.0 1e-06 
0.0 0.2462 0 -2.0 1e-06 
0.0 0.2463 0 -2.0 1e-06 
0.0 0.2464 0 -2.0 1e-06 
0.0 0.2465 0 -2.0 1e-06 
0.0 0.2466 0 -2.0 1e-06 
0.0 0.2467 0 -2.0 1e-06 
0.0 0.2468 0 -2.0 1e-06 
0.0 0.2469 0 -2.0 1e-06 
0.0 0.247 0 -2.0 1e-06 
0.0 0.2471 0 -2.0 1e-06 
0.0 0.2472 0 -2.0 1e-06 
0.0 0.2473 0 -2.0 1e-06 
0.0 0.2474 0 -2.0 1e-06 
0.0 0.2475 0 -2.0 1e-06 
0.0 0.2476 0 -2.0 1e-06 
0.0 0.2477 0 -2.0 1e-06 
0.0 0.2478 0 -2.0 1e-06 
0.0 0.2479 0 -2.0 1e-06 
0.0 0.248 0 -2.0 1e-06 
0.0 0.2481 0 -2.0 1e-06 
0.0 0.2482 0 -2.0 1e-06 
0.0 0.2483 0 -2.0 1e-06 
0.0 0.2484 0 -2.0 1e-06 
0.0 0.2485 0 -2.0 1e-06 
0.0 0.2486 0 -2.0 1e-06 
0.0 0.2487 0 -2.0 1e-06 
0.0 0.2488 0 -2.0 1e-06 
0.0 0.2489 0 -2.0 1e-06 
0.0 0.249 0 -2.0 1e-06 
0.0 0.2491 0 -2.0 1e-06 
0.0 0.2492 0 -2.0 1e-06 
0.0 0.2493 0 -2.0 1e-06 
0.0 0.2494 0 -2.0 1e-06 
0.0 0.2495 0 -2.0 1e-06 
0.0 0.2496 0 -2.0 1e-06 
0.0 0.2497 0 -2.0 1e-06 
0.0 0.2498 0 -2.0 1e-06 
0.0 0.2499 0 -2.0 1e-06 
0.0 0.25 0 -2.0 1e-06 
0.0 0.2501 0 -2.0 1e-06 
0.0 0.2502 0 -2.0 1e-06 
0.0 0.2503 0 -2.0 1e-06 
0.0 0.2504 0 -2.0 1e-06 
0.0 0.2505 0 -2.0 1e-06 
0.0 0.2506 0 -2.0 1e-06 
0.0 0.2507 0 -2.0 1e-06 
0.0 0.2508 0 -2.0 1e-06 
0.0 0.2509 0 -2.0 1e-06 
0.0 0.251 0 -2.0 1e-06 
0.0 0.2511 0 -2.0 1e-06 
0.0 0.2512 0 -2.0 1e-06 
0.0 0.2513 0 -2.0 1e-06 
0.0 0.2514 0 -2.0 1e-06 
0.0 0.2515 0 -2.0 1e-06 
0.0 0.2516 0 -2.0 1e-06 
0.0 0.2517 0 -2.0 1e-06 
0.0 0.2518 0 -2.0 1e-06 
0.0 0.2519 0 -2.0 1e-06 
0.0 0.252 0 -2.0 1e-06 
0.0 0.2521 0 -2.0 1e-06 
0.0 0.2522 0 -2.0 1e-06 
0.0 0.2523 0 -2.0 1e-06 
0.0 0.2524 0 -2.0 1e-06 
0.0 0.2525 0 -2.0 1e-06 
0.0 0.2526 0 -2.0 1e-06 
0.0 0.2527 0 -2.0 1e-06 
0.0 0.2528 0 -2.0 1e-06 
0.0 0.2529 0 -2.0 1e-06 
0.0 0.253 0 -2.0 1e-06 
0.0 0.2531 0 -2.0 1e-06 
0.0 0.2532 0 -2.0 1e-06 
0.0 0.2533 0 -2.0 1e-06 
0.0 0.2534 0 -2.0 1e-06 
0.0 0.2535 0 -2.0 1e-06 
0.0 0.2536 0 -2.0 1e-06 
0.0 0.2537 0 -2.0 1e-06 
0.0 0.2538 0 -2.0 1e-06 
0.0 0.2539 0 -2.0 1e-06 
0.0 0.254 0 -2.0 1e-06 
0.0 0.2541 0 -2.0 1e-06 
0.0 0.2542 0 -2.0 1e-06 
0.0 0.2543 0 -2.0 1e-06 
0.0 0.2544 0 -2.0 1e-06 
0.0 0.2545 0 -2.0 1e-06 
0.0 0.2546 0 -2.0 1e-06 
0.0 0.2547 0 -2.0 1e-06 
0.0 0.2548 0 -2.0 1e-06 
0.0 0.2549 0 -2.0 1e-06 
0.0 0.255 0 -2.0 1e-06 
0.0 0.2551 0 -2.0 1e-06 
0.0 0.2552 0 -2.0 1e-06 
0.0 0.2553 0 -2.0 1e-06 
0.0 0.2554 0 -2.0 1e-06 
0.0 0.2555 0 -2.0 1e-06 
0.0 0.2556 0 -2.0 1e-06 
0.0 0.2557 0 -2.0 1e-06 
0.0 0.2558 0 -2.0 1e-06 
0.0 0.2559 0 -2.0 1e-06 
0.0 0.256 0 -2.0 1e-06 
0.0 0.2561 0 -2.0 1e-06 
0.0 0.2562 0 -2.0 1e-06 
0.0 0.2563 0 -2.0 1e-06 
0.0 0.2564 0 -2.0 1e-06 
0.0 0.2565 0 -2.0 1e-06 
0.0 0.2566 0 -2.0 1e-06 
0.0 0.2567 0 -2.0 1e-06 
0.0 0.2568 0 -2.0 1e-06 
0.0 0.2569 0 -2.0 1e-06 
0.0 0.257 0 -2.0 1e-06 
0.0 0.2571 0 -2.0 1e-06 
0.0 0.2572 0 -2.0 1e-06 
0.0 0.2573 0 -2.0 1e-06 
0.0 0.2574 0 -2.0 1e-06 
0.0 0.2575 0 -2.0 1e-06 
0.0 0.2576 0 -2.0 1e-06 
0.0 0.2577 0 -2.0 1e-06 
0.0 0.2578 0 -2.0 1e-06 
0.0 0.2579 0 -2.0 1e-06 
0.0 0.258 0 -2.0 1e-06 
0.0 0.2581 0 -2.0 1e-06 
0.0 0.2582 0 -2.0 1e-06 
0.0 0.2583 0 -2.0 1e-06 
0.0 0.2584 0 -2.0 1e-06 
0.0 0.2585 0 -2.0 1e-06 
0.0 0.2586 0 -2.0 1e-06 
0.0 0.2587 0 -2.0 1e-06 
0.0 0.2588 0 -2.0 1e-06 
0.0 0.2589 0 -2.0 1e-06 
0.0 0.259 0 -2.0 1e-06 
0.0 0.2591 0 -2.0 1e-06 
0.0 0.2592 0 -2.0 1e-06 
0.0 0.2593 0 -2.0 1e-06 
0.0 0.2594 0 -2.0 1e-06 
0.0 0.2595 0 -2.0 1e-06 
0.0 0.2596 0 -2.0 1e-06 
0.0 0.2597 0 -2.0 1e-06 
0.0 0.2598 0 -2.0 1e-06 
0.0 0.2599 0 -2.0 1e-06 
0.0 0.26 0 -2.0 1e-06 
0.0 0.2601 0 -2.0 1e-06 
0.0 0.2602 0 -2.0 1e-06 
0.0 0.2603 0 -2.0 1e-06 
0.0 0.2604 0 -2.0 1e-06 
0.0 0.2605 0 -2.0 1e-06 
0.0 0.2606 0 -2.0 1e-06 
0.0 0.2607 0 -2.0 1e-06 
0.0 0.2608 0 -2.0 1e-06 
0.0 0.2609 0 -2.0 1e-06 
0.0 0.261 0 -2.0 1e-06 
0.0 0.2611 0 -2.0 1e-06 
0.0 0.2612 0 -2.0 1e-06 
0.0 0.2613 0 -2.0 1e-06 
0.0 0.2614 0 -2.0 1e-06 
0.0 0.2615 0 -2.0 1e-06 
0.0 0.2616 0 -2.0 1e-06 
0.0 0.2617 0 -2.0 1e-06 
0.0 0.2618 0 -2.0 1e-06 
0.0 0.2619 0 -2.0 1e-06 
0.0 0.262 0 -2.0 1e-06 
0.0 0.2621 0 -2.0 1e-06 
0.0 0.2622 0 -2.0 1e-06 
0.0 0.2623 0 -2.0 1e-06 
0.0 0.2624 0 -2.0 1e-06 
0.0 0.2625 0 -2.0 1e-06 
0.0 0.2626 0 -2.0 1e-06 
0.0 0.2627 0 -2.0 1e-06 
0.0 0.2628 0 -2.0 1e-06 
0.0 0.2629 0 -2.0 1e-06 
0.0 0.263 0 -2.0 1e-06 
0.0 0.2631 0 -2.0 1e-06 
0.0 0.2632 0 -2.0 1e-06 
0.0 0.2633 0 -2.0 1e-06 
0.0 0.2634 0 -2.0 1e-06 
0.0 0.2635 0 -2.0 1e-06 
0.0 0.2636 0 -2.0 1e-06 
0.0 0.2637 0 -2.0 1e-06 
0.0 0.2638 0 -2.0 1e-06 
0.0 0.2639 0 -2.0 1e-06 
0.0 0.264 0 -2.0 1e-06 
0.0 0.2641 0 -2.0 1e-06 
0.0 0.2642 0 -2.0 1e-06 
0.0 0.2643 0 -2.0 1e-06 
0.0 0.2644 0 -2.0 1e-06 
0.0 0.2645 0 -2.0 1e-06 
0.0 0.2646 0 -2.0 1e-06 
0.0 0.2647 0 -2.0 1e-06 
0.0 0.2648 0 -2.0 1e-06 
0.0 0.2649 0 -2.0 1e-06 
0.0 0.265 0 -2.0 1e-06 
0.0 0.2651 0 -2.0 1e-06 
0.0 0.2652 0 -2.0 1e-06 
0.0 0.2653 0 -2.0 1e-06 
0.0 0.2654 0 -2.0 1e-06 
0.0 0.2655 0 -2.0 1e-06 
0.0 0.2656 0 -2.0 1e-06 
0.0 0.2657 0 -2.0 1e-06 
0.0 0.2658 0 -2.0 1e-06 
0.0 0.2659 0 -2.0 1e-06 
0.0 0.266 0 -2.0 1e-06 
0.0 0.2661 0 -2.0 1e-06 
0.0 0.2662 0 -2.0 1e-06 
0.0 0.2663 0 -2.0 1e-06 
0.0 0.2664 0 -2.0 1e-06 
0.0 0.2665 0 -2.0 1e-06 
0.0 0.2666 0 -2.0 1e-06 
0.0 0.2667 0 -2.0 1e-06 
0.0 0.2668 0 -2.0 1e-06 
0.0 0.2669 0 -2.0 1e-06 
0.0 0.267 0 -2.0 1e-06 
0.0 0.2671 0 -2.0 1e-06 
0.0 0.2672 0 -2.0 1e-06 
0.0 0.2673 0 -2.0 1e-06 
0.0 0.2674 0 -2.0 1e-06 
0.0 0.2675 0 -2.0 1e-06 
0.0 0.2676 0 -2.0 1e-06 
0.0 0.2677 0 -2.0 1e-06 
0.0 0.2678 0 -2.0 1e-06 
0.0 0.2679 0 -2.0 1e-06 
0.0 0.268 0 -2.0 1e-06 
0.0 0.2681 0 -2.0 1e-06 
0.0 0.2682 0 -2.0 1e-06 
0.0 0.2683 0 -2.0 1e-06 
0.0 0.2684 0 -2.0 1e-06 
0.0 0.2685 0 -2.0 1e-06 
0.0 0.2686 0 -2.0 1e-06 
0.0 0.2687 0 -2.0 1e-06 
0.0 0.2688 0 -2.0 1e-06 
0.0 0.2689 0 -2.0 1e-06 
0.0 0.269 0 -2.0 1e-06 
0.0 0.2691 0 -2.0 1e-06 
0.0 0.2692 0 -2.0 1e-06 
0.0 0.2693 0 -2.0 1e-06 
0.0 0.2694 0 -2.0 1e-06 
0.0 0.2695 0 -2.0 1e-06 
0.0 0.2696 0 -2.0 1e-06 
0.0 0.2697 0 -2.0 1e-06 
0.0 0.2698 0 -2.0 1e-06 
0.0 0.2699 0 -2.0 1e-06 
0.0 0.27 0 -2.0 1e-06 
0.0 0.2701 0 -2.0 1e-06 
0.0 0.2702 0 -2.0 1e-06 
0.0 0.2703 0 -2.0 1e-06 
0.0 0.2704 0 -2.0 1e-06 
0.0 0.2705 0 -2.0 1e-06 
0.0 0.2706 0 -2.0 1e-06 
0.0 0.2707 0 -2.0 1e-06 
0.0 0.2708 0 -2.0 1e-06 
0.0 0.2709 0 -2.0 1e-06 
0.0 0.271 0 -2.0 1e-06 
0.0 0.2711 0 -2.0 1e-06 
0.0 0.2712 0 -2.0 1e-06 
0.0 0.2713 0 -2.0 1e-06 
0.0 0.2714 0 -2.0 1e-06 
0.0 0.2715 0 -2.0 1e-06 
0.0 0.2716 0 -2.0 1e-06 
0.0 0.2717 0 -2.0 1e-06 
0.0 0.2718 0 -2.0 1e-06 
0.0 0.2719 0 -2.0 1e-06 
0.0 0.272 0 -2.0 1e-06 
0.0 0.2721 0 -2.0 1e-06 
0.0 0.2722 0 -2.0 1e-06 
0.0 0.2723 0 -2.0 1e-06 
0.0 0.2724 0 -2.0 1e-06 
0.0 0.2725 0 -2.0 1e-06 
0.0 0.2726 0 -2.0 1e-06 
0.0 0.2727 0 -2.0 1e-06 
0.0 0.2728 0 -2.0 1e-06 
0.0 0.2729 0 -2.0 1e-06 
0.0 0.273 0 -2.0 1e-06 
0.0 0.2731 0 -2.0 1e-06 
0.0 0.2732 0 -2.0 1e-06 
0.0 0.2733 0 -2.0 1e-06 
0.0 0.2734 0 -2.0 1e-06 
0.0 0.2735 0 -2.0 1e-06 
0.0 0.2736 0 -2.0 1e-06 
0.0 0.2737 0 -2.0 1e-06 
0.0 0.2738 0 -2.0 1e-06 
0.0 0.2739 0 -2.0 1e-06 
0.0 0.274 0 -2.0 1e-06 
0.0 0.2741 0 -2.0 1e-06 
0.0 0.2742 0 -2.0 1e-06 
0.0 0.2743 0 -2.0 1e-06 
0.0 0.2744 0 -2.0 1e-06 
0.0 0.2745 0 -2.0 1e-06 
0.0 0.2746 0 -2.0 1e-06 
0.0 0.2747 0 -2.0 1e-06 
0.0 0.2748 0 -2.0 1e-06 
0.0 0.2749 0 -2.0 1e-06 
0.0 0.275 0 -2.0 1e-06 
0.0 0.2751 0 -2.0 1e-06 
0.0 0.2752 0 -2.0 1e-06 
0.0 0.2753 0 -2.0 1e-06 
0.0 0.2754 0 -2.0 1e-06 
0.0 0.2755 0 -2.0 1e-06 
0.0 0.2756 0 -2.0 1e-06 
0.0 0.2757 0 -2.0 1e-06 
0.0 0.2758 0 -2.0 1e-06 
0.0 0.2759 0 -2.0 1e-06 
0.0 0.276 0 -2.0 1e-06 
0.0 0.2761 0 -2.0 1e-06 
0.0 0.2762 0 -2.0 1e-06 
0.0 0.2763 0 -2.0 1e-06 
0.0 0.2764 0 -2.0 1e-06 
0.0 0.2765 0 -2.0 1e-06 
0.0 0.2766 0 -2.0 1e-06 
0.0 0.2767 0 -2.0 1e-06 
0.0 0.2768 0 -2.0 1e-06 
0.0 0.2769 0 -2.0 1e-06 
0.0 0.277 0 -2.0 1e-06 
0.0 0.2771 0 -2.0 1e-06 
0.0 0.2772 0 -2.0 1e-06 
0.0 0.2773 0 -2.0 1e-06 
0.0 0.2774 0 -2.0 1e-06 
0.0 0.2775 0 -2.0 1e-06 
0.0 0.2776 0 -2.0 1e-06 
0.0 0.2777 0 -2.0 1e-06 
0.0 0.2778 0 -2.0 1e-06 
0.0 0.2779 0 -2.0 1e-06 
0.0 0.278 0 -2.0 1e-06 
0.0 0.2781 0 -2.0 1e-06 
0.0 0.2782 0 -2.0 1e-06 
0.0 0.2783 0 -2.0 1e-06 
0.0 0.2784 0 -2.0 1e-06 
0.0 0.2785 0 -2.0 1e-06 
0.0 0.2786 0 -2.0 1e-06 
0.0 0.2787 0 -2.0 1e-06 
0.0 0.2788 0 -2.0 1e-06 
0.0 0.2789 0 -2.0 1e-06 
0.0 0.279 0 -2.0 1e-06 
0.0 0.2791 0 -2.0 1e-06 
0.0 0.2792 0 -2.0 1e-06 
0.0 0.2793 0 -2.0 1e-06 
0.0 0.2794 0 -2.0 1e-06 
0.0 0.2795 0 -2.0 1e-06 
0.0 0.2796 0 -2.0 1e-06 
0.0 0.2797 0 -2.0 1e-06 
0.0 0.2798 0 -2.0 1e-06 
0.0 0.2799 0 -2.0 1e-06 
0.0 0.28 0 -2.0 1e-06 
0.0 0.2801 0 -2.0 1e-06 
0.0 0.2802 0 -2.0 1e-06 
0.0 0.2803 0 -2.0 1e-06 
0.0 0.2804 0 -2.0 1e-06 
0.0 0.2805 0 -2.0 1e-06 
0.0 0.2806 0 -2.0 1e-06 
0.0 0.2807 0 -2.0 1e-06 
0.0 0.2808 0 -2.0 1e-06 
0.0 0.2809 0 -2.0 1e-06 
0.0 0.281 0 -2.0 1e-06 
0.0 0.2811 0 -2.0 1e-06 
0.0 0.2812 0 -2.0 1e-06 
0.0 0.2813 0 -2.0 1e-06 
0.0 0.2814 0 -2.0 1e-06 
0.0 0.2815 0 -2.0 1e-06 
0.0 0.2816 0 -2.0 1e-06 
0.0 0.2817 0 -2.0 1e-06 
0.0 0.2818 0 -2.0 1e-06 
0.0 0.2819 0 -2.0 1e-06 
0.0 0.282 0 -2.0 1e-06 
0.0 0.2821 0 -2.0 1e-06 
0.0 0.2822 0 -2.0 1e-06 
0.0 0.2823 0 -2.0 1e-06 
0.0 0.2824 0 -2.0 1e-06 
0.0 0.2825 0 -2.0 1e-06 
0.0 0.2826 0 -2.0 1e-06 
0.0 0.2827 0 -2.0 1e-06 
0.0 0.2828 0 -2.0 1e-06 
0.0 0.2829 0 -2.0 1e-06 
0.0 0.283 0 -2.0 1e-06 
0.0 0.2831 0 -2.0 1e-06 
0.0 0.2832 0 -2.0 1e-06 
0.0 0.2833 0 -2.0 1e-06 
0.0 0.2834 0 -2.0 1e-06 
0.0 0.2835 0 -2.0 1e-06 
0.0 0.2836 0 -2.0 1e-06 
0.0 0.2837 0 -2.0 1e-06 
0.0 0.2838 0 -2.0 1e-06 
0.0 0.2839 0 -2.0 1e-06 
0.0 0.284 0 -2.0 1e-06 
0.0 0.2841 0 -2.0 1e-06 
0.0 0.2842 0 -2.0 1e-06 
0.0 0.2843 0 -2.0 1e-06 
0.0 0.2844 0 -2.0 1e-06 
0.0 0.2845 0 -2.0 1e-06 
0.0 0.2846 0 -2.0 1e-06 
0.0 0.2847 0 -2.0 1e-06 
0.0 0.2848 0 -2.0 1e-06 
0.0 0.2849 0 -2.0 1e-06 
0.0 0.285 0 -2.0 1e-06 
0.0 0.2851 0 -2.0 1e-06 
0.0 0.2852 0 -2.0 1e-06 
0.0 0.2853 0 -2.0 1e-06 
0.0 0.2854 0 -2.0 1e-06 
0.0 0.2855 0 -2.0 1e-06 
0.0 0.2856 0 -2.0 1e-06 
0.0 0.2857 0 -2.0 1e-06 
0.0 0.2858 0 -2.0 1e-06 
0.0 0.2859 0 -2.0 1e-06 
0.0 0.286 0 -2.0 1e-06 
0.0 0.2861 0 -2.0 1e-06 
0.0 0.2862 0 -2.0 1e-06 
0.0 0.2863 0 -2.0 1e-06 
0.0 0.2864 0 -2.0 1e-06 
0.0 0.2865 0 -2.0 1e-06 
0.0 0.2866 0 -2.0 1e-06 
0.0 0.2867 0 -2.0 1e-06 
0.0 0.2868 0 -2.0 1e-06 
0.0 0.2869 0 -2.0 1e-06 
0.0 0.287 0 -2.0 1e-06 
0.0 0.2871 0 -2.0 1e-06 
0.0 0.2872 0 -2.0 1e-06 
0.0 0.2873 0 -2.0 1e-06 
0.0 0.2874 0 -2.0 1e-06 
0.0 0.2875 0 -2.0 1e-06 
0.0 0.2876 0 -2.0 1e-06 
0.0 0.2877 0 -2.0 1e-06 
0.0 0.2878 0 -2.0 1e-06 
0.0 0.2879 0 -2.0 1e-06 
0.0 0.288 0 -2.0 1e-06 
0.0 0.2881 0 -2.0 1e-06 
0.0 0.2882 0 -2.0 1e-06 
0.0 0.2883 0 -2.0 1e-06 
0.0 0.2884 0 -2.0 1e-06 
0.0 0.2885 0 -2.0 1e-06 
0.0 0.2886 0 -2.0 1e-06 
0.0 0.2887 0 -2.0 1e-06 
0.0 0.2888 0 -2.0 1e-06 
0.0 0.2889 0 -2.0 1e-06 
0.0 0.289 0 -2.0 1e-06 
0.0 0.2891 0 -2.0 1e-06 
0.0 0.2892 0 -2.0 1e-06 
0.0 0.2893 0 -2.0 1e-06 
0.0 0.2894 0 -2.0 1e-06 
0.0 0.2895 0 -2.0 1e-06 
0.0 0.2896 0 -2.0 1e-06 
0.0 0.2897 0 -2.0 1e-06 
0.0 0.2898 0 -2.0 1e-06 
0.0 0.2899 0 -2.0 1e-06 
0.0 0.29 0 -2.0 1e-06 
0.0 0.2901 0 -2.0 1e-06 
0.0 0.2902 0 -2.0 1e-06 
0.0 0.2903 0 -2.0 1e-06 
0.0 0.2904 0 -2.0 1e-06 
0.0 0.2905 0 -2.0 1e-06 
0.0 0.2906 0 -2.0 1e-06 
0.0 0.2907 0 -2.0 1e-06 
0.0 0.2908 0 -2.0 1e-06 
0.0 0.2909 0 -2.0 1e-06 
0.0 0.291 0 -2.0 1e-06 
0.0 0.2911 0 -2.0 1e-06 
0.0 0.2912 0 -2.0 1e-06 
0.0 0.2913 0 -2.0 1e-06 
0.0 0.2914 0 -2.0 1e-06 
0.0 0.2915 0 -2.0 1e-06 
0.0 0.2916 0 -2.0 1e-06 
0.0 0.2917 0 -2.0 1e-06 
0.0 0.2918 0 -2.0 1e-06 
0.0 0.2919 0 -2.0 1e-06 
0.0 0.292 0 -2.0 1e-06 
0.0 0.2921 0 -2.0 1e-06 
0.0 0.2922 0 -2.0 1e-06 
0.0 0.2923 0 -2.0 1e-06 
0.0 0.2924 0 -2.0 1e-06 
0.0 0.2925 0 -2.0 1e-06 
0.0 0.2926 0 -2.0 1e-06 
0.0 0.2927 0 -2.0 1e-06 
0.0 0.2928 0 -2.0 1e-06 
0.0 0.2929 0 -2.0 1e-06 
0.0 0.293 0 -2.0 1e-06 
0.0 0.2931 0 -2.0 1e-06 
0.0 0.2932 0 -2.0 1e-06 
0.0 0.2933 0 -2.0 1e-06 
0.0 0.2934 0 -2.0 1e-06 
0.0 0.2935 0 -2.0 1e-06 
0.0 0.2936 0 -2.0 1e-06 
0.0 0.2937 0 -2.0 1e-06 
0.0 0.2938 0 -2.0 1e-06 
0.0 0.2939 0 -2.0 1e-06 
0.0 0.294 0 -2.0 1e-06 
0.0 0.2941 0 -2.0 1e-06 
0.0 0.2942 0 -2.0 1e-06 
0.0 0.2943 0 -2.0 1e-06 
0.0 0.2944 0 -2.0 1e-06 
0.0 0.2945 0 -2.0 1e-06 
0.0 0.2946 0 -2.0 1e-06 
0.0 0.2947 0 -2.0 1e-06 
0.0 0.2948 0 -2.0 1e-06 
0.0 0.2949 0 -2.0 1e-06 
0.0 0.295 0 -2.0 1e-06 
0.0 0.2951 0 -2.0 1e-06 
0.0 0.2952 0 -2.0 1e-06 
0.0 0.2953 0 -2.0 1e-06 
0.0 0.2954 0 -2.0 1e-06 
0.0 0.2955 0 -2.0 1e-06 
0.0 0.2956 0 -2.0 1e-06 
0.0 0.2957 0 -2.0 1e-06 
0.0 0.2958 0 -2.0 1e-06 
0.0 0.2959 0 -2.0 1e-06 
0.0 0.296 0 -2.0 1e-06 
0.0 0.2961 0 -2.0 1e-06 
0.0 0.2962 0 -2.0 1e-06 
0.0 0.2963 0 -2.0 1e-06 
0.0 0.2964 0 -2.0 1e-06 
0.0 0.2965 0 -2.0 1e-06 
0.0 0.2966 0 -2.0 1e-06 
0.0 0.2967 0 -2.0 1e-06 
0.0 0.2968 0 -2.0 1e-06 
0.0 0.2969 0 -2.0 1e-06 
0.0 0.297 0 -2.0 1e-06 
0.0 0.2971 0 -2.0 1e-06 
0.0 0.2972 0 -2.0 1e-06 
0.0 0.2973 0 -2.0 1e-06 
0.0 0.2974 0 -2.0 1e-06 
0.0 0.2975 0 -2.0 1e-06 
0.0 0.2976 0 -2.0 1e-06 
0.0 0.2977 0 -2.0 1e-06 
0.0 0.2978 0 -2.0 1e-06 
0.0 0.2979 0 -2.0 1e-06 
0.0 0.298 0 -2.0 1e-06 
0.0 0.2981 0 -2.0 1e-06 
0.0 0.2982 0 -2.0 1e-06 
0.0 0.2983 0 -2.0 1e-06 
0.0 0.2984 0 -2.0 1e-06 
0.0 0.2985 0 -2.0 1e-06 
0.0 0.2986 0 -2.0 1e-06 
0.0 0.2987 0 -2.0 1e-06 
0.0 0.2988 0 -2.0 1e-06 
0.0 0.2989 0 -2.0 1e-06 
0.0 0.299 0 -2.0 1e-06 
0.0 0.2991 0 -2.0 1e-06 
0.0 0.2992 0 -2.0 1e-06 
0.0 0.2993 0 -2.0 1e-06 
0.0 0.2994 0 -2.0 1e-06 
0.0 0.2995 0 -2.0 1e-06 
0.0 0.2996 0 -2.0 1e-06 
0.0 0.2997 0 -2.0 1e-06 
0.0 0.2998 0 -2.0 1e-06 
0.0 0.2999 0 -2.0 1e-06 
0.0 0.3 0 -2.0 1e-06 
0.0 0.3001 0 -2.0 1e-06 
0.0 0.3002 0 -2.0 1e-06 
0.0 0.3003 0 -2.0 1e-06 
0.0 0.3004 0 -2.0 1e-06 
0.0 0.3005 0 -2.0 1e-06 
0.0 0.3006 0 -2.0 1e-06 
0.0 0.3007 0 -2.0 1e-06 
0.0 0.3008 0 -2.0 1e-06 
0.0 0.3009 0 -2.0 1e-06 
0.0 0.301 0 -2.0 1e-06 
0.0 0.3011 0 -2.0 1e-06 
0.0 0.3012 0 -2.0 1e-06 
0.0 0.3013 0 -2.0 1e-06 
0.0 0.3014 0 -2.0 1e-06 
0.0 0.3015 0 -2.0 1e-06 
0.0 0.3016 0 -2.0 1e-06 
0.0 0.3017 0 -2.0 1e-06 
0.0 0.3018 0 -2.0 1e-06 
0.0 0.3019 0 -2.0 1e-06 
0.0 0.302 0 -2.0 1e-06 
0.0 0.3021 0 -2.0 1e-06 
0.0 0.3022 0 -2.0 1e-06 
0.0 0.3023 0 -2.0 1e-06 
0.0 0.3024 0 -2.0 1e-06 
0.0 0.3025 0 -2.0 1e-06 
0.0 0.3026 0 -2.0 1e-06 
0.0 0.3027 0 -2.0 1e-06 
0.0 0.3028 0 -2.0 1e-06 
0.0 0.3029 0 -2.0 1e-06 
0.0 0.303 0 -2.0 1e-06 
0.0 0.3031 0 -2.0 1e-06 
0.0 0.3032 0 -2.0 1e-06 
0.0 0.3033 0 -2.0 1e-06 
0.0 0.3034 0 -2.0 1e-06 
0.0 0.3035 0 -2.0 1e-06 
0.0 0.3036 0 -2.0 1e-06 
0.0 0.3037 0 -2.0 1e-06 
0.0 0.3038 0 -2.0 1e-06 
0.0 0.3039 0 -2.0 1e-06 
0.0 0.304 0 -2.0 1e-06 
0.0 0.3041 0 -2.0 1e-06 
0.0 0.3042 0 -2.0 1e-06 
0.0 0.3043 0 -2.0 1e-06 
0.0 0.3044 0 -2.0 1e-06 
0.0 0.3045 0 -2.0 1e-06 
0.0 0.3046 0 -2.0 1e-06 
0.0 0.3047 0 -2.0 1e-06 
0.0 0.3048 0 -2.0 1e-06 
0.0 0.3049 0 -2.0 1e-06 
0.0 0.305 0 -2.0 1e-06 
0.0 0.3051 0 -2.0 1e-06 
0.0 0.3052 0 -2.0 1e-06 
0.0 0.3053 0 -2.0 1e-06 
0.0 0.3054 0 -2.0 1e-06 
0.0 0.3055 0 -2.0 1e-06 
0.0 0.3056 0 -2.0 1e-06 
0.0 0.3057 0 -2.0 1e-06 
0.0 0.3058 0 -2.0 1e-06 
0.0 0.3059 0 -2.0 1e-06 
0.0 0.306 0 -2.0 1e-06 
0.0 0.3061 0 -2.0 1e-06 
0.0 0.3062 0 -2.0 1e-06 
0.0 0.3063 0 -2.0 1e-06 
0.0 0.3064 0 -2.0 1e-06 
0.0 0.3065 0 -2.0 1e-06 
0.0 0.3066 0 -2.0 1e-06 
0.0 0.3067 0 -2.0 1e-06 
0.0 0.3068 0 -2.0 1e-06 
0.0 0.3069 0 -2.0 1e-06 
0.0 0.307 0 -2.0 1e-06 
0.0 0.3071 0 -2.0 1e-06 
0.0 0.3072 0 -2.0 1e-06 
0.0 0.3073 0 -2.0 1e-06 
0.0 0.3074 0 -2.0 1e-06 
0.0 0.3075 0 -2.0 1e-06 
0.0 0.3076 0 -2.0 1e-06 
0.0 0.3077 0 -2.0 1e-06 
0.0 0.3078 0 -2.0 1e-06 
0.0 0.3079 0 -2.0 1e-06 
0.0 0.308 0 -2.0 1e-06 
0.0 0.3081 0 -2.0 1e-06 
0.0 0.3082 0 -2.0 1e-06 
0.0 0.3083 0 -2.0 1e-06 
0.0 0.3084 0 -2.0 1e-06 
0.0 0.3085 0 -2.0 1e-06 
0.0 0.3086 0 -2.0 1e-06 
0.0 0.3087 0 -2.0 1e-06 
0.0 0.3088 0 -2.0 1e-06 
0.0 0.3089 0 -2.0 1e-06 
0.0 0.309 0 -2.0 1e-06 
0.0 0.3091 0 -2.0 1e-06 
0.0 0.3092 0 -2.0 1e-06 
0.0 0.3093 0 -2.0 1e-06 
0.0 0.3094 0 -2.0 1e-06 
0.0 0.3095 0 -2.0 1e-06 
0.0 0.3096 0 -2.0 1e-06 
0.0 0.3097 0 -2.0 1e-06 
0.0 0.3098 0 -2.0 1e-06 
0.0 0.3099 0 -2.0 1e-06 
0.0 0.31 0 -2.0 1e-06 
0.0 0.3101 0 -2.0 1e-06 
0.0 0.3102 0 -2.0 1e-06 
0.0 0.3103 0 -2.0 1e-06 
0.0 0.3104 0 -2.0 1e-06 
0.0 0.3105 0 -2.0 1e-06 
0.0 0.3106 0 -2.0 1e-06 
0.0 0.3107 0 -2.0 1e-06 
0.0 0.3108 0 -2.0 1e-06 
0.0 0.3109 0 -2.0 1e-06 
0.0 0.311 0 -2.0 1e-06 
0.0 0.3111 0 -2.0 1e-06 
0.0 0.3112 0 -2.0 1e-06 
0.0 0.3113 0 -2.0 1e-06 
0.0 0.3114 0 -2.0 1e-06 
0.0 0.3115 0 -2.0 1e-06 
0.0 0.3116 0 -2.0 1e-06 
0.0 0.3117 0 -2.0 1e-06 
0.0 0.3118 0 -2.0 1e-06 
0.0 0.3119 0 -2.0 1e-06 
0.0 0.312 0 -2.0 1e-06 
0.0 0.3121 0 -2.0 1e-06 
0.0 0.3122 0 -2.0 1e-06 
0.0 0.3123 0 -2.0 1e-06 
0.0 0.3124 0 -2.0 1e-06 
0.0 0.3125 0 -2.0 1e-06 
0.0 0.3126 0 -2.0 1e-06 
0.0 0.3127 0 -2.0 1e-06 
0.0 0.3128 0 -2.0 1e-06 
0.0 0.3129 0 -2.0 1e-06 
0.0 0.313 0 -2.0 1e-06 
0.0 0.3131 0 -2.0 1e-06 
0.0 0.3132 0 -2.0 1e-06 
0.0 0.3133 0 -2.0 1e-06 
0.0 0.3134 0 -2.0 1e-06 
0.0 0.3135 0 -2.0 1e-06 
0.0 0.3136 0 -2.0 1e-06 
0.0 0.3137 0 -2.0 1e-06 
0.0 0.3138 0 -2.0 1e-06 
0.0 0.3139 0 -2.0 1e-06 
0.0 0.314 0 -2.0 1e-06 
0.0 0.3141 0 -2.0 1e-06 
0.0 0.3142 0 -2.0 1e-06 
0.0 0.3143 0 -2.0 1e-06 
0.0 0.3144 0 -2.0 1e-06 
0.0 0.3145 0 -2.0 1e-06 
0.0 0.3146 0 -2.0 1e-06 
0.0 0.3147 0 -2.0 1e-06 
0.0 0.3148 0 -2.0 1e-06 
0.0 0.3149 0 -2.0 1e-06 
0.0 0.315 0 -2.0 1e-06 
0.0 0.3151 0 -2.0 1e-06 
0.0 0.3152 0 -2.0 1e-06 
0.0 0.3153 0 -2.0 1e-06 
0.0 0.3154 0 -2.0 1e-06 
0.0 0.3155 0 -2.0 1e-06 
0.0 0.3156 0 -2.0 1e-06 
0.0 0.3157 0 -2.0 1e-06 
0.0 0.3158 0 -2.0 1e-06 
0.0 0.3159 0 -2.0 1e-06 
0.0 0.316 0 -2.0 1e-06 
0.0 0.3161 0 -2.0 1e-06 
0.0 0.3162 0 -2.0 1e-06 
0.0 0.3163 0 -2.0 1e-06 
0.0 0.3164 0 -2.0 1e-06 
0.0 0.3165 0 -2.0 1e-06 
0.0 0.3166 0 -2.0 1e-06 
0.0 0.3167 0 -2.0 1e-06 
0.0 0.3168 0 -2.0 1e-06 
0.0 0.3169 0 -2.0 1e-06 
0.0 0.317 0 -2.0 1e-06 
0.0 0.3171 0 -2.0 1e-06 
0.0 0.3172 0 -2.0 1e-06 
0.0 0.3173 0 -2.0 1e-06 
0.0 0.3174 0 -2.0 1e-06 
0.0 0.3175 0 -2.0 1e-06 
0.0 0.3176 0 -2.0 1e-06 
0.0 0.3177 0 -2.0 1e-06 
0.0 0.3178 0 -2.0 1e-06 
0.0 0.3179 0 -2.0 1e-06 
0.0 0.318 0 -2.0 1e-06 
0.0 0.3181 0 -2.0 1e-06 
0.0 0.3182 0 -2.0 1e-06 
0.0 0.3183 0 -2.0 1e-06 
0.0 0.3184 0 -2.0 1e-06 
0.0 0.3185 0 -2.0 1e-06 
0.0 0.3186 0 -2.0 1e-06 
0.0 0.3187 0 -2.0 1e-06 
0.0 0.3188 0 -2.0 1e-06 
0.0 0.3189 0 -2.0 1e-06 
0.0 0.319 0 -2.0 1e-06 
0.0 0.3191 0 -2.0 1e-06 
0.0 0.3192 0 -2.0 1e-06 
0.0 0.3193 0 -2.0 1e-06 
0.0 0.3194 0 -2.0 1e-06 
0.0 0.3195 0 -2.0 1e-06 
0.0 0.3196 0 -2.0 1e-06 
0.0 0.3197 0 -2.0 1e-06 
0.0 0.3198 0 -2.0 1e-06 
0.0 0.3199 0 -2.0 1e-06 
0.0 0.32 0 -2.0 1e-06 
0.0 0.3201 0 -2.0 1e-06 
0.0 0.3202 0 -2.0 1e-06 
0.0 0.3203 0 -2.0 1e-06 
0.0 0.3204 0 -2.0 1e-06 
0.0 0.3205 0 -2.0 1e-06 
0.0 0.3206 0 -2.0 1e-06 
0.0 0.3207 0 -2.0 1e-06 
0.0 0.3208 0 -2.0 1e-06 
0.0 0.3209 0 -2.0 1e-06 
0.0 0.321 0 -2.0 1e-06 
0.0 0.3211 0 -2.0 1e-06 
0.0 0.3212 0 -2.0 1e-06 
0.0 0.3213 0 -2.0 1e-06 
0.0 0.3214 0 -2.0 1e-06 
0.0 0.3215 0 -2.0 1e-06 
0.0 0.3216 0 -2.0 1e-06 
0.0 0.3217 0 -2.0 1e-06 
0.0 0.3218 0 -2.0 1e-06 
0.0 0.3219 0 -2.0 1e-06 
0.0 0.322 0 -2.0 1e-06 
0.0 0.3221 0 -2.0 1e-06 
0.0 0.3222 0 -2.0 1e-06 
0.0 0.3223 0 -2.0 1e-06 
0.0 0.3224 0 -2.0 1e-06 
0.0 0.3225 0 -2.0 1e-06 
0.0 0.3226 0 -2.0 1e-06 
0.0 0.3227 0 -2.0 1e-06 
0.0 0.3228 0 -2.0 1e-06 
0.0 0.3229 0 -2.0 1e-06 
0.0 0.323 0 -2.0 1e-06 
0.0 0.3231 0 -2.0 1e-06 
0.0 0.3232 0 -2.0 1e-06 
0.0 0.3233 0 -2.0 1e-06 
0.0 0.3234 0 -2.0 1e-06 
0.0 0.3235 0 -2.0 1e-06 
0.0 0.3236 0 -2.0 1e-06 
0.0 0.3237 0 -2.0 1e-06 
0.0 0.3238 0 -2.0 1e-06 
0.0 0.3239 0 -2.0 1e-06 
0.0 0.324 0 -2.0 1e-06 
0.0 0.3241 0 -2.0 1e-06 
0.0 0.3242 0 -2.0 1e-06 
0.0 0.3243 0 -2.0 1e-06 
0.0 0.3244 0 -2.0 1e-06 
0.0 0.3245 0 -2.0 1e-06 
0.0 0.3246 0 -2.0 1e-06 
0.0 0.3247 0 -2.0 1e-06 
0.0 0.3248 0 -2.0 1e-06 
0.0 0.3249 0 -2.0 1e-06 
0.0 0.325 0 -2.0 1e-06 
0.0 0.3251 0 -2.0 1e-06 
0.0 0.3252 0 -2.0 1e-06 
0.0 0.3253 0 -2.0 1e-06 
0.0 0.3254 0 -2.0 1e-06 
0.0 0.3255 0 -2.0 1e-06 
0.0 0.3256 0 -2.0 1e-06 
0.0 0.3257 0 -2.0 1e-06 
0.0 0.3258 0 -2.0 1e-06 
0.0 0.3259 0 -2.0 1e-06 
0.0 0.326 0 -2.0 1e-06 
0.0 0.3261 0 -2.0 1e-06 
0.0 0.3262 0 -2.0 1e-06 
0.0 0.3263 0 -2.0 1e-06 
0.0 0.3264 0 -2.0 1e-06 
0.0 0.3265 0 -2.0 1e-06 
0.0 0.3266 0 -2.0 1e-06 
0.0 0.3267 0 -2.0 1e-06 
0.0 0.3268 0 -2.0 1e-06 
0.0 0.3269 0 -2.0 1e-06 
0.0 0.327 0 -2.0 1e-06 
0.0 0.3271 0 -2.0 1e-06 
0.0 0.3272 0 -2.0 1e-06 
0.0 0.3273 0 -2.0 1e-06 
0.0 0.3274 0 -2.0 1e-06 
0.0 0.3275 0 -2.0 1e-06 
0.0 0.3276 0 -2.0 1e-06 
0.0 0.3277 0 -2.0 1e-06 
0.0 0.3278 0 -2.0 1e-06 
0.0 0.3279 0 -2.0 1e-06 
0.0 0.328 0 -2.0 1e-06 
0.0 0.3281 0 -2.0 1e-06 
0.0 0.3282 0 -2.0 1e-06 
0.0 0.3283 0 -2.0 1e-06 
0.0 0.3284 0 -2.0 1e-06 
0.0 0.3285 0 -2.0 1e-06 
0.0 0.3286 0 -2.0 1e-06 
0.0 0.3287 0 -2.0 1e-06 
0.0 0.3288 0 -2.0 1e-06 
0.0 0.3289 0 -2.0 1e-06 
0.0 0.329 0 -2.0 1e-06 
0.0 0.3291 0 -2.0 1e-06 
0.0 0.3292 0 -2.0 1e-06 
0.0 0.3293 0 -2.0 1e-06 
0.0 0.3294 0 -2.0 1e-06 
0.0 0.3295 0 -2.0 1e-06 
0.0 0.3296 0 -2.0 1e-06 
0.0 0.3297 0 -2.0 1e-06 
0.0 0.3298 0 -2.0 1e-06 
0.0 0.3299 0 -2.0 1e-06 
0.0 0.33 0 -2.0 1e-06 
0.0 0.3301 0 -2.0 1e-06 
0.0 0.3302 0 -2.0 1e-06 
0.0 0.3303 0 -2.0 1e-06 
0.0 0.3304 0 -2.0 1e-06 
0.0 0.3305 0 -2.0 1e-06 
0.0 0.3306 0 -2.0 1e-06 
0.0 0.3307 0 -2.0 1e-06 
0.0 0.3308 0 -2.0 1e-06 
0.0 0.3309 0 -2.0 1e-06 
0.0 0.331 0 -2.0 1e-06 
0.0 0.3311 0 -2.0 1e-06 
0.0 0.3312 0 -2.0 1e-06 
0.0 0.3313 0 -2.0 1e-06 
0.0 0.3314 0 -2.0 1e-06 
0.0 0.3315 0 -2.0 1e-06 
0.0 0.3316 0 -2.0 1e-06 
0.0 0.3317 0 -2.0 1e-06 
0.0 0.3318 0 -2.0 1e-06 
0.0 0.3319 0 -2.0 1e-06 
0.0 0.332 0 -2.0 1e-06 
0.0 0.3321 0 -2.0 1e-06 
0.0 0.3322 0 -2.0 1e-06 
0.0 0.3323 0 -2.0 1e-06 
0.0 0.3324 0 -2.0 1e-06 
0.0 0.3325 0 -2.0 1e-06 
0.0 0.3326 0 -2.0 1e-06 
0.0 0.3327 0 -2.0 1e-06 
0.0 0.3328 0 -2.0 1e-06 
0.0 0.3329 0 -2.0 1e-06 
0.0 0.333 0 -2.0 1e-06 
0.0 0.3331 0 -2.0 1e-06 
0.0 0.3332 0 -2.0 1e-06 
0.0 0.3333 0 -2.0 1e-06 
0.0 0.3334 0 -2.0 1e-06 
0.0 0.3335 0 -2.0 1e-06 
0.0 0.3336 0 -2.0 1e-06 
0.0 0.3337 0 -2.0 1e-06 
0.0 0.3338 0 -2.0 1e-06 
0.0 0.3339 0 -2.0 1e-06 
0.0 0.334 0 -2.0 1e-06 
0.0 0.3341 0 -2.0 1e-06 
0.0 0.3342 0 -2.0 1e-06 
0.0 0.3343 0 -2.0 1e-06 
0.0 0.3344 0 -2.0 1e-06 
0.0 0.3345 0 -2.0 1e-06 
0.0 0.3346 0 -2.0 1e-06 
0.0 0.3347 0 -2.0 1e-06 
0.0 0.3348 0 -2.0 1e-06 
0.0 0.3349 0 -2.0 1e-06 
0.0 0.335 0 -2.0 1e-06 
0.0 0.3351 0 -2.0 1e-06 
0.0 0.3352 0 -2.0 1e-06 
0.0 0.3353 0 -2.0 1e-06 
0.0 0.3354 0 -2.0 1e-06 
0.0 0.3355 0 -2.0 1e-06 
0.0 0.3356 0 -2.0 1e-06 
0.0 0.3357 0 -2.0 1e-06 
0.0 0.3358 0 -2.0 1e-06 
0.0 0.3359 0 -2.0 1e-06 
0.0 0.336 0 -2.0 1e-06 
0.0 0.3361 0 -2.0 1e-06 
0.0 0.3362 0 -2.0 1e-06 
0.0 0.3363 0 -2.0 1e-06 
0.0 0.3364 0 -2.0 1e-06 
0.0 0.3365 0 -2.0 1e-06 
0.0 0.3366 0 -2.0 1e-06 
0.0 0.3367 0 -2.0 1e-06 
0.0 0.3368 0 -2.0 1e-06 
0.0 0.3369 0 -2.0 1e-06 
0.0 0.337 0 -2.0 1e-06 
0.0 0.3371 0 -2.0 1e-06 
0.0 0.3372 0 -2.0 1e-06 
0.0 0.3373 0 -2.0 1e-06 
0.0 0.3374 0 -2.0 1e-06 
0.0 0.3375 0 -2.0 1e-06 
0.0 0.3376 0 -2.0 1e-06 
0.0 0.3377 0 -2.0 1e-06 
0.0 0.3378 0 -2.0 1e-06 
0.0 0.3379 0 -2.0 1e-06 
0.0 0.338 0 -2.0 1e-06 
0.0 0.3381 0 -2.0 1e-06 
0.0 0.3382 0 -2.0 1e-06 
0.0 0.3383 0 -2.0 1e-06 
0.0 0.3384 0 -2.0 1e-06 
0.0 0.3385 0 -2.0 1e-06 
0.0 0.3386 0 -2.0 1e-06 
0.0 0.3387 0 -2.0 1e-06 
0.0 0.3388 0 -2.0 1e-06 
0.0 0.3389 0 -2.0 1e-06 
0.0 0.339 0 -2.0 1e-06 
0.0 0.3391 0 -2.0 1e-06 
0.0 0.3392 0 -2.0 1e-06 
0.0 0.3393 0 -2.0 1e-06 
0.0 0.3394 0 -2.0 1e-06 
0.0 0.3395 0 -2.0 1e-06 
0.0 0.3396 0 -2.0 1e-06 
0.0 0.3397 0 -2.0 1e-06 
0.0 0.3398 0 -2.0 1e-06 
0.0 0.3399 0 -2.0 1e-06 
0.0 0.34 0 -2.0 1e-06 
0.0 0.3401 0 -2.0 1e-06 
0.0 0.3402 0 -2.0 1e-06 
0.0 0.3403 0 -2.0 1e-06 
0.0 0.3404 0 -2.0 1e-06 
0.0 0.3405 0 -2.0 1e-06 
0.0 0.3406 0 -2.0 1e-06 
0.0 0.3407 0 -2.0 1e-06 
0.0 0.3408 0 -2.0 1e-06 
0.0 0.3409 0 -2.0 1e-06 
0.0 0.341 0 -2.0 1e-06 
0.0 0.3411 0 -2.0 1e-06 
0.0 0.3412 0 -2.0 1e-06 
0.0 0.3413 0 -2.0 1e-06 
0.0 0.3414 0 -2.0 1e-06 
0.0 0.3415 0 -2.0 1e-06 
0.0 0.3416 0 -2.0 1e-06 
0.0 0.3417 0 -2.0 1e-06 
0.0 0.3418 0 -2.0 1e-06 
0.0 0.3419 0 -2.0 1e-06 
0.0 0.342 0 -2.0 1e-06 
0.0 0.3421 0 -2.0 1e-06 
0.0 0.3422 0 -2.0 1e-06 
0.0 0.3423 0 -2.0 1e-06 
0.0 0.3424 0 -2.0 1e-06 
0.0 0.3425 0 -2.0 1e-06 
0.0 0.3426 0 -2.0 1e-06 
0.0 0.3427 0 -2.0 1e-06 
0.0 0.3428 0 -2.0 1e-06 
0.0 0.3429 0 -2.0 1e-06 
0.0 0.343 0 -2.0 1e-06 
0.0 0.3431 0 -2.0 1e-06 
0.0 0.3432 0 -2.0 1e-06 
0.0 0.3433 0 -2.0 1e-06 
0.0 0.3434 0 -2.0 1e-06 
0.0 0.3435 0 -2.0 1e-06 
0.0 0.3436 0 -2.0 1e-06 
0.0 0.3437 0 -2.0 1e-06 
0.0 0.3438 0 -2.0 1e-06 
0.0 0.3439 0 -2.0 1e-06 
0.0 0.344 0 -2.0 1e-06 
0.0 0.3441 0 -2.0 1e-06 
0.0 0.3442 0 -2.0 1e-06 
0.0 0.3443 0 -2.0 1e-06 
0.0 0.3444 0 -2.0 1e-06 
0.0 0.3445 0 -2.0 1e-06 
0.0 0.3446 0 -2.0 1e-06 
0.0 0.3447 0 -2.0 1e-06 
0.0 0.3448 0 -2.0 1e-06 
0.0 0.3449 0 -2.0 1e-06 
0.0 0.345 0 -2.0 1e-06 
0.0 0.3451 0 -2.0 1e-06 
0.0 0.3452 0 -2.0 1e-06 
0.0 0.3453 0 -2.0 1e-06 
0.0 0.3454 0 -2.0 1e-06 
0.0 0.3455 0 -2.0 1e-06 
0.0 0.3456 0 -2.0 1e-06 
0.0 0.3457 0 -2.0 1e-06 
0.0 0.3458 0 -2.0 1e-06 
0.0 0.3459 0 -2.0 1e-06 
0.0 0.346 0 -2.0 1e-06 
0.0 0.3461 0 -2.0 1e-06 
0.0 0.3462 0 -2.0 1e-06 
0.0 0.3463 0 -2.0 1e-06 
0.0 0.3464 0 -2.0 1e-06 
0.0 0.3465 0 -2.0 1e-06 
0.0 0.3466 0 -2.0 1e-06 
0.0 0.3467 0 -2.0 1e-06 
0.0 0.3468 0 -2.0 1e-06 
0.0 0.3469 0 -2.0 1e-06 
0.0 0.347 0 -2.0 1e-06 
0.0 0.3471 0 -2.0 1e-06 
0.0 0.3472 0 -2.0 1e-06 
0.0 0.3473 0 -2.0 1e-06 
0.0 0.3474 0 -2.0 1e-06 
0.0 0.3475 0 -2.0 1e-06 
0.0 0.3476 0 -2.0 1e-06 
0.0 0.3477 0 -2.0 1e-06 
0.0 0.3478 0 -2.0 1e-06 
0.0 0.3479 0 -2.0 1e-06 
0.0 0.348 0 -2.0 1e-06 
0.0 0.3481 0 -2.0 1e-06 
0.0 0.3482 0 -2.0 1e-06 
0.0 0.3483 0 -2.0 1e-06 
0.0 0.3484 0 -2.0 1e-06 
0.0 0.3485 0 -2.0 1e-06 
0.0 0.3486 0 -2.0 1e-06 
0.0 0.3487 0 -2.0 1e-06 
0.0 0.3488 0 -2.0 1e-06 
0.0 0.3489 0 -2.0 1e-06 
0.0 0.349 0 -2.0 1e-06 
0.0 0.3491 0 -2.0 1e-06 
0.0 0.3492 0 -2.0 1e-06 
0.0 0.3493 0 -2.0 1e-06 
0.0 0.3494 0 -2.0 1e-06 
0.0 0.3495 0 -2.0 1e-06 
0.0 0.3496 0 -2.0 1e-06 
0.0 0.3497 0 -2.0 1e-06 
0.0 0.3498 0 -2.0 1e-06 
0.0 0.3499 0 -2.0 1e-06 
0.0 0.35 0 -2.0 1e-06 
0.0 0.3501 0 -2.0 1e-06 
0.0 0.3502 0 -2.0 1e-06 
0.0 0.3503 0 -2.0 1e-06 
0.0 0.3504 0 -2.0 1e-06 
0.0 0.3505 0 -2.0 1e-06 
0.0 0.3506 0 -2.0 1e-06 
0.0 0.3507 0 -2.0 1e-06 
0.0 0.3508 0 -2.0 1e-06 
0.0 0.3509 0 -2.0 1e-06 
0.0 0.351 0 -2.0 1e-06 
0.0 0.3511 0 -2.0 1e-06 
0.0 0.3512 0 -2.0 1e-06 
0.0 0.3513 0 -2.0 1e-06 
0.0 0.3514 0 -2.0 1e-06 
0.0 0.3515 0 -2.0 1e-06 
0.0 0.3516 0 -2.0 1e-06 
0.0 0.3517 0 -2.0 1e-06 
0.0 0.3518 0 -2.0 1e-06 
0.0 0.3519 0 -2.0 1e-06 
0.0 0.352 0 -2.0 1e-06 
0.0 0.3521 0 -2.0 1e-06 
0.0 0.3522 0 -2.0 1e-06 
0.0 0.3523 0 -2.0 1e-06 
0.0 0.3524 0 -2.0 1e-06 
0.0 0.3525 0 -2.0 1e-06 
0.0 0.3526 0 -2.0 1e-06 
0.0 0.3527 0 -2.0 1e-06 
0.0 0.3528 0 -2.0 1e-06 
0.0 0.3529 0 -2.0 1e-06 
0.0 0.353 0 -2.0 1e-06 
0.0 0.3531 0 -2.0 1e-06 
0.0 0.3532 0 -2.0 1e-06 
0.0 0.3533 0 -2.0 1e-06 
0.0 0.3534 0 -2.0 1e-06 
0.0 0.3535 0 -2.0 1e-06 
0.0 0.3536 0 -2.0 1e-06 
0.0 0.3537 0 -2.0 1e-06 
0.0 0.3538 0 -2.0 1e-06 
0.0 0.3539 0 -2.0 1e-06 
0.0 0.354 0 -2.0 1e-06 
0.0 0.3541 0 -2.0 1e-06 
0.0 0.3542 0 -2.0 1e-06 
0.0 0.3543 0 -2.0 1e-06 
0.0 0.3544 0 -2.0 1e-06 
0.0 0.3545 0 -2.0 1e-06 
0.0 0.3546 0 -2.0 1e-06 
0.0 0.3547 0 -2.0 1e-06 
0.0 0.3548 0 -2.0 1e-06 
0.0 0.3549 0 -2.0 1e-06 
0.0 0.355 0 -2.0 1e-06 
0.0 0.3551 0 -2.0 1e-06 
0.0 0.3552 0 -2.0 1e-06 
0.0 0.3553 0 -2.0 1e-06 
0.0 0.3554 0 -2.0 1e-06 
0.0 0.3555 0 -2.0 1e-06 
0.0 0.3556 0 -2.0 1e-06 
0.0 0.3557 0 -2.0 1e-06 
0.0 0.3558 0 -2.0 1e-06 
0.0 0.3559 0 -2.0 1e-06 
0.0 0.356 0 -2.0 1e-06 
0.0 0.3561 0 -2.0 1e-06 
0.0 0.3562 0 -2.0 1e-06 
0.0 0.3563 0 -2.0 1e-06 
0.0 0.3564 0 -2.0 1e-06 
0.0 0.3565 0 -2.0 1e-06 
0.0 0.3566 0 -2.0 1e-06 
0.0 0.3567 0 -2.0 1e-06 
0.0 0.3568 0 -2.0 1e-06 
0.0 0.3569 0 -2.0 1e-06 
0.0 0.357 0 -2.0 1e-06 
0.0 0.3571 0 -2.0 1e-06 
0.0 0.3572 0 -2.0 1e-06 
0.0 0.3573 0 -2.0 1e-06 
0.0 0.3574 0 -2.0 1e-06 
0.0 0.3575 0 -2.0 1e-06 
0.0 0.3576 0 -2.0 1e-06 
0.0 0.3577 0 -2.0 1e-06 
0.0 0.3578 0 -2.0 1e-06 
0.0 0.3579 0 -2.0 1e-06 
0.0 0.358 0 -2.0 1e-06 
0.0 0.3581 0 -2.0 1e-06 
0.0 0.3582 0 -2.0 1e-06 
0.0 0.3583 0 -2.0 1e-06 
0.0 0.3584 0 -2.0 1e-06 
0.0 0.3585 0 -2.0 1e-06 
0.0 0.3586 0 -2.0 1e-06 
0.0 0.3587 0 -2.0 1e-06 
0.0 0.3588 0 -2.0 1e-06 
0.0 0.3589 0 -2.0 1e-06 
0.0 0.359 0 -2.0 1e-06 
0.0 0.3591 0 -2.0 1e-06 
0.0 0.3592 0 -2.0 1e-06 
0.0 0.3593 0 -2.0 1e-06 
0.0 0.3594 0 -2.0 1e-06 
0.0 0.3595 0 -2.0 1e-06 
0.0 0.3596 0 -2.0 1e-06 
0.0 0.3597 0 -2.0 1e-06 
0.0 0.3598 0 -2.0 1e-06 
0.0 0.3599 0 -2.0 1e-06 
0.0 0.36 0 -2.0 1e-06 
0.0 0.3601 0 -2.0 1e-06 
0.0 0.3602 0 -2.0 1e-06 
0.0 0.3603 0 -2.0 1e-06 
0.0 0.3604 0 -2.0 1e-06 
0.0 0.3605 0 -2.0 1e-06 
0.0 0.3606 0 -2.0 1e-06 
0.0 0.3607 0 -2.0 1e-06 
0.0 0.3608 0 -2.0 1e-06 
0.0 0.3609 0 -2.0 1e-06 
0.0 0.361 0 -2.0 1e-06 
0.0 0.3611 0 -2.0 1e-06 
0.0 0.3612 0 -2.0 1e-06 
0.0 0.3613 0 -2.0 1e-06 
0.0 0.3614 0 -2.0 1e-06 
0.0 0.3615 0 -2.0 1e-06 
0.0 0.3616 0 -2.0 1e-06 
0.0 0.3617 0 -2.0 1e-06 
0.0 0.3618 0 -2.0 1e-06 
0.0 0.3619 0 -2.0 1e-06 
0.0 0.362 0 -2.0 1e-06 
0.0 0.3621 0 -2.0 1e-06 
0.0 0.3622 0 -2.0 1e-06 
0.0 0.3623 0 -2.0 1e-06 
0.0 0.3624 0 -2.0 1e-06 
0.0 0.3625 0 -2.0 1e-06 
0.0 0.3626 0 -2.0 1e-06 
0.0 0.3627 0 -2.0 1e-06 
0.0 0.3628 0 -2.0 1e-06 
0.0 0.3629 0 -2.0 1e-06 
0.0 0.363 0 -2.0 1e-06 
0.0 0.3631 0 -2.0 1e-06 
0.0 0.3632 0 -2.0 1e-06 
0.0 0.3633 0 -2.0 1e-06 
0.0 0.3634 0 -2.0 1e-06 
0.0 0.3635 0 -2.0 1e-06 
0.0 0.3636 0 -2.0 1e-06 
0.0 0.3637 0 -2.0 1e-06 
0.0 0.3638 0 -2.0 1e-06 
0.0 0.3639 0 -2.0 1e-06 
0.0 0.364 0 -2.0 1e-06 
0.0 0.3641 0 -2.0 1e-06 
0.0 0.3642 0 -2.0 1e-06 
0.0 0.3643 0 -2.0 1e-06 
0.0 0.3644 0 -2.0 1e-06 
0.0 0.3645 0 -2.0 1e-06 
0.0 0.3646 0 -2.0 1e-06 
0.0 0.3647 0 -2.0 1e-06 
0.0 0.3648 0 -2.0 1e-06 
0.0 0.3649 0 -2.0 1e-06 
0.0 0.365 0 -2.0 1e-06 
0.0 0.3651 0 -2.0 1e-06 
0.0 0.3652 0 -2.0 1e-06 
0.0 0.3653 0 -2.0 1e-06 
0.0 0.3654 0 -2.0 1e-06 
0.0 0.3655 0 -2.0 1e-06 
0.0 0.3656 0 -2.0 1e-06 
0.0 0.3657 0 -2.0 1e-06 
0.0 0.3658 0 -2.0 1e-06 
0.0 0.3659 0 -2.0 1e-06 
0.0 0.366 0 -2.0 1e-06 
0.0 0.3661 0 -2.0 1e-06 
0.0 0.3662 0 -2.0 1e-06 
0.0 0.3663 0 -2.0 1e-06 
0.0 0.3664 0 -2.0 1e-06 
0.0 0.3665 0 -2.0 1e-06 
0.0 0.3666 0 -2.0 1e-06 
0.0 0.3667 0 -2.0 1e-06 
0.0 0.3668 0 -2.0 1e-06 
0.0 0.3669 0 -2.0 1e-06 
0.0 0.367 0 -2.0 1e-06 
0.0 0.3671 0 -2.0 1e-06 
0.0 0.3672 0 -2.0 1e-06 
0.0 0.3673 0 -2.0 1e-06 
0.0 0.3674 0 -2.0 1e-06 
0.0 0.3675 0 -2.0 1e-06 
0.0 0.3676 0 -2.0 1e-06 
0.0 0.3677 0 -2.0 1e-06 
0.0 0.3678 0 -2.0 1e-06 
0.0 0.3679 0 -2.0 1e-06 
0.0 0.368 0 -2.0 1e-06 
0.0 0.3681 0 -2.0 1e-06 
0.0 0.3682 0 -2.0 1e-06 
0.0 0.3683 0 -2.0 1e-06 
0.0 0.3684 0 -2.0 1e-06 
0.0 0.3685 0 -2.0 1e-06 
0.0 0.3686 0 -2.0 1e-06 
0.0 0.3687 0 -2.0 1e-06 
0.0 0.3688 0 -2.0 1e-06 
0.0 0.3689 0 -2.0 1e-06 
0.0 0.369 0 -2.0 1e-06 
0.0 0.3691 0 -2.0 1e-06 
0.0 0.3692 0 -2.0 1e-06 
0.0 0.3693 0 -2.0 1e-06 
0.0 0.3694 0 -2.0 1e-06 
0.0 0.3695 0 -2.0 1e-06 
0.0 0.3696 0 -2.0 1e-06 
0.0 0.3697 0 -2.0 1e-06 
0.0 0.3698 0 -2.0 1e-06 
0.0 0.3699 0 -2.0 1e-06 
0.0 0.37 0 -2.0 1e-06 
0.0 0.3701 0 -2.0 1e-06 
0.0 0.3702 0 -2.0 1e-06 
0.0 0.3703 0 -2.0 1e-06 
0.0 0.3704 0 -2.0 1e-06 
0.0 0.3705 0 -2.0 1e-06 
0.0 0.3706 0 -2.0 1e-06 
0.0 0.3707 0 -2.0 1e-06 
0.0 0.3708 0 -2.0 1e-06 
0.0 0.3709 0 -2.0 1e-06 
0.0 0.371 0 -2.0 1e-06 
0.0 0.3711 0 -2.0 1e-06 
0.0 0.3712 0 -2.0 1e-06 
0.0 0.3713 0 -2.0 1e-06 
0.0 0.3714 0 -2.0 1e-06 
0.0 0.3715 0 -2.0 1e-06 
0.0 0.3716 0 -2.0 1e-06 
0.0 0.3717 0 -2.0 1e-06 
0.0 0.3718 0 -2.0 1e-06 
0.0 0.3719 0 -2.0 1e-06 
0.0 0.372 0 -2.0 1e-06 
0.0 0.3721 0 -2.0 1e-06 
0.0 0.3722 0 -2.0 1e-06 
0.0 0.3723 0 -2.0 1e-06 
0.0 0.3724 0 -2.0 1e-06 
0.0 0.3725 0 -2.0 1e-06 
0.0 0.3726 0 -2.0 1e-06 
0.0 0.3727 0 -2.0 1e-06 
0.0 0.3728 0 -2.0 1e-06 
0.0 0.3729 0 -2.0 1e-06 
0.0 0.373 0 -2.0 1e-06 
0.0 0.3731 0 -2.0 1e-06 
0.0 0.3732 0 -2.0 1e-06 
0.0 0.3733 0 -2.0 1e-06 
0.0 0.3734 0 -2.0 1e-06 
0.0 0.3735 0 -2.0 1e-06 
0.0 0.3736 0 -2.0 1e-06 
0.0 0.3737 0 -2.0 1e-06 
0.0 0.3738 0 -2.0 1e-06 
0.0 0.3739 0 -2.0 1e-06 
0.0 0.374 0 -2.0 1e-06 
0.0 0.3741 0 -2.0 1e-06 
0.0 0.3742 0 -2.0 1e-06 
0.0 0.3743 0 -2.0 1e-06 
0.0 0.3744 0 -2.0 1e-06 
0.0 0.3745 0 -2.0 1e-06 
0.0 0.3746 0 -2.0 1e-06 
0.0 0.3747 0 -2.0 1e-06 
0.0 0.3748 0 -2.0 1e-06 
0.0 0.3749 0 -2.0 1e-06 
0.0 0.375 0 -2.0 1e-06 
0.0 0.3751 0 -2.0 1e-06 
0.0 0.3752 0 -2.0 1e-06 
0.0 0.3753 0 -2.0 1e-06 
0.0 0.3754 0 -2.0 1e-06 
0.0 0.3755 0 -2.0 1e-06 
0.0 0.3756 0 -2.0 1e-06 
0.0 0.3757 0 -2.0 1e-06 
0.0 0.3758 0 -2.0 1e-06 
0.0 0.3759 0 -2.0 1e-06 
0.0 0.376 0 -2.0 1e-06 
0.0 0.3761 0 -2.0 1e-06 
0.0 0.3762 0 -2.0 1e-06 
0.0 0.3763 0 -2.0 1e-06 
0.0 0.3764 0 -2.0 1e-06 
0.0 0.3765 0 -2.0 1e-06 
0.0 0.3766 0 -2.0 1e-06 
0.0 0.3767 0 -2.0 1e-06 
0.0 0.3768 0 -2.0 1e-06 
0.0 0.3769 0 -2.0 1e-06 
0.0 0.377 0 -2.0 1e-06 
0.0 0.3771 0 -2.0 1e-06 
0.0 0.3772 0 -2.0 1e-06 
0.0 0.3773 0 -2.0 1e-06 
0.0 0.3774 0 -2.0 1e-06 
0.0 0.3775 0 -2.0 1e-06 
0.0 0.3776 0 -2.0 1e-06 
0.0 0.3777 0 -2.0 1e-06 
0.0 0.3778 0 -2.0 1e-06 
0.0 0.3779 0 -2.0 1e-06 
0.0 0.378 0 -2.0 1e-06 
0.0 0.3781 0 -2.0 1e-06 
0.0 0.3782 0 -2.0 1e-06 
0.0 0.3783 0 -2.0 1e-06 
0.0 0.3784 0 -2.0 1e-06 
0.0 0.3785 0 -2.0 1e-06 
0.0 0.3786 0 -2.0 1e-06 
0.0 0.3787 0 -2.0 1e-06 
0.0 0.3788 0 -2.0 1e-06 
0.0 0.3789 0 -2.0 1e-06 
0.0 0.379 0 -2.0 1e-06 
0.0 0.3791 0 -2.0 1e-06 
0.0 0.3792 0 -2.0 1e-06 
0.0 0.3793 0 -2.0 1e-06 
0.0 0.3794 0 -2.0 1e-06 
0.0 0.3795 0 -2.0 1e-06 
0.0 0.3796 0 -2.0 1e-06 
0.0 0.3797 0 -2.0 1e-06 
0.0 0.3798 0 -2.0 1e-06 
0.0 0.3799 0 -2.0 1e-06 
0.0 0.38 0 -2.0 1e-06 
0.0 0.3801 0 -2.0 1e-06 
0.0 0.3802 0 -2.0 1e-06 
0.0 0.3803 0 -2.0 1e-06 
0.0 0.3804 0 -2.0 1e-06 
0.0 0.3805 0 -2.0 1e-06 
0.0 0.3806 0 -2.0 1e-06 
0.0 0.3807 0 -2.0 1e-06 
0.0 0.3808 0 -2.0 1e-06 
0.0 0.3809 0 -2.0 1e-06 
0.0 0.381 0 -2.0 1e-06 
0.0 0.3811 0 -2.0 1e-06 
0.0 0.3812 0 -2.0 1e-06 
0.0 0.3813 0 -2.0 1e-06 
0.0 0.3814 0 -2.0 1e-06 
0.0 0.3815 0 -2.0 1e-06 
0.0 0.3816 0 -2.0 1e-06 
0.0 0.3817 0 -2.0 1e-06 
0.0 0.3818 0 -2.0 1e-06 
0.0 0.3819 0 -2.0 1e-06 
0.0 0.382 0 -2.0 1e-06 
0.0 0.3821 0 -2.0 1e-06 
0.0 0.3822 0 -2.0 1e-06 
0.0 0.3823 0 -2.0 1e-06 
0.0 0.3824 0 -2.0 1e-06 
0.0 0.3825 0 -2.0 1e-06 
0.0 0.3826 0 -2.0 1e-06 
0.0 0.3827 0 -2.0 1e-06 
0.0 0.3828 0 -2.0 1e-06 
0.0 0.3829 0 -2.0 1e-06 
0.0 0.383 0 -2.0 1e-06 
0.0 0.3831 0 -2.0 1e-06 
0.0 0.3832 0 -2.0 1e-06 
0.0 0.3833 0 -2.0 1e-06 
0.0 0.3834 0 -2.0 1e-06 
0.0 0.3835 0 -2.0 1e-06 
0.0 0.3836 0 -2.0 1e-06 
0.0 0.3837 0 -2.0 1e-06 
0.0 0.3838 0 -2.0 1e-06 
0.0 0.3839 0 -2.0 1e-06 
0.0 0.384 0 -2.0 1e-06 
0.0 0.3841 0 -2.0 1e-06 
0.0 0.3842 0 -2.0 1e-06 
0.0 0.3843 0 -2.0 1e-06 
0.0 0.3844 0 -2.0 1e-06 
0.0 0.3845 0 -2.0 1e-06 
0.0 0.3846 0 -2.0 1e-06 
0.0 0.3847 0 -2.0 1e-06 
0.0 0.3848 0 -2.0 1e-06 
0.0 0.3849 0 -2.0 1e-06 
0.0 0.385 0 -2.0 1e-06 
0.0 0.3851 0 -2.0 1e-06 
0.0 0.3852 0 -2.0 1e-06 
0.0 0.3853 0 -2.0 1e-06 
0.0 0.3854 0 -2.0 1e-06 
0.0 0.3855 0 -2.0 1e-06 
0.0 0.3856 0 -2.0 1e-06 
0.0 0.3857 0 -2.0 1e-06 
0.0 0.3858 0 -2.0 1e-06 
0.0 0.3859 0 -2.0 1e-06 
0.0 0.386 0 -2.0 1e-06 
0.0 0.3861 0 -2.0 1e-06 
0.0 0.3862 0 -2.0 1e-06 
0.0 0.3863 0 -2.0 1e-06 
0.0 0.3864 0 -2.0 1e-06 
0.0 0.3865 0 -2.0 1e-06 
0.0 0.3866 0 -2.0 1e-06 
0.0 0.3867 0 -2.0 1e-06 
0.0 0.3868 0 -2.0 1e-06 
0.0 0.3869 0 -2.0 1e-06 
0.0 0.387 0 -2.0 1e-06 
0.0 0.3871 0 -2.0 1e-06 
0.0 0.3872 0 -2.0 1e-06 
0.0 0.3873 0 -2.0 1e-06 
0.0 0.3874 0 -2.0 1e-06 
0.0 0.3875 0 -2.0 1e-06 
0.0 0.3876 0 -2.0 1e-06 
0.0 0.3877 0 -2.0 1e-06 
0.0 0.3878 0 -2.0 1e-06 
0.0 0.3879 0 -2.0 1e-06 
0.0 0.388 0 -2.0 1e-06 
0.0 0.3881 0 -2.0 1e-06 
0.0 0.3882 0 -2.0 1e-06 
0.0 0.3883 0 -2.0 1e-06 
0.0 0.3884 0 -2.0 1e-06 
0.0 0.3885 0 -2.0 1e-06 
0.0 0.3886 0 -2.0 1e-06 
0.0 0.3887 0 -2.0 1e-06 
0.0 0.3888 0 -2.0 1e-06 
0.0 0.3889 0 -2.0 1e-06 
0.0 0.389 0 -2.0 1e-06 
0.0 0.3891 0 -2.0 1e-06 
0.0 0.3892 0 -2.0 1e-06 
0.0 0.3893 0 -2.0 1e-06 
0.0 0.3894 0 -2.0 1e-06 
0.0 0.3895 0 -2.0 1e-06 
0.0 0.3896 0 -2.0 1e-06 
0.0 0.3897 0 -2.0 1e-06 
0.0 0.3898 0 -2.0 1e-06 
0.0 0.3899 0 -2.0 1e-06 
0.0 0.39 0 -2.0 1e-06 
0.0 0.3901 0 -2.0 1e-06 
0.0 0.3902 0 -2.0 1e-06 
0.0 0.3903 0 -2.0 1e-06 
0.0 0.3904 0 -2.0 1e-06 
0.0 0.3905 0 -2.0 1e-06 
0.0 0.3906 0 -2.0 1e-06 
0.0 0.3907 0 -2.0 1e-06 
0.0 0.3908 0 -2.0 1e-06 
0.0 0.3909 0 -2.0 1e-06 
0.0 0.391 0 -2.0 1e-06 
0.0 0.3911 0 -2.0 1e-06 
0.0 0.3912 0 -2.0 1e-06 
0.0 0.3913 0 -2.0 1e-06 
0.0 0.3914 0 -2.0 1e-06 
0.0 0.3915 0 -2.0 1e-06 
0.0 0.3916 0 -2.0 1e-06 
0.0 0.3917 0 -2.0 1e-06 
0.0 0.3918 0 -2.0 1e-06 
0.0 0.3919 0 -2.0 1e-06 
0.0 0.392 0 -2.0 1e-06 
0.0 0.3921 0 -2.0 1e-06 
0.0 0.3922 0 -2.0 1e-06 
0.0 0.3923 0 -2.0 1e-06 
0.0 0.3924 0 -2.0 1e-06 
0.0 0.3925 0 -2.0 1e-06 
0.0 0.3926 0 -2.0 1e-06 
0.0 0.3927 0 -2.0 1e-06 
0.0 0.3928 0 -2.0 1e-06 
0.0 0.3929 0 -2.0 1e-06 
0.0 0.393 0 -2.0 1e-06 
0.0 0.3931 0 -2.0 1e-06 
0.0 0.3932 0 -2.0 1e-06 
0.0 0.3933 0 -2.0 1e-06 
0.0 0.3934 0 -2.0 1e-06 
0.0 0.3935 0 -2.0 1e-06 
0.0 0.3936 0 -2.0 1e-06 
0.0 0.3937 0 -2.0 1e-06 
0.0 0.3938 0 -2.0 1e-06 
0.0 0.3939 0 -2.0 1e-06 
0.0 0.394 0 -2.0 1e-06 
0.0 0.3941 0 -2.0 1e-06 
0.0 0.3942 0 -2.0 1e-06 
0.0 0.3943 0 -2.0 1e-06 
0.0 0.3944 0 -2.0 1e-06 
0.0 0.3945 0 -2.0 1e-06 
0.0 0.3946 0 -2.0 1e-06 
0.0 0.3947 0 -2.0 1e-06 
0.0 0.3948 0 -2.0 1e-06 
0.0 0.3949 0 -2.0 1e-06 
0.0 0.395 0 -2.0 1e-06 
0.0 0.3951 0 -2.0 1e-06 
0.0 0.3952 0 -2.0 1e-06 
0.0 0.3953 0 -2.0 1e-06 
0.0 0.3954 0 -2.0 1e-06 
0.0 0.3955 0 -2.0 1e-06 
0.0 0.3956 0 -2.0 1e-06 
0.0 0.3957 0 -2.0 1e-06 
0.0 0.3958 0 -2.0 1e-06 
0.0 0.3959 0 -2.0 1e-06 
0.0 0.396 0 -2.0 1e-06 
0.0 0.3961 0 -2.0 1e-06 
0.0 0.3962 0 -2.0 1e-06 
0.0 0.3963 0 -2.0 1e-06 
0.0 0.3964 0 -2.0 1e-06 
0.0 0.3965 0 -2.0 1e-06 
0.0 0.3966 0 -2.0 1e-06 
0.0 0.3967 0 -2.0 1e-06 
0.0 0.3968 0 -2.0 1e-06 
0.0 0.3969 0 -2.0 1e-06 
0.0 0.397 0 -2.0 1e-06 
0.0 0.3971 0 -2.0 1e-06 
0.0 0.3972 0 -2.0 1e-06 
0.0 0.3973 0 -2.0 1e-06 
0.0 0.3974 0 -2.0 1e-06 
0.0 0.3975 0 -2.0 1e-06 
0.0 0.3976 0 -2.0 1e-06 
0.0 0.3977 0 -2.0 1e-06 
0.0 0.3978 0 -2.0 1e-06 
0.0 0.3979 0 -2.0 1e-06 
0.0 0.398 0 -2.0 1e-06 
0.0 0.3981 0 -2.0 1e-06 
0.0 0.3982 0 -2.0 1e-06 
0.0 0.3983 0 -2.0 1e-06 
0.0 0.3984 0 -2.0 1e-06 
0.0 0.3985 0 -2.0 1e-06 
0.0 0.3986 0 -2.0 1e-06 
0.0 0.3987 0 -2.0 1e-06 
0.0 0.3988 0 -2.0 1e-06 
0.0 0.3989 0 -2.0 1e-06 
0.0 0.399 0 -2.0 1e-06 
0.0 0.3991 0 -2.0 1e-06 
0.0 0.3992 0 -2.0 1e-06 
0.0 0.3993 0 -2.0 1e-06 
0.0 0.3994 0 -2.0 1e-06 
0.0 0.3995 0 -2.0 1e-06 
0.0 0.3996 0 -2.0 1e-06 
0.0 0.3997 0 -2.0 1e-06 
0.0 0.3998 0 -2.0 1e-06 
0.0 0.3999 0 -2.0 1e-06 
0.0 0.4 0 -2.0 1e-06 
0.0 0.4001 0 -2.0 1e-06 
0.0 0.4002 0 -2.0 1e-06 
0.0 0.4003 0 -2.0 1e-06 
0.0 0.4004 0 -2.0 1e-06 
0.0 0.4005 0 -2.0 1e-06 
0.0 0.4006 0 -2.0 1e-06 
0.0 0.4007 0 -2.0 1e-06 
0.0 0.4008 0 -2.0 1e-06 
0.0 0.4009 0 -2.0 1e-06 
0.0 0.401 0 -2.0 1e-06 
0.0 0.4011 0 -2.0 1e-06 
0.0 0.4012 0 -2.0 1e-06 
0.0 0.4013 0 -2.0 1e-06 
0.0 0.4014 0 -2.0 1e-06 
0.0 0.4015 0 -2.0 1e-06 
0.0 0.4016 0 -2.0 1e-06 
0.0 0.4017 0 -2.0 1e-06 
0.0 0.4018 0 -2.0 1e-06 
0.0 0.4019 0 -2.0 1e-06 
0.0 0.402 0 -2.0 1e-06 
0.0 0.4021 0 -2.0 1e-06 
0.0 0.4022 0 -2.0 1e-06 
0.0 0.4023 0 -2.0 1e-06 
0.0 0.4024 0 -2.0 1e-06 
0.0 0.4025 0 -2.0 1e-06 
0.0 0.4026 0 -2.0 1e-06 
0.0 0.4027 0 -2.0 1e-06 
0.0 0.4028 0 -2.0 1e-06 
0.0 0.4029 0 -2.0 1e-06 
0.0 0.403 0 -2.0 1e-06 
0.0 0.4031 0 -2.0 1e-06 
0.0 0.4032 0 -2.0 1e-06 
0.0 0.4033 0 -2.0 1e-06 
0.0 0.4034 0 -2.0 1e-06 
0.0 0.4035 0 -2.0 1e-06 
0.0 0.4036 0 -2.0 1e-06 
0.0 0.4037 0 -2.0 1e-06 
0.0 0.4038 0 -2.0 1e-06 
0.0 0.4039 0 -2.0 1e-06 
0.0 0.404 0 -2.0 1e-06 
0.0 0.4041 0 -2.0 1e-06 
0.0 0.4042 0 -2.0 1e-06 
0.0 0.4043 0 -2.0 1e-06 
0.0 0.4044 0 -2.0 1e-06 
0.0 0.4045 0 -2.0 1e-06 
0.0 0.4046 0 -2.0 1e-06 
0.0 0.4047 0 -2.0 1e-06 
0.0 0.4048 0 -2.0 1e-06 
0.0 0.4049 0 -2.0 1e-06 
0.0 0.405 0 -2.0 1e-06 
0.0 0.4051 0 -2.0 1e-06 
0.0 0.4052 0 -2.0 1e-06 
0.0 0.4053 0 -2.0 1e-06 
0.0 0.4054 0 -2.0 1e-06 
0.0 0.4055 0 -2.0 1e-06 
0.0 0.4056 0 -2.0 1e-06 
0.0 0.4057 0 -2.0 1e-06 
0.0 0.4058 0 -2.0 1e-06 
0.0 0.4059 0 -2.0 1e-06 
0.0 0.406 0 -2.0 1e-06 
0.0 0.4061 0 -2.0 1e-06 
0.0 0.4062 0 -2.0 1e-06 
0.0 0.4063 0 -2.0 1e-06 
0.0 0.4064 0 -2.0 1e-06 
0.0 0.4065 0 -2.0 1e-06 
0.0 0.4066 0 -2.0 1e-06 
0.0 0.4067 0 -2.0 1e-06 
0.0 0.4068 0 -2.0 1e-06 
0.0 0.4069 0 -2.0 1e-06 
0.0 0.407 0 -2.0 1e-06 
0.0 0.4071 0 -2.0 1e-06 
0.0 0.4072 0 -2.0 1e-06 
0.0 0.4073 0 -2.0 1e-06 
0.0 0.4074 0 -2.0 1e-06 
0.0 0.4075 0 -2.0 1e-06 
0.0 0.4076 0 -2.0 1e-06 
0.0 0.4077 0 -2.0 1e-06 
0.0 0.4078 0 -2.0 1e-06 
0.0 0.4079 0 -2.0 1e-06 
0.0 0.408 0 -2.0 1e-06 
0.0 0.4081 0 -2.0 1e-06 
0.0 0.4082 0 -2.0 1e-06 
0.0 0.4083 0 -2.0 1e-06 
0.0 0.4084 0 -2.0 1e-06 
0.0 0.4085 0 -2.0 1e-06 
0.0 0.4086 0 -2.0 1e-06 
0.0 0.4087 0 -2.0 1e-06 
0.0 0.4088 0 -2.0 1e-06 
0.0 0.4089 0 -2.0 1e-06 
0.0 0.409 0 -2.0 1e-06 
0.0 0.4091 0 -2.0 1e-06 
0.0 0.4092 0 -2.0 1e-06 
0.0 0.4093 0 -2.0 1e-06 
0.0 0.4094 0 -2.0 1e-06 
0.0 0.4095 0 -2.0 1e-06 
0.0 0.4096 0 -2.0 1e-06 
0.0 0.4097 0 -2.0 1e-06 
0.0 0.4098 0 -2.0 1e-06 
0.0 0.4099 0 -2.0 1e-06 
0.0 0.41 0 -2.0 1e-06 
0.0 0.4101 0 -2.0 1e-06 
0.0 0.4102 0 -2.0 1e-06 
0.0 0.4103 0 -2.0 1e-06 
0.0 0.4104 0 -2.0 1e-06 
0.0 0.4105 0 -2.0 1e-06 
0.0 0.4106 0 -2.0 1e-06 
0.0 0.4107 0 -2.0 1e-06 
0.0 0.4108 0 -2.0 1e-06 
0.0 0.4109 0 -2.0 1e-06 
0.0 0.411 0 -2.0 1e-06 
0.0 0.4111 0 -2.0 1e-06 
0.0 0.4112 0 -2.0 1e-06 
0.0 0.4113 0 -2.0 1e-06 
0.0 0.4114 0 -2.0 1e-06 
0.0 0.4115 0 -2.0 1e-06 
0.0 0.4116 0 -2.0 1e-06 
0.0 0.4117 0 -2.0 1e-06 
0.0 0.4118 0 -2.0 1e-06 
0.0 0.4119 0 -2.0 1e-06 
0.0 0.412 0 -2.0 1e-06 
0.0 0.4121 0 -2.0 1e-06 
0.0 0.4122 0 -2.0 1e-06 
0.0 0.4123 0 -2.0 1e-06 
0.0 0.4124 0 -2.0 1e-06 
0.0 0.4125 0 -2.0 1e-06 
0.0 0.4126 0 -2.0 1e-06 
0.0 0.4127 0 -2.0 1e-06 
0.0 0.4128 0 -2.0 1e-06 
0.0 0.4129 0 -2.0 1e-06 
0.0 0.413 0 -2.0 1e-06 
0.0 0.4131 0 -2.0 1e-06 
0.0 0.4132 0 -2.0 1e-06 
0.0 0.4133 0 -2.0 1e-06 
0.0 0.4134 0 -2.0 1e-06 
0.0 0.4135 0 -2.0 1e-06 
0.0 0.4136 0 -2.0 1e-06 
0.0 0.4137 0 -2.0 1e-06 
0.0 0.4138 0 -2.0 1e-06 
0.0 0.4139 0 -2.0 1e-06 
0.0 0.414 0 -2.0 1e-06 
0.0 0.4141 0 -2.0 1e-06 
0.0 0.4142 0 -2.0 1e-06 
0.0 0.4143 0 -2.0 1e-06 
0.0 0.4144 0 -2.0 1e-06 
0.0 0.4145 0 -2.0 1e-06 
0.0 0.4146 0 -2.0 1e-06 
0.0 0.4147 0 -2.0 1e-06 
0.0 0.4148 0 -2.0 1e-06 
0.0 0.4149 0 -2.0 1e-06 
0.0 0.415 0 -2.0 1e-06 
0.0 0.4151 0 -2.0 1e-06 
0.0 0.4152 0 -2.0 1e-06 
0.0 0.4153 0 -2.0 1e-06 
0.0 0.4154 0 -2.0 1e-06 
0.0 0.4155 0 -2.0 1e-06 
0.0 0.4156 0 -2.0 1e-06 
0.0 0.4157 0 -2.0 1e-06 
0.0 0.4158 0 -2.0 1e-06 
0.0 0.4159 0 -2.0 1e-06 
0.0 0.416 0 -2.0 1e-06 
0.0 0.4161 0 -2.0 1e-06 
0.0 0.4162 0 -2.0 1e-06 
0.0 0.4163 0 -2.0 1e-06 
0.0 0.4164 0 -2.0 1e-06 
0.0 0.4165 0 -2.0 1e-06 
0.0 0.4166 0 -2.0 1e-06 
0.0 0.4167 0 -2.0 1e-06 
0.0 0.4168 0 -2.0 1e-06 
0.0 0.4169 0 -2.0 1e-06 
0.0 0.417 0 -2.0 1e-06 
0.0 0.4171 0 -2.0 1e-06 
0.0 0.4172 0 -2.0 1e-06 
0.0 0.4173 0 -2.0 1e-06 
0.0 0.4174 0 -2.0 1e-06 
0.0 0.4175 0 -2.0 1e-06 
0.0 0.4176 0 -2.0 1e-06 
0.0 0.4177 0 -2.0 1e-06 
0.0 0.4178 0 -2.0 1e-06 
0.0 0.4179 0 -2.0 1e-06 
0.0 0.418 0 -2.0 1e-06 
0.0 0.4181 0 -2.0 1e-06 
0.0 0.4182 0 -2.0 1e-06 
0.0 0.4183 0 -2.0 1e-06 
0.0 0.4184 0 -2.0 1e-06 
0.0 0.4185 0 -2.0 1e-06 
0.0 0.4186 0 -2.0 1e-06 
0.0 0.4187 0 -2.0 1e-06 
0.0 0.4188 0 -2.0 1e-06 
0.0 0.4189 0 -2.0 1e-06 
0.0 0.419 0 -2.0 1e-06 
0.0 0.4191 0 -2.0 1e-06 
0.0 0.4192 0 -2.0 1e-06 
0.0 0.4193 0 -2.0 1e-06 
0.0 0.4194 0 -2.0 1e-06 
0.0 0.4195 0 -2.0 1e-06 
0.0 0.4196 0 -2.0 1e-06 
0.0 0.4197 0 -2.0 1e-06 
0.0 0.4198 0 -2.0 1e-06 
0.0 0.4199 0 -2.0 1e-06 
0.0 0.42 0 -2.0 1e-06 
0.0 0.4201 0 -2.0 1e-06 
0.0 0.4202 0 -2.0 1e-06 
0.0 0.4203 0 -2.0 1e-06 
0.0 0.4204 0 -2.0 1e-06 
0.0 0.4205 0 -2.0 1e-06 
0.0 0.4206 0 -2.0 1e-06 
0.0 0.4207 0 -2.0 1e-06 
0.0 0.4208 0 -2.0 1e-06 
0.0 0.4209 0 -2.0 1e-06 
0.0 0.421 0 -2.0 1e-06 
0.0 0.4211 0 -2.0 1e-06 
0.0 0.4212 0 -2.0 1e-06 
0.0 0.4213 0 -2.0 1e-06 
0.0 0.4214 0 -2.0 1e-06 
0.0 0.4215 0 -2.0 1e-06 
0.0 0.4216 0 -2.0 1e-06 
0.0 0.4217 0 -2.0 1e-06 
0.0 0.4218 0 -2.0 1e-06 
0.0 0.4219 0 -2.0 1e-06 
0.0 0.422 0 -2.0 1e-06 
0.0 0.4221 0 -2.0 1e-06 
0.0 0.4222 0 -2.0 1e-06 
0.0 0.4223 0 -2.0 1e-06 
0.0 0.4224 0 -2.0 1e-06 
0.0 0.4225 0 -2.0 1e-06 
0.0 0.4226 0 -2.0 1e-06 
0.0 0.4227 0 -2.0 1e-06 
0.0 0.4228 0 -2.0 1e-06 
0.0 0.4229 0 -2.0 1e-06 
0.0 0.423 0 -2.0 1e-06 
0.0 0.4231 0 -2.0 1e-06 
0.0 0.4232 0 -2.0 1e-06 
0.0 0.4233 0 -2.0 1e-06 
0.0 0.4234 0 -2.0 1e-06 
0.0 0.4235 0 -2.0 1e-06 
0.0 0.4236 0 -2.0 1e-06 
0.0 0.4237 0 -2.0 1e-06 
0.0 0.4238 0 -2.0 1e-06 
0.0 0.4239 0 -2.0 1e-06 
0.0 0.424 0 -2.0 1e-06 
0.0 0.4241 0 -2.0 1e-06 
0.0 0.4242 0 -2.0 1e-06 
0.0 0.4243 0 -2.0 1e-06 
0.0 0.4244 0 -2.0 1e-06 
0.0 0.4245 0 -2.0 1e-06 
0.0 0.4246 0 -2.0 1e-06 
0.0 0.4247 0 -2.0 1e-06 
0.0 0.4248 0 -2.0 1e-06 
0.0 0.4249 0 -2.0 1e-06 
0.0 0.425 0 -2.0 1e-06 
0.0 0.4251 0 -2.0 1e-06 
0.0 0.4252 0 -2.0 1e-06 
0.0 0.4253 0 -2.0 1e-06 
0.0 0.4254 0 -2.0 1e-06 
0.0 0.4255 0 -2.0 1e-06 
0.0 0.4256 0 -2.0 1e-06 
0.0 0.4257 0 -2.0 1e-06 
0.0 0.4258 0 -2.0 1e-06 
0.0 0.4259 0 -2.0 1e-06 
0.0 0.426 0 -2.0 1e-06 
0.0 0.4261 0 -2.0 1e-06 
0.0 0.4262 0 -2.0 1e-06 
0.0 0.4263 0 -2.0 1e-06 
0.0 0.4264 0 -2.0 1e-06 
0.0 0.4265 0 -2.0 1e-06 
0.0 0.4266 0 -2.0 1e-06 
0.0 0.4267 0 -2.0 1e-06 
0.0 0.4268 0 -2.0 1e-06 
0.0 0.4269 0 -2.0 1e-06 
0.0 0.427 0 -2.0 1e-06 
0.0 0.4271 0 -2.0 1e-06 
0.0 0.4272 0 -2.0 1e-06 
0.0 0.4273 0 -2.0 1e-06 
0.0 0.4274 0 -2.0 1e-06 
0.0 0.4275 0 -2.0 1e-06 
0.0 0.4276 0 -2.0 1e-06 
0.0 0.4277 0 -2.0 1e-06 
0.0 0.4278 0 -2.0 1e-06 
0.0 0.4279 0 -2.0 1e-06 
0.0 0.428 0 -2.0 1e-06 
0.0 0.4281 0 -2.0 1e-06 
0.0 0.4282 0 -2.0 1e-06 
0.0 0.4283 0 -2.0 1e-06 
0.0 0.4284 0 -2.0 1e-06 
0.0 0.4285 0 -2.0 1e-06 
0.0 0.4286 0 -2.0 1e-06 
0.0 0.4287 0 -2.0 1e-06 
0.0 0.4288 0 -2.0 1e-06 
0.0 0.4289 0 -2.0 1e-06 
0.0 0.429 0 -2.0 1e-06 
0.0 0.4291 0 -2.0 1e-06 
0.0 0.4292 0 -2.0 1e-06 
0.0 0.4293 0 -2.0 1e-06 
0.0 0.4294 0 -2.0 1e-06 
0.0 0.4295 0 -2.0 1e-06 
0.0 0.4296 0 -2.0 1e-06 
0.0 0.4297 0 -2.0 1e-06 
0.0 0.4298 0 -2.0 1e-06 
0.0 0.4299 0 -2.0 1e-06 
0.0 0.43 0 -2.0 1e-06 
0.0 0.4301 0 -2.0 1e-06 
0.0 0.4302 0 -2.0 1e-06 
0.0 0.4303 0 -2.0 1e-06 
0.0 0.4304 0 -2.0 1e-06 
0.0 0.4305 0 -2.0 1e-06 
0.0 0.4306 0 -2.0 1e-06 
0.0 0.4307 0 -2.0 1e-06 
0.0 0.4308 0 -2.0 1e-06 
0.0 0.4309 0 -2.0 1e-06 
0.0 0.431 0 -2.0 1e-06 
0.0 0.4311 0 -2.0 1e-06 
0.0 0.4312 0 -2.0 1e-06 
0.0 0.4313 0 -2.0 1e-06 
0.0 0.4314 0 -2.0 1e-06 
0.0 0.4315 0 -2.0 1e-06 
0.0 0.4316 0 -2.0 1e-06 
0.0 0.4317 0 -2.0 1e-06 
0.0 0.4318 0 -2.0 1e-06 
0.0 0.4319 0 -2.0 1e-06 
0.0 0.432 0 -2.0 1e-06 
0.0 0.4321 0 -2.0 1e-06 
0.0 0.4322 0 -2.0 1e-06 
0.0 0.4323 0 -2.0 1e-06 
0.0 0.4324 0 -2.0 1e-06 
0.0 0.4325 0 -2.0 1e-06 
0.0 0.4326 0 -2.0 1e-06 
0.0 0.4327 0 -2.0 1e-06 
0.0 0.4328 0 -2.0 1e-06 
0.0 0.4329 0 -2.0 1e-06 
0.0 0.433 0 -2.0 1e-06 
0.0 0.4331 0 -2.0 1e-06 
0.0 0.4332 0 -2.0 1e-06 
0.0 0.4333 0 -2.0 1e-06 
0.0 0.4334 0 -2.0 1e-06 
0.0 0.4335 0 -2.0 1e-06 
0.0 0.4336 0 -2.0 1e-06 
0.0 0.4337 0 -2.0 1e-06 
0.0 0.4338 0 -2.0 1e-06 
0.0 0.4339 0 -2.0 1e-06 
0.0 0.434 0 -2.0 1e-06 
0.0 0.4341 0 -2.0 1e-06 
0.0 0.4342 0 -2.0 1e-06 
0.0 0.4343 0 -2.0 1e-06 
0.0 0.4344 0 -2.0 1e-06 
0.0 0.4345 0 -2.0 1e-06 
0.0 0.4346 0 -2.0 1e-06 
0.0 0.4347 0 -2.0 1e-06 
0.0 0.4348 0 -2.0 1e-06 
0.0 0.4349 0 -2.0 1e-06 
0.0 0.435 0 -2.0 1e-06 
0.0 0.4351 0 -2.0 1e-06 
0.0 0.4352 0 -2.0 1e-06 
0.0 0.4353 0 -2.0 1e-06 
0.0 0.4354 0 -2.0 1e-06 
0.0 0.4355 0 -2.0 1e-06 
0.0 0.4356 0 -2.0 1e-06 
0.0 0.4357 0 -2.0 1e-06 
0.0 0.4358 0 -2.0 1e-06 
0.0 0.4359 0 -2.0 1e-06 
0.0 0.436 0 -2.0 1e-06 
0.0 0.4361 0 -2.0 1e-06 
0.0 0.4362 0 -2.0 1e-06 
0.0 0.4363 0 -2.0 1e-06 
0.0 0.4364 0 -2.0 1e-06 
0.0 0.4365 0 -2.0 1e-06 
0.0 0.4366 0 -2.0 1e-06 
0.0 0.4367 0 -2.0 1e-06 
0.0 0.4368 0 -2.0 1e-06 
0.0 0.4369 0 -2.0 1e-06 
0.0 0.437 0 -2.0 1e-06 
0.0 0.4371 0 -2.0 1e-06 
0.0 0.4372 0 -2.0 1e-06 
0.0 0.4373 0 -2.0 1e-06 
0.0 0.4374 0 -2.0 1e-06 
0.0 0.4375 0 -2.0 1e-06 
0.0 0.4376 0 -2.0 1e-06 
0.0 0.4377 0 -2.0 1e-06 
0.0 0.4378 0 -2.0 1e-06 
0.0 0.4379 0 -2.0 1e-06 
0.0 0.438 0 -2.0 1e-06 
0.0 0.4381 0 -2.0 1e-06 
0.0 0.4382 0 -2.0 1e-06 
0.0 0.4383 0 -2.0 1e-06 
0.0 0.4384 0 -2.0 1e-06 
0.0 0.4385 0 -2.0 1e-06 
0.0 0.4386 0 -2.0 1e-06 
0.0 0.4387 0 -2.0 1e-06 
0.0 0.4388 0 -2.0 1e-06 
0.0 0.4389 0 -2.0 1e-06 
0.0 0.439 0 -2.0 1e-06 
0.0 0.4391 0 -2.0 1e-06 
0.0 0.4392 0 -2.0 1e-06 
0.0 0.4393 0 -2.0 1e-06 
0.0 0.4394 0 -2.0 1e-06 
0.0 0.4395 0 -2.0 1e-06 
0.0 0.4396 0 -2.0 1e-06 
0.0 0.4397 0 -2.0 1e-06 
0.0 0.4398 0 -2.0 1e-06 
0.0 0.4399 0 -2.0 1e-06 
0.0 0.44 0 -2.0 1e-06 
0.0 0.4401 0 -2.0 1e-06 
0.0 0.4402 0 -2.0 1e-06 
0.0 0.4403 0 -2.0 1e-06 
0.0 0.4404 0 -2.0 1e-06 
0.0 0.4405 0 -2.0 1e-06 
0.0 0.4406 0 -2.0 1e-06 
0.0 0.4407 0 -2.0 1e-06 
0.0 0.4408 0 -2.0 1e-06 
0.0 0.4409 0 -2.0 1e-06 
0.0 0.441 0 -2.0 1e-06 
0.0 0.4411 0 -2.0 1e-06 
0.0 0.4412 0 -2.0 1e-06 
0.0 0.4413 0 -2.0 1e-06 
0.0 0.4414 0 -2.0 1e-06 
0.0 0.4415 0 -2.0 1e-06 
0.0 0.4416 0 -2.0 1e-06 
0.0 0.4417 0 -2.0 1e-06 
0.0 0.4418 0 -2.0 1e-06 
0.0 0.4419 0 -2.0 1e-06 
0.0 0.442 0 -2.0 1e-06 
0.0 0.4421 0 -2.0 1e-06 
0.0 0.4422 0 -2.0 1e-06 
0.0 0.4423 0 -2.0 1e-06 
0.0 0.4424 0 -2.0 1e-06 
0.0 0.4425 0 -2.0 1e-06 
0.0 0.4426 0 -2.0 1e-06 
0.0 0.4427 0 -2.0 1e-06 
0.0 0.4428 0 -2.0 1e-06 
0.0 0.4429 0 -2.0 1e-06 
0.0 0.443 0 -2.0 1e-06 
0.0 0.4431 0 -2.0 1e-06 
0.0 0.4432 0 -2.0 1e-06 
0.0 0.4433 0 -2.0 1e-06 
0.0 0.4434 0 -2.0 1e-06 
0.0 0.4435 0 -2.0 1e-06 
0.0 0.4436 0 -2.0 1e-06 
0.0 0.4437 0 -2.0 1e-06 
0.0 0.4438 0 -2.0 1e-06 
0.0 0.4439 0 -2.0 1e-06 
0.0 0.444 0 -2.0 1e-06 
0.0 0.4441 0 -2.0 1e-06 
0.0 0.4442 0 -2.0 1e-06 
0.0 0.4443 0 -2.0 1e-06 
0.0 0.4444 0 -2.0 1e-06 
0.0 0.4445 0 -2.0 1e-06 
0.0 0.4446 0 -2.0 1e-06 
0.0 0.4447 0 -2.0 1e-06 
0.0 0.4448 0 -2.0 1e-06 
0.0 0.4449 0 -2.0 1e-06 
0.0 0.445 0 -2.0 1e-06 
0.0 0.4451 0 -2.0 1e-06 
0.0 0.4452 0 -2.0 1e-06 
0.0 0.4453 0 -2.0 1e-06 
0.0 0.4454 0 -2.0 1e-06 
0.0 0.4455 0 -2.0 1e-06 
0.0 0.4456 0 -2.0 1e-06 
0.0 0.4457 0 -2.0 1e-06 
0.0 0.4458 0 -2.0 1e-06 
0.0 0.4459 0 -2.0 1e-06 
0.0 0.446 0 -2.0 1e-06 
0.0 0.4461 0 -2.0 1e-06 
0.0 0.4462 0 -2.0 1e-06 
0.0 0.4463 0 -2.0 1e-06 
0.0 0.4464 0 -2.0 1e-06 
0.0 0.4465 0 -2.0 1e-06 
0.0 0.4466 0 -2.0 1e-06 
0.0 0.4467 0 -2.0 1e-06 
0.0 0.4468 0 -2.0 1e-06 
0.0 0.4469 0 -2.0 1e-06 
0.0 0.447 0 -2.0 1e-06 
0.0 0.4471 0 -2.0 1e-06 
0.0 0.4472 0 -2.0 1e-06 
0.0 0.4473 0 -2.0 1e-06 
0.0 0.4474 0 -2.0 1e-06 
0.0 0.4475 0 -2.0 1e-06 
0.0 0.4476 0 -2.0 1e-06 
0.0 0.4477 0 -2.0 1e-06 
0.0 0.4478 0 -2.0 1e-06 
0.0 0.4479 0 -2.0 1e-06 
0.0 0.448 0 -2.0 1e-06 
0.0 0.4481 0 -2.0 1e-06 
0.0 0.4482 0 -2.0 1e-06 
0.0 0.4483 0 -2.0 1e-06 
0.0 0.4484 0 -2.0 1e-06 
0.0 0.4485 0 -2.0 1e-06 
0.0 0.4486 0 -2.0 1e-06 
0.0 0.4487 0 -2.0 1e-06 
0.0 0.4488 0 -2.0 1e-06 
0.0 0.4489 0 -2.0 1e-06 
0.0 0.449 0 -2.0 1e-06 
0.0 0.4491 0 -2.0 1e-06 
0.0 0.4492 0 -2.0 1e-06 
0.0 0.4493 0 -2.0 1e-06 
0.0 0.4494 0 -2.0 1e-06 
0.0 0.4495 0 -2.0 1e-06 
0.0 0.4496 0 -2.0 1e-06 
0.0 0.4497 0 -2.0 1e-06 
0.0 0.4498 0 -2.0 1e-06 
0.0 0.4499 0 -2.0 1e-06 
0.0 0.45 0 -2.0 1e-06 
0.0 0.4501 0 -2.0 1e-06 
0.0 0.4502 0 -2.0 1e-06 
0.0 0.4503 0 -2.0 1e-06 
0.0 0.4504 0 -2.0 1e-06 
0.0 0.4505 0 -2.0 1e-06 
0.0 0.4506 0 -2.0 1e-06 
0.0 0.4507 0 -2.0 1e-06 
0.0 0.4508 0 -2.0 1e-06 
0.0 0.4509 0 -2.0 1e-06 
0.0 0.451 0 -2.0 1e-06 
0.0 0.4511 0 -2.0 1e-06 
0.0 0.4512 0 -2.0 1e-06 
0.0 0.4513 0 -2.0 1e-06 
0.0 0.4514 0 -2.0 1e-06 
0.0 0.4515 0 -2.0 1e-06 
0.0 0.4516 0 -2.0 1e-06 
0.0 0.4517 0 -2.0 1e-06 
0.0 0.4518 0 -2.0 1e-06 
0.0 0.4519 0 -2.0 1e-06 
0.0 0.452 0 -2.0 1e-06 
0.0 0.4521 0 -2.0 1e-06 
0.0 0.4522 0 -2.0 1e-06 
0.0 0.4523 0 -2.0 1e-06 
0.0 0.4524 0 -2.0 1e-06 
0.0 0.4525 0 -2.0 1e-06 
0.0 0.4526 0 -2.0 1e-06 
0.0 0.4527 0 -2.0 1e-06 
0.0 0.4528 0 -2.0 1e-06 
0.0 0.4529 0 -2.0 1e-06 
0.0 0.453 0 -2.0 1e-06 
0.0 0.4531 0 -2.0 1e-06 
0.0 0.4532 0 -2.0 1e-06 
0.0 0.4533 0 -2.0 1e-06 
0.0 0.4534 0 -2.0 1e-06 
0.0 0.4535 0 -2.0 1e-06 
0.0 0.4536 0 -2.0 1e-06 
0.0 0.4537 0 -2.0 1e-06 
0.0 0.4538 0 -2.0 1e-06 
0.0 0.4539 0 -2.0 1e-06 
0.0 0.454 0 -2.0 1e-06 
0.0 0.4541 0 -2.0 1e-06 
0.0 0.4542 0 -2.0 1e-06 
0.0 0.4543 0 -2.0 1e-06 
0.0 0.4544 0 -2.0 1e-06 
0.0 0.4545 0 -2.0 1e-06 
0.0 0.4546 0 -2.0 1e-06 
0.0 0.4547 0 -2.0 1e-06 
0.0 0.4548 0 -2.0 1e-06 
0.0 0.4549 0 -2.0 1e-06 
0.0 0.455 0 -2.0 1e-06 
0.0 0.4551 0 -2.0 1e-06 
0.0 0.4552 0 -2.0 1e-06 
0.0 0.4553 0 -2.0 1e-06 
0.0 0.4554 0 -2.0 1e-06 
0.0 0.4555 0 -2.0 1e-06 
0.0 0.4556 0 -2.0 1e-06 
0.0 0.4557 0 -2.0 1e-06 
0.0 0.4558 0 -2.0 1e-06 
0.0 0.4559 0 -2.0 1e-06 
0.0 0.456 0 -2.0 1e-06 
0.0 0.4561 0 -2.0 1e-06 
0.0 0.4562 0 -2.0 1e-06 
0.0 0.4563 0 -2.0 1e-06 
0.0 0.4564 0 -2.0 1e-06 
0.0 0.4565 0 -2.0 1e-06 
0.0 0.4566 0 -2.0 1e-06 
0.0 0.4567 0 -2.0 1e-06 
0.0 0.4568 0 -2.0 1e-06 
0.0 0.4569 0 -2.0 1e-06 
0.0 0.457 0 -2.0 1e-06 
0.0 0.4571 0 -2.0 1e-06 
0.0 0.4572 0 -2.0 1e-06 
0.0 0.4573 0 -2.0 1e-06 
0.0 0.4574 0 -2.0 1e-06 
0.0 0.4575 0 -2.0 1e-06 
0.0 0.4576 0 -2.0 1e-06 
0.0 0.4577 0 -2.0 1e-06 
0.0 0.4578 0 -2.0 1e-06 
0.0 0.4579 0 -2.0 1e-06 
0.0 0.458 0 -2.0 1e-06 
0.0 0.4581 0 -2.0 1e-06 
0.0 0.4582 0 -2.0 1e-06 
0.0 0.4583 0 -2.0 1e-06 
0.0 0.4584 0 -2.0 1e-06 
0.0 0.4585 0 -2.0 1e-06 
0.0 0.4586 0 -2.0 1e-06 
0.0 0.4587 0 -2.0 1e-06 
0.0 0.4588 0 -2.0 1e-06 
0.0 0.4589 0 -2.0 1e-06 
0.0 0.459 0 -2.0 1e-06 
0.0 0.4591 0 -2.0 1e-06 
0.0 0.4592 0 -2.0 1e-06 
0.0 0.4593 0 -2.0 1e-06 
0.0 0.4594 0 -2.0 1e-06 
0.0 0.4595 0 -2.0 1e-06 
0.0 0.4596 0 -2.0 1e-06 
0.0 0.4597 0 -2.0 1e-06 
0.0 0.4598 0 -2.0 1e-06 
0.0 0.4599 0 -2.0 1e-06 
0.0 0.46 0 -2.0 1e-06 
0.0 0.4601 0 -2.0 1e-06 
0.0 0.4602 0 -2.0 1e-06 
0.0 0.4603 0 -2.0 1e-06 
0.0 0.4604 0 -2.0 1e-06 
0.0 0.4605 0 -2.0 1e-06 
0.0 0.4606 0 -2.0 1e-06 
0.0 0.4607 0 -2.0 1e-06 
0.0 0.4608 0 -2.0 1e-06 
0.0 0.4609 0 -2.0 1e-06 
0.0 0.461 0 -2.0 1e-06 
0.0 0.4611 0 -2.0 1e-06 
0.0 0.4612 0 -2.0 1e-06 
0.0 0.4613 0 -2.0 1e-06 
0.0 0.4614 0 -2.0 1e-06 
0.0 0.4615 0 -2.0 1e-06 
0.0 0.4616 0 -2.0 1e-06 
0.0 0.4617 0 -2.0 1e-06 
0.0 0.4618 0 -2.0 1e-06 
0.0 0.4619 0 -2.0 1e-06 
0.0 0.462 0 -2.0 1e-06 
0.0 0.4621 0 -2.0 1e-06 
0.0 0.4622 0 -2.0 1e-06 
0.0 0.4623 0 -2.0 1e-06 
0.0 0.4624 0 -2.0 1e-06 
0.0 0.4625 0 -2.0 1e-06 
0.0 0.4626 0 -2.0 1e-06 
0.0 0.4627 0 -2.0 1e-06 
0.0 0.4628 0 -2.0 1e-06 
0.0 0.4629 0 -2.0 1e-06 
0.0 0.463 0 -2.0 1e-06 
0.0 0.4631 0 -2.0 1e-06 
0.0 0.4632 0 -2.0 1e-06 
0.0 0.4633 0 -2.0 1e-06 
0.0 0.4634 0 -2.0 1e-06 
0.0 0.4635 0 -2.0 1e-06 
0.0 0.4636 0 -2.0 1e-06 
0.0 0.4637 0 -2.0 1e-06 
0.0 0.4638 0 -2.0 1e-06 
0.0 0.4639 0 -2.0 1e-06 
0.0 0.464 0 -2.0 1e-06 
0.0 0.4641 0 -2.0 1e-06 
0.0 0.4642 0 -2.0 1e-06 
0.0 0.4643 0 -2.0 1e-06 
0.0 0.4644 0 -2.0 1e-06 
0.0 0.4645 0 -2.0 1e-06 
0.0 0.4646 0 -2.0 1e-06 
0.0 0.4647 0 -2.0 1e-06 
0.0 0.4648 0 -2.0 1e-06 
0.0 0.4649 0 -2.0 1e-06 
0.0 0.465 0 -2.0 1e-06 
0.0 0.4651 0 -2.0 1e-06 
0.0 0.4652 0 -2.0 1e-06 
0.0 0.4653 0 -2.0 1e-06 
0.0 0.4654 0 -2.0 1e-06 
0.0 0.4655 0 -2.0 1e-06 
0.0 0.4656 0 -2.0 1e-06 
0.0 0.4657 0 -2.0 1e-06 
0.0 0.4658 0 -2.0 1e-06 
0.0 0.4659 0 -2.0 1e-06 
0.0 0.466 0 -2.0 1e-06 
0.0 0.4661 0 -2.0 1e-06 
0.0 0.4662 0 -2.0 1e-06 
0.0 0.4663 0 -2.0 1e-06 
0.0 0.4664 0 -2.0 1e-06 
0.0 0.4665 0 -2.0 1e-06 
0.0 0.4666 0 -2.0 1e-06 
0.0 0.4667 0 -2.0 1e-06 
0.0 0.4668 0 -2.0 1e-06 
0.0 0.4669 0 -2.0 1e-06 
0.0 0.467 0 -2.0 1e-06 
0.0 0.4671 0 -2.0 1e-06 
0.0 0.4672 0 -2.0 1e-06 
0.0 0.4673 0 -2.0 1e-06 
0.0 0.4674 0 -2.0 1e-06 
0.0 0.4675 0 -2.0 1e-06 
0.0 0.4676 0 -2.0 1e-06 
0.0 0.4677 0 -2.0 1e-06 
0.0 0.4678 0 -2.0 1e-06 
0.0 0.4679 0 -2.0 1e-06 
0.0 0.468 0 -2.0 1e-06 
0.0 0.4681 0 -2.0 1e-06 
0.0 0.4682 0 -2.0 1e-06 
0.0 0.4683 0 -2.0 1e-06 
0.0 0.4684 0 -2.0 1e-06 
0.0 0.4685 0 -2.0 1e-06 
0.0 0.4686 0 -2.0 1e-06 
0.0 0.4687 0 -2.0 1e-06 
0.0 0.4688 0 -2.0 1e-06 
0.0 0.4689 0 -2.0 1e-06 
0.0 0.469 0 -2.0 1e-06 
0.0 0.4691 0 -2.0 1e-06 
0.0 0.4692 0 -2.0 1e-06 
0.0 0.4693 0 -2.0 1e-06 
0.0 0.4694 0 -2.0 1e-06 
0.0 0.4695 0 -2.0 1e-06 
0.0 0.4696 0 -2.0 1e-06 
0.0 0.4697 0 -2.0 1e-06 
0.0 0.4698 0 -2.0 1e-06 
0.0 0.4699 0 -2.0 1e-06 
0.0 0.47 0 -2.0 1e-06 
0.0 0.4701 0 -2.0 1e-06 
0.0 0.4702 0 -2.0 1e-06 
0.0 0.4703 0 -2.0 1e-06 
0.0 0.4704 0 -2.0 1e-06 
0.0 0.4705 0 -2.0 1e-06 
0.0 0.4706 0 -2.0 1e-06 
0.0 0.4707 0 -2.0 1e-06 
0.0 0.4708 0 -2.0 1e-06 
0.0 0.4709 0 -2.0 1e-06 
0.0 0.471 0 -2.0 1e-06 
0.0 0.4711 0 -2.0 1e-06 
0.0 0.4712 0 -2.0 1e-06 
0.0 0.4713 0 -2.0 1e-06 
0.0 0.4714 0 -2.0 1e-06 
0.0 0.4715 0 -2.0 1e-06 
0.0 0.4716 0 -2.0 1e-06 
0.0 0.4717 0 -2.0 1e-06 
0.0 0.4718 0 -2.0 1e-06 
0.0 0.4719 0 -2.0 1e-06 
0.0 0.472 0 -2.0 1e-06 
0.0 0.4721 0 -2.0 1e-06 
0.0 0.4722 0 -2.0 1e-06 
0.0 0.4723 0 -2.0 1e-06 
0.0 0.4724 0 -2.0 1e-06 
0.0 0.4725 0 -2.0 1e-06 
0.0 0.4726 0 -2.0 1e-06 
0.0 0.4727 0 -2.0 1e-06 
0.0 0.4728 0 -2.0 1e-06 
0.0 0.4729 0 -2.0 1e-06 
0.0 0.473 0 -2.0 1e-06 
0.0 0.4731 0 -2.0 1e-06 
0.0 0.4732 0 -2.0 1e-06 
0.0 0.4733 0 -2.0 1e-06 
0.0 0.4734 0 -2.0 1e-06 
0.0 0.4735 0 -2.0 1e-06 
0.0 0.4736 0 -2.0 1e-06 
0.0 0.4737 0 -2.0 1e-06 
0.0 0.4738 0 -2.0 1e-06 
0.0 0.4739 0 -2.0 1e-06 
0.0 0.474 0 -2.0 1e-06 
0.0 0.4741 0 -2.0 1e-06 
0.0 0.4742 0 -2.0 1e-06 
0.0 0.4743 0 -2.0 1e-06 
0.0 0.4744 0 -2.0 1e-06 
0.0 0.4745 0 -2.0 1e-06 
0.0 0.4746 0 -2.0 1e-06 
0.0 0.4747 0 -2.0 1e-06 
0.0 0.4748 0 -2.0 1e-06 
0.0 0.4749 0 -2.0 1e-06 
0.0 0.475 0 -2.0 1e-06 
0.0 0.4751 0 -2.0 1e-06 
0.0 0.4752 0 -2.0 1e-06 
0.0 0.4753 0 -2.0 1e-06 
0.0 0.4754 0 -2.0 1e-06 
0.0 0.4755 0 -2.0 1e-06 
0.0 0.4756 0 -2.0 1e-06 
0.0 0.4757 0 -2.0 1e-06 
0.0 0.4758 0 -2.0 1e-06 
0.0 0.4759 0 -2.0 1e-06 
0.0 0.476 0 -2.0 1e-06 
0.0 0.4761 0 -2.0 1e-06 
0.0 0.4762 0 -2.0 1e-06 
0.0 0.4763 0 -2.0 1e-06 
0.0 0.4764 0 -2.0 1e-06 
0.0 0.4765 0 -2.0 1e-06 
0.0 0.4766 0 -2.0 1e-06 
0.0 0.4767 0 -2.0 1e-06 
0.0 0.4768 0 -2.0 1e-06 
0.0 0.4769 0 -2.0 1e-06 
0.0 0.477 0 -2.0 1e-06 
0.0 0.4771 0 -2.0 1e-06 
0.0 0.4772 0 -2.0 1e-06 
0.0 0.4773 0 -2.0 1e-06 
0.0 0.4774 0 -2.0 1e-06 
0.0 0.4775 0 -2.0 1e-06 
0.0 0.4776 0 -2.0 1e-06 
0.0 0.4777 0 -2.0 1e-06 
0.0 0.4778 0 -2.0 1e-06 
0.0 0.4779 0 -2.0 1e-06 
0.0 0.478 0 -2.0 1e-06 
0.0 0.4781 0 -2.0 1e-06 
0.0 0.4782 0 -2.0 1e-06 
0.0 0.4783 0 -2.0 1e-06 
0.0 0.4784 0 -2.0 1e-06 
0.0 0.4785 0 -2.0 1e-06 
0.0 0.4786 0 -2.0 1e-06 
0.0 0.4787 0 -2.0 1e-06 
0.0 0.4788 0 -2.0 1e-06 
0.0 0.4789 0 -2.0 1e-06 
0.0 0.479 0 -2.0 1e-06 
0.0 0.4791 0 -2.0 1e-06 
0.0 0.4792 0 -2.0 1e-06 
0.0 0.4793 0 -2.0 1e-06 
0.0 0.4794 0 -2.0 1e-06 
0.0 0.4795 0 -2.0 1e-06 
0.0 0.4796 0 -2.0 1e-06 
0.0 0.4797 0 -2.0 1e-06 
0.0 0.4798 0 -2.0 1e-06 
0.0 0.4799 0 -2.0 1e-06 
0.0 0.48 0 -2.0 1e-06 
0.0 0.4801 0 -2.0 1e-06 
0.0 0.4802 0 -2.0 1e-06 
0.0 0.4803 0 -2.0 1e-06 
0.0 0.4804 0 -2.0 1e-06 
0.0 0.4805 0 -2.0 1e-06 
0.0 0.4806 0 -2.0 1e-06 
0.0 0.4807 0 -2.0 1e-06 
0.0 0.4808 0 -2.0 1e-06 
0.0 0.4809 0 -2.0 1e-06 
0.0 0.481 0 -2.0 1e-06 
0.0 0.4811 0 -2.0 1e-06 
0.0 0.4812 0 -2.0 1e-06 
0.0 0.4813 0 -2.0 1e-06 
0.0 0.4814 0 -2.0 1e-06 
0.0 0.4815 0 -2.0 1e-06 
0.0 0.4816 0 -2.0 1e-06 
0.0 0.4817 0 -2.0 1e-06 
0.0 0.4818 0 -2.0 1e-06 
0.0 0.4819 0 -2.0 1e-06 
0.0 0.482 0 -2.0 1e-06 
0.0 0.4821 0 -2.0 1e-06 
0.0 0.4822 0 -2.0 1e-06 
0.0 0.4823 0 -2.0 1e-06 
0.0 0.4824 0 -2.0 1e-06 
0.0 0.4825 0 -2.0 1e-06 
0.0 0.4826 0 -2.0 1e-06 
0.0 0.4827 0 -2.0 1e-06 
0.0 0.4828 0 -2.0 1e-06 
0.0 0.4829 0 -2.0 1e-06 
0.0 0.483 0 -2.0 1e-06 
0.0 0.4831 0 -2.0 1e-06 
0.0 0.4832 0 -2.0 1e-06 
0.0 0.4833 0 -2.0 1e-06 
0.0 0.4834 0 -2.0 1e-06 
0.0 0.4835 0 -2.0 1e-06 
0.0 0.4836 0 -2.0 1e-06 
0.0 0.4837 0 -2.0 1e-06 
0.0 0.4838 0 -2.0 1e-06 
0.0 0.4839 0 -2.0 1e-06 
0.0 0.484 0 -2.0 1e-06 
0.0 0.4841 0 -2.0 1e-06 
0.0 0.4842 0 -2.0 1e-06 
0.0 0.4843 0 -2.0 1e-06 
0.0 0.4844 0 -2.0 1e-06 
0.0 0.4845 0 -2.0 1e-06 
0.0 0.4846 0 -2.0 1e-06 
0.0 0.4847 0 -2.0 1e-06 
0.0 0.4848 0 -2.0 1e-06 
0.0 0.4849 0 -2.0 1e-06 
0.0 0.485 0 -2.0 1e-06 
0.0 0.4851 0 -2.0 1e-06 
0.0 0.4852 0 -2.0 1e-06 
0.0 0.4853 0 -2.0 1e-06 
0.0 0.4854 0 -2.0 1e-06 
0.0 0.4855 0 -2.0 1e-06 
0.0 0.4856 0 -2.0 1e-06 
0.0 0.4857 0 -2.0 1e-06 
0.0 0.4858 0 -2.0 1e-06 
0.0 0.4859 0 -2.0 1e-06 
0.0 0.486 0 -2.0 1e-06 
0.0 0.4861 0 -2.0 1e-06 
0.0 0.4862 0 -2.0 1e-06 
0.0 0.4863 0 -2.0 1e-06 
0.0 0.4864 0 -2.0 1e-06 
0.0 0.4865 0 -2.0 1e-06 
0.0 0.4866 0 -2.0 1e-06 
0.0 0.4867 0 -2.0 1e-06 
0.0 0.4868 0 -2.0 1e-06 
0.0 0.4869 0 -2.0 1e-06 
0.0 0.487 0 -2.0 1e-06 
0.0 0.4871 0 -2.0 1e-06 
0.0 0.4872 0 -2.0 1e-06 
0.0 0.4873 0 -2.0 1e-06 
0.0 0.4874 0 -2.0 1e-06 
0.0 0.4875 0 -2.0 1e-06 
0.0 0.4876 0 -2.0 1e-06 
0.0 0.4877 0 -2.0 1e-06 
0.0 0.4878 0 -2.0 1e-06 
0.0 0.4879 0 -2.0 1e-06 
0.0 0.488 0 -2.0 1e-06 
0.0 0.4881 0 -2.0 1e-06 
0.0 0.4882 0 -2.0 1e-06 
0.0 0.4883 0 -2.0 1e-06 
0.0 0.4884 0 -2.0 1e-06 
0.0 0.4885 0 -2.0 1e-06 
0.0 0.4886 0 -2.0 1e-06 
0.0 0.4887 0 -2.0 1e-06 
0.0 0.4888 0 -2.0 1e-06 
0.0 0.4889 0 -2.0 1e-06 
0.0 0.489 0 -2.0 1e-06 
0.0 0.4891 0 -2.0 1e-06 
0.0 0.4892 0 -2.0 1e-06 
0.0 0.4893 0 -2.0 1e-06 
0.0 0.4894 0 -2.0 1e-06 
0.0 0.4895 0 -2.0 1e-06 
0.0 0.4896 0 -2.0 1e-06 
0.0 0.4897 0 -2.0 1e-06 
0.0 0.4898 0 -2.0 1e-06 
0.0 0.4899 0 -2.0 1e-06 
0.0 0.49 0 -2.0 1e-06 
0.0 0.4901 0 -2.0 1e-06 
0.0 0.4902 0 -2.0 1e-06 
0.0 0.4903 0 -2.0 1e-06 
0.0 0.4904 0 -2.0 1e-06 
0.0 0.4905 0 -2.0 1e-06 
0.0 0.4906 0 -2.0 1e-06 
0.0 0.4907 0 -2.0 1e-06 
0.0 0.4908 0 -2.0 1e-06 
0.0 0.4909 0 -2.0 1e-06 
0.0 0.491 0 -2.0 1e-06 
0.0 0.4911 0 -2.0 1e-06 
0.0 0.4912 0 -2.0 1e-06 
0.0 0.4913 0 -2.0 1e-06 
0.0 0.4914 0 -2.0 1e-06 
0.0 0.4915 0 -2.0 1e-06 
0.0 0.4916 0 -2.0 1e-06 
0.0 0.4917 0 -2.0 1e-06 
0.0 0.4918 0 -2.0 1e-06 
0.0 0.4919 0 -2.0 1e-06 
0.0 0.492 0 -2.0 1e-06 
0.0 0.4921 0 -2.0 1e-06 
0.0 0.4922 0 -2.0 1e-06 
0.0 0.4923 0 -2.0 1e-06 
0.0 0.4924 0 -2.0 1e-06 
0.0 0.4925 0 -2.0 1e-06 
0.0 0.4926 0 -2.0 1e-06 
0.0 0.4927 0 -2.0 1e-06 
0.0 0.4928 0 -2.0 1e-06 
0.0 0.4929 0 -2.0 1e-06 
0.0 0.493 0 -2.0 1e-06 
0.0 0.4931 0 -2.0 1e-06 
0.0 0.4932 0 -2.0 1e-06 
0.0 0.4933 0 -2.0 1e-06 
0.0 0.4934 0 -2.0 1e-06 
0.0 0.4935 0 -2.0 1e-06 
0.0 0.4936 0 -2.0 1e-06 
0.0 0.4937 0 -2.0 1e-06 
0.0 0.4938 0 -2.0 1e-06 
0.0 0.4939 0 -2.0 1e-06 
0.0 0.494 0 -2.0 1e-06 
0.0 0.4941 0 -2.0 1e-06 
0.0 0.4942 0 -2.0 1e-06 
0.0 0.4943 0 -2.0 1e-06 
0.0 0.4944 0 -2.0 1e-06 
0.0 0.4945 0 -2.0 1e-06 
0.0 0.4946 0 -2.0 1e-06 
0.0 0.4947 0 -2.0 1e-06 
0.0 0.4948 0 -2.0 1e-06 
0.0 0.4949 0 -2.0 1e-06 
0.0 0.495 0 -2.0 1e-06 
0.0 0.4951 0 -2.0 1e-06 
0.0 0.4952 0 -2.0 1e-06 
0.0 0.4953 0 -2.0 1e-06 
0.0 0.4954 0 -2.0 1e-06 
0.0 0.4955 0 -2.0 1e-06 
0.0 0.4956 0 -2.0 1e-06 
0.0 0.4957 0 -2.0 1e-06 
0.0 0.4958 0 -2.0 1e-06 
0.0 0.4959 0 -2.0 1e-06 
0.0 0.496 0 -2.0 1e-06 
0.0 0.4961 0 -2.0 1e-06 
0.0 0.4962 0 -2.0 1e-06 
0.0 0.4963 0 -2.0 1e-06 
0.0 0.4964 0 -2.0 1e-06 
0.0 0.4965 0 -2.0 1e-06 
0.0 0.4966 0 -2.0 1e-06 
0.0 0.4967 0 -2.0 1e-06 
0.0 0.4968 0 -2.0 1e-06 
0.0 0.4969 0 -2.0 1e-06 
0.0 0.497 0 -2.0 1e-06 
0.0 0.4971 0 -2.0 1e-06 
0.0 0.4972 0 -2.0 1e-06 
0.0 0.4973 0 -2.0 1e-06 
0.0 0.4974 0 -2.0 1e-06 
0.0 0.4975 0 -2.0 1e-06 
0.0 0.4976 0 -2.0 1e-06 
0.0 0.4977 0 -2.0 1e-06 
0.0 0.4978 0 -2.0 1e-06 
0.0 0.4979 0 -2.0 1e-06 
0.0 0.498 0 -2.0 1e-06 
0.0 0.4981 0 -2.0 1e-06 
0.0 0.4982 0 -2.0 1e-06 
0.0 0.4983 0 -2.0 1e-06 
0.0 0.4984 0 -2.0 1e-06 
0.0 0.4985 0 -2.0 1e-06 
0.0 0.4986 0 -2.0 1e-06 
0.0 0.4987 0 -2.0 1e-06 
0.0 0.4988 0 -2.0 1e-06 
0.0 0.4989 0 -2.0 1e-06 
0.0 0.499 0 -2.0 1e-06 
0.0 0.4991 0 -2.0 1e-06 
0.0 0.4992 0 -2.0 1e-06 
0.0 0.4993 0 -2.0 1e-06 
0.0 0.4994 0 -2.0 1e-06 
0.0 0.4995 0 -2.0 1e-06 
0.0 0.4996 0 -2.0 1e-06 
0.0 0.4997 0 -2.0 1e-06 
0.0 0.4998 0 -2.0 1e-06 
0.0 0.4999 0 -2.0 1e-06 
0.0 0.5 0 -2.0 1e-06 
0.0 0.5001 0 -2.0 1e-06 
0.0 0.5002 0 -2.0 1e-06 
0.0 0.5003 0 -2.0 1e-06 
0.0 0.5004 0 -2.0 1e-06 
0.0 0.5005 0 -2.0 1e-06 
0.0 0.5006 0 -2.0 1e-06 
0.0 0.5007 0 -2.0 1e-06 
0.0 0.5008 0 -2.0 1e-06 
0.0 0.5009 0 -2.0 1e-06 
0.0 0.501 0 -2.0 1e-06 
0.0 0.5011 0 -2.0 1e-06 
0.0 0.5012 0 -2.0 1e-06 
0.0 0.5013 0 -2.0 1e-06 
0.0 0.5014 0 -2.0 1e-06 
0.0 0.5015 0 -2.0 1e-06 
0.0 0.5016 0 -2.0 1e-06 
0.0 0.5017 0 -2.0 1e-06 
0.0 0.5018 0 -2.0 1e-06 
0.0 0.5019 0 -2.0 1e-06 
0.0 0.502 0 -2.0 1e-06 
0.0 0.5021 0 -2.0 1e-06 
0.0 0.5022 0 -2.0 1e-06 
0.0 0.5023 0 -2.0 1e-06 
0.0 0.5024 0 -2.0 1e-06 
0.0 0.5025 0 -2.0 1e-06 
0.0 0.5026 0 -2.0 1e-06 
0.0 0.5027 0 -2.0 1e-06 
0.0 0.5028 0 -2.0 1e-06 
0.0 0.5029 0 -2.0 1e-06 
0.0 0.503 0 -2.0 1e-06 
0.0 0.5031 0 -2.0 1e-06 
0.0 0.5032 0 -2.0 1e-06 
0.0 0.5033 0 -2.0 1e-06 
0.0 0.5034 0 -2.0 1e-06 
0.0 0.5035 0 -2.0 1e-06 
0.0 0.5036 0 -2.0 1e-06 
0.0 0.5037 0 -2.0 1e-06 
0.0 0.5038 0 -2.0 1e-06 
0.0 0.5039 0 -2.0 1e-06 
0.0 0.504 0 -2.0 1e-06 
0.0 0.5041 0 -2.0 1e-06 
0.0 0.5042 0 -2.0 1e-06 
0.0 0.5043 0 -2.0 1e-06 
0.0 0.5044 0 -2.0 1e-06 
0.0 0.5045 0 -2.0 1e-06 
0.0 0.5046 0 -2.0 1e-06 
0.0 0.5047 0 -2.0 1e-06 
0.0 0.5048 0 -2.0 1e-06 
0.0 0.5049 0 -2.0 1e-06 
0.0 0.505 0 -2.0 1e-06 
0.0 0.5051 0 -2.0 1e-06 
0.0 0.5052 0 -2.0 1e-06 
0.0 0.5053 0 -2.0 1e-06 
0.0 0.5054 0 -2.0 1e-06 
0.0 0.5055 0 -2.0 1e-06 
0.0 0.5056 0 -2.0 1e-06 
0.0 0.5057 0 -2.0 1e-06 
0.0 0.5058 0 -2.0 1e-06 
0.0 0.5059 0 -2.0 1e-06 
0.0 0.506 0 -2.0 1e-06 
0.0 0.5061 0 -2.0 1e-06 
0.0 0.5062 0 -2.0 1e-06 
0.0 0.5063 0 -2.0 1e-06 
0.0 0.5064 0 -2.0 1e-06 
0.0 0.5065 0 -2.0 1e-06 
0.0 0.5066 0 -2.0 1e-06 
0.0 0.5067 0 -2.0 1e-06 
0.0 0.5068 0 -2.0 1e-06 
0.0 0.5069 0 -2.0 1e-06 
0.0 0.507 0 -2.0 1e-06 
0.0 0.5071 0 -2.0 1e-06 
0.0 0.5072 0 -2.0 1e-06 
0.0 0.5073 0 -2.0 1e-06 
0.0 0.5074 0 -2.0 1e-06 
0.0 0.5075 0 -2.0 1e-06 
0.0 0.5076 0 -2.0 1e-06 
0.0 0.5077 0 -2.0 1e-06 
0.0 0.5078 0 -2.0 1e-06 
0.0 0.5079 0 -2.0 1e-06 
0.0 0.508 0 -2.0 1e-06 
0.0 0.5081 0 -2.0 1e-06 
0.0 0.5082 0 -2.0 1e-06 
0.0 0.5083 0 -2.0 1e-06 
0.0 0.5084 0 -2.0 1e-06 
0.0 0.5085 0 -2.0 1e-06 
0.0 0.5086 0 -2.0 1e-06 
0.0 0.5087 0 -2.0 1e-06 
0.0 0.5088 0 -2.0 1e-06 
0.0 0.5089 0 -2.0 1e-06 
0.0 0.509 0 -2.0 1e-06 
0.0 0.5091 0 -2.0 1e-06 
0.0 0.5092 0 -2.0 1e-06 
0.0 0.5093 0 -2.0 1e-06 
0.0 0.5094 0 -2.0 1e-06 
0.0 0.5095 0 -2.0 1e-06 
0.0 0.5096 0 -2.0 1e-06 
0.0 0.5097 0 -2.0 1e-06 
0.0 0.5098 0 -2.0 1e-06 
0.0 0.5099 0 -2.0 1e-06 
0.0 0.51 0 -2.0 1e-06 
0.0 0.5101 0 -2.0 1e-06 
0.0 0.5102 0 -2.0 1e-06 
0.0 0.5103 0 -2.0 1e-06 
0.0 0.5104 0 -2.0 1e-06 
0.0 0.5105 0 -2.0 1e-06 
0.0 0.5106 0 -2.0 1e-06 
0.0 0.5107 0 -2.0 1e-06 
0.0 0.5108 0 -2.0 1e-06 
0.0 0.5109 0 -2.0 1e-06 
0.0 0.511 0 -2.0 1e-06 
0.0 0.5111 0 -2.0 1e-06 
0.0 0.5112 0 -2.0 1e-06 
0.0 0.5113 0 -2.0 1e-06 
0.0 0.5114 0 -2.0 1e-06 
0.0 0.5115 0 -2.0 1e-06 
0.0 0.5116 0 -2.0 1e-06 
0.0 0.5117 0 -2.0 1e-06 
0.0 0.5118 0 -2.0 1e-06 
0.0 0.5119 0 -2.0 1e-06 
0.0 0.512 0 -2.0 1e-06 
0.0 0.5121 0 -2.0 1e-06 
0.0 0.5122 0 -2.0 1e-06 
0.0 0.5123 0 -2.0 1e-06 
0.0 0.5124 0 -2.0 1e-06 
0.0 0.5125 0 -2.0 1e-06 
0.0 0.5126 0 -2.0 1e-06 
0.0 0.5127 0 -2.0 1e-06 
0.0 0.5128 0 -2.0 1e-06 
0.0 0.5129 0 -2.0 1e-06 
0.0 0.513 0 -2.0 1e-06 
0.0 0.5131 0 -2.0 1e-06 
0.0 0.5132 0 -2.0 1e-06 
0.0 0.5133 0 -2.0 1e-06 
0.0 0.5134 0 -2.0 1e-06 
0.0 0.5135 0 -2.0 1e-06 
0.0 0.5136 0 -2.0 1e-06 
0.0 0.5137 0 -2.0 1e-06 
0.0 0.5138 0 -2.0 1e-06 
0.0 0.5139 0 -2.0 1e-06 
0.0 0.514 0 -2.0 1e-06 
0.0 0.5141 0 -2.0 1e-06 
0.0 0.5142 0 -2.0 1e-06 
0.0 0.5143 0 -2.0 1e-06 
0.0 0.5144 0 -2.0 1e-06 
0.0 0.5145 0 -2.0 1e-06 
0.0 0.5146 0 -2.0 1e-06 
0.0 0.5147 0 -2.0 1e-06 
0.0 0.5148 0 -2.0 1e-06 
0.0 0.5149 0 -2.0 1e-06 
0.0 0.515 0 -2.0 1e-06 
0.0 0.5151 0 -2.0 1e-06 
0.0 0.5152 0 -2.0 1e-06 
0.0 0.5153 0 -2.0 1e-06 
0.0 0.5154 0 -2.0 1e-06 
0.0 0.5155 0 -2.0 1e-06 
0.0 0.5156 0 -2.0 1e-06 
0.0 0.5157 0 -2.0 1e-06 
0.0 0.5158 0 -2.0 1e-06 
0.0 0.5159 0 -2.0 1e-06 
0.0 0.516 0 -2.0 1e-06 
0.0 0.5161 0 -2.0 1e-06 
0.0 0.5162 0 -2.0 1e-06 
0.0 0.5163 0 -2.0 1e-06 
0.0 0.5164 0 -2.0 1e-06 
0.0 0.5165 0 -2.0 1e-06 
0.0 0.5166 0 -2.0 1e-06 
0.0 0.5167 0 -2.0 1e-06 
0.0 0.5168 0 -2.0 1e-06 
0.0 0.5169 0 -2.0 1e-06 
0.0 0.517 0 -2.0 1e-06 
0.0 0.5171 0 -2.0 1e-06 
0.0 0.5172 0 -2.0 1e-06 
0.0 0.5173 0 -2.0 1e-06 
0.0 0.5174 0 -2.0 1e-06 
0.0 0.5175 0 -2.0 1e-06 
0.0 0.5176 0 -2.0 1e-06 
0.0 0.5177 0 -2.0 1e-06 
0.0 0.5178 0 -2.0 1e-06 
0.0 0.5179 0 -2.0 1e-06 
0.0 0.518 0 -2.0 1e-06 
0.0 0.5181 0 -2.0 1e-06 
0.0 0.5182 0 -2.0 1e-06 
0.0 0.5183 0 -2.0 1e-06 
0.0 0.5184 0 -2.0 1e-06 
0.0 0.5185 0 -2.0 1e-06 
0.0 0.5186 0 -2.0 1e-06 
0.0 0.5187 0 -2.0 1e-06 
0.0 0.5188 0 -2.0 1e-06 
0.0 0.5189 0 -2.0 1e-06 
0.0 0.519 0 -2.0 1e-06 
0.0 0.5191 0 -2.0 1e-06 
0.0 0.5192 0 -2.0 1e-06 
0.0 0.5193 0 -2.0 1e-06 
0.0 0.5194 0 -2.0 1e-06 
0.0 0.5195 0 -2.0 1e-06 
0.0 0.5196 0 -2.0 1e-06 
0.0 0.5197 0 -2.0 1e-06 
0.0 0.5198 0 -2.0 1e-06 
0.0 0.5199 0 -2.0 1e-06 
0.0 0.52 0 -2.0 1e-06 
0.0 0.5201 0 -2.0 1e-06 
0.0 0.5202 0 -2.0 1e-06 
0.0 0.5203 0 -2.0 1e-06 
0.0 0.5204 0 -2.0 1e-06 
0.0 0.5205 0 -2.0 1e-06 
0.0 0.5206 0 -2.0 1e-06 
0.0 0.5207 0 -2.0 1e-06 
0.0 0.5208 0 -2.0 1e-06 
0.0 0.5209 0 -2.0 1e-06 
0.0 0.521 0 -2.0 1e-06 
0.0 0.5211 0 -2.0 1e-06 
0.0 0.5212 0 -2.0 1e-06 
0.0 0.5213 0 -2.0 1e-06 
0.0 0.5214 0 -2.0 1e-06 
0.0 0.5215 0 -2.0 1e-06 
0.0 0.5216 0 -2.0 1e-06 
0.0 0.5217 0 -2.0 1e-06 
0.0 0.5218 0 -2.0 1e-06 
0.0 0.5219 0 -2.0 1e-06 
0.0 0.522 0 -2.0 1e-06 
0.0 0.5221 0 -2.0 1e-06 
0.0 0.5222 0 -2.0 1e-06 
0.0 0.5223 0 -2.0 1e-06 
0.0 0.5224 0 -2.0 1e-06 
0.0 0.5225 0 -2.0 1e-06 
0.0 0.5226 0 -2.0 1e-06 
0.0 0.5227 0 -2.0 1e-06 
0.0 0.5228 0 -2.0 1e-06 
0.0 0.5229 0 -2.0 1e-06 
0.0 0.523 0 -2.0 1e-06 
0.0 0.5231 0 -2.0 1e-06 
0.0 0.5232 0 -2.0 1e-06 
0.0 0.5233 0 -2.0 1e-06 
0.0 0.5234 0 -2.0 1e-06 
0.0 0.5235 0 -2.0 1e-06 
0.0 0.5236 0 -2.0 1e-06 
0.0 0.5237 0 -2.0 1e-06 
0.0 0.5238 0 -2.0 1e-06 
0.0 0.5239 0 -2.0 1e-06 
0.0 0.524 0 -2.0 1e-06 
0.0 0.5241 0 -2.0 1e-06 
0.0 0.5242 0 -2.0 1e-06 
0.0 0.5243 0 -2.0 1e-06 
0.0 0.5244 0 -2.0 1e-06 
0.0 0.5245 0 -2.0 1e-06 
0.0 0.5246 0 -2.0 1e-06 
0.0 0.5247 0 -2.0 1e-06 
0.0 0.5248 0 -2.0 1e-06 
0.0 0.5249 0 -2.0 1e-06 
0.0 0.525 0 -2.0 1e-06 
0.0 0.5251 0 -2.0 1e-06 
0.0 0.5252 0 -2.0 1e-06 
0.0 0.5253 0 -2.0 1e-06 
0.0 0.5254 0 -2.0 1e-06 
0.0 0.5255 0 -2.0 1e-06 
0.0 0.5256 0 -2.0 1e-06 
0.0 0.5257 0 -2.0 1e-06 
0.0 0.5258 0 -2.0 1e-06 
0.0 0.5259 0 -2.0 1e-06 
0.0 0.526 0 -2.0 1e-06 
0.0 0.5261 0 -2.0 1e-06 
0.0 0.5262 0 -2.0 1e-06 
0.0 0.5263 0 -2.0 1e-06 
0.0 0.5264 0 -2.0 1e-06 
0.0 0.5265 0 -2.0 1e-06 
0.0 0.5266 0 -2.0 1e-06 
0.0 0.5267 0 -2.0 1e-06 
0.0 0.5268 0 -2.0 1e-06 
0.0 0.5269 0 -2.0 1e-06 
0.0 0.527 0 -2.0 1e-06 
0.0 0.5271 0 -2.0 1e-06 
0.0 0.5272 0 -2.0 1e-06 
0.0 0.5273 0 -2.0 1e-06 
0.0 0.5274 0 -2.0 1e-06 
0.0 0.5275 0 -2.0 1e-06 
0.0 0.5276 0 -2.0 1e-06 
0.0 0.5277 0 -2.0 1e-06 
0.0 0.5278 0 -2.0 1e-06 
0.0 0.5279 0 -2.0 1e-06 
0.0 0.528 0 -2.0 1e-06 
0.0 0.5281 0 -2.0 1e-06 
0.0 0.5282 0 -2.0 1e-06 
0.0 0.5283 0 -2.0 1e-06 
0.0 0.5284 0 -2.0 1e-06 
0.0 0.5285 0 -2.0 1e-06 
0.0 0.5286 0 -2.0 1e-06 
0.0 0.5287 0 -2.0 1e-06 
0.0 0.5288 0 -2.0 1e-06 
0.0 0.5289 0 -2.0 1e-06 
0.0 0.529 0 -2.0 1e-06 
0.0 0.5291 0 -2.0 1e-06 
0.0 0.5292 0 -2.0 1e-06 
0.0 0.5293 0 -2.0 1e-06 
0.0 0.5294 0 -2.0 1e-06 
0.0 0.5295 0 -2.0 1e-06 
0.0 0.5296 0 -2.0 1e-06 
0.0 0.5297 0 -2.0 1e-06 
0.0 0.5298 0 -2.0 1e-06 
0.0 0.5299 0 -2.0 1e-06 
0.0 0.53 0 -2.0 1e-06 
0.0 0.5301 0 -2.0 1e-06 
0.0 0.5302 0 -2.0 1e-06 
0.0 0.5303 0 -2.0 1e-06 
0.0 0.5304 0 -2.0 1e-06 
0.0 0.5305 0 -2.0 1e-06 
0.0 0.5306 0 -2.0 1e-06 
0.0 0.5307 0 -2.0 1e-06 
0.0 0.5308 0 -2.0 1e-06 
0.0 0.5309 0 -2.0 1e-06 
0.0 0.531 0 -2.0 1e-06 
0.0 0.5311 0 -2.0 1e-06 
0.0 0.5312 0 -2.0 1e-06 
0.0 0.5313 0 -2.0 1e-06 
0.0 0.5314 0 -2.0 1e-06 
0.0 0.5315 0 -2.0 1e-06 
0.0 0.5316 0 -2.0 1e-06 
0.0 0.5317 0 -2.0 1e-06 
0.0 0.5318 0 -2.0 1e-06 
0.0 0.5319 0 -2.0 1e-06 
0.0 0.532 0 -2.0 1e-06 
0.0 0.5321 0 -2.0 1e-06 
0.0 0.5322 0 -2.0 1e-06 
0.0 0.5323 0 -2.0 1e-06 
0.0 0.5324 0 -2.0 1e-06 
0.0 0.5325 0 -2.0 1e-06 
0.0 0.5326 0 -2.0 1e-06 
0.0 0.5327 0 -2.0 1e-06 
0.0 0.5328 0 -2.0 1e-06 
0.0 0.5329 0 -2.0 1e-06 
0.0 0.533 0 -2.0 1e-06 
0.0 0.5331 0 -2.0 1e-06 
0.0 0.5332 0 -2.0 1e-06 
0.0 0.5333 0 -2.0 1e-06 
0.0 0.5334 0 -2.0 1e-06 
0.0 0.5335 0 -2.0 1e-06 
0.0 0.5336 0 -2.0 1e-06 
0.0 0.5337 0 -2.0 1e-06 
0.0 0.5338 0 -2.0 1e-06 
0.0 0.5339 0 -2.0 1e-06 
0.0 0.534 0 -2.0 1e-06 
0.0 0.5341 0 -2.0 1e-06 
0.0 0.5342 0 -2.0 1e-06 
0.0 0.5343 0 -2.0 1e-06 
0.0 0.5344 0 -2.0 1e-06 
0.0 0.5345 0 -2.0 1e-06 
0.0 0.5346 0 -2.0 1e-06 
0.0 0.5347 0 -2.0 1e-06 
0.0 0.5348 0 -2.0 1e-06 
0.0 0.5349 0 -2.0 1e-06 
0.0 0.535 0 -2.0 1e-06 
0.0 0.5351 0 -2.0 1e-06 
0.0 0.5352 0 -2.0 1e-06 
0.0 0.5353 0 -2.0 1e-06 
0.0 0.5354 0 -2.0 1e-06 
0.0 0.5355 0 -2.0 1e-06 
0.0 0.5356 0 -2.0 1e-06 
0.0 0.5357 0 -2.0 1e-06 
0.0 0.5358 0 -2.0 1e-06 
0.0 0.5359 0 -2.0 1e-06 
0.0 0.536 0 -2.0 1e-06 
0.0 0.5361 0 -2.0 1e-06 
0.0 0.5362 0 -2.0 1e-06 
0.0 0.5363 0 -2.0 1e-06 
0.0 0.5364 0 -2.0 1e-06 
0.0 0.5365 0 -2.0 1e-06 
0.0 0.5366 0 -2.0 1e-06 
0.0 0.5367 0 -2.0 1e-06 
0.0 0.5368 0 -2.0 1e-06 
0.0 0.5369 0 -2.0 1e-06 
0.0 0.537 0 -2.0 1e-06 
0.0 0.5371 0 -2.0 1e-06 
0.0 0.5372 0 -2.0 1e-06 
0.0 0.5373 0 -2.0 1e-06 
0.0 0.5374 0 -2.0 1e-06 
0.0 0.5375 0 -2.0 1e-06 
0.0 0.5376 0 -2.0 1e-06 
0.0 0.5377 0 -2.0 1e-06 
0.0 0.5378 0 -2.0 1e-06 
0.0 0.5379 0 -2.0 1e-06 
0.0 0.538 0 -2.0 1e-06 
0.0 0.5381 0 -2.0 1e-06 
0.0 0.5382 0 -2.0 1e-06 
0.0 0.5383 0 -2.0 1e-06 
0.0 0.5384 0 -2.0 1e-06 
0.0 0.5385 0 -2.0 1e-06 
0.0 0.5386 0 -2.0 1e-06 
0.0 0.5387 0 -2.0 1e-06 
0.0 0.5388 0 -2.0 1e-06 
0.0 0.5389 0 -2.0 1e-06 
0.0 0.539 0 -2.0 1e-06 
0.0 0.5391 0 -2.0 1e-06 
0.0 0.5392 0 -2.0 1e-06 
0.0 0.5393 0 -2.0 1e-06 
0.0 0.5394 0 -2.0 1e-06 
0.0 0.5395 0 -2.0 1e-06 
0.0 0.5396 0 -2.0 1e-06 
0.0 0.5397 0 -2.0 1e-06 
0.0 0.5398 0 -2.0 1e-06 
0.0 0.5399 0 -2.0 1e-06 
0.0 0.54 0 -2.0 1e-06 
0.0 0.5401 0 -2.0 1e-06 
0.0 0.5402 0 -2.0 1e-06 
0.0 0.5403 0 -2.0 1e-06 
0.0 0.5404 0 -2.0 1e-06 
0.0 0.5405 0 -2.0 1e-06 
0.0 0.5406 0 -2.0 1e-06 
0.0 0.5407 0 -2.0 1e-06 
0.0 0.5408 0 -2.0 1e-06 
0.0 0.5409 0 -2.0 1e-06 
0.0 0.541 0 -2.0 1e-06 
0.0 0.5411 0 -2.0 1e-06 
0.0 0.5412 0 -2.0 1e-06 
0.0 0.5413 0 -2.0 1e-06 
0.0 0.5414 0 -2.0 1e-06 
0.0 0.5415 0 -2.0 1e-06 
0.0 0.5416 0 -2.0 1e-06 
0.0 0.5417 0 -2.0 1e-06 
0.0 0.5418 0 -2.0 1e-06 
0.0 0.5419 0 -2.0 1e-06 
0.0 0.542 0 -2.0 1e-06 
0.0 0.5421 0 -2.0 1e-06 
0.0 0.5422 0 -2.0 1e-06 
0.0 0.5423 0 -2.0 1e-06 
0.0 0.5424 0 -2.0 1e-06 
0.0 0.5425 0 -2.0 1e-06 
0.0 0.5426 0 -2.0 1e-06 
0.0 0.5427 0 -2.0 1e-06 
0.0 0.5428 0 -2.0 1e-06 
0.0 0.5429 0 -2.0 1e-06 
0.0 0.543 0 -2.0 1e-06 
0.0 0.5431 0 -2.0 1e-06 
0.0 0.5432 0 -2.0 1e-06 
0.0 0.5433 0 -2.0 1e-06 
0.0 0.5434 0 -2.0 1e-06 
0.0 0.5435 0 -2.0 1e-06 
0.0 0.5436 0 -2.0 1e-06 
0.0 0.5437 0 -2.0 1e-06 
0.0 0.5438 0 -2.0 1e-06 
0.0 0.5439 0 -2.0 1e-06 
0.0 0.544 0 -2.0 1e-06 
0.0 0.5441 0 -2.0 1e-06 
0.0 0.5442 0 -2.0 1e-06 
0.0 0.5443 0 -2.0 1e-06 
0.0 0.5444 0 -2.0 1e-06 
0.0 0.5445 0 -2.0 1e-06 
0.0 0.5446 0 -2.0 1e-06 
0.0 0.5447 0 -2.0 1e-06 
0.0 0.5448 0 -2.0 1e-06 
0.0 0.5449 0 -2.0 1e-06 
0.0 0.545 0 -2.0 1e-06 
0.0 0.5451 0 -2.0 1e-06 
0.0 0.5452 0 -2.0 1e-06 
0.0 0.5453 0 -2.0 1e-06 
0.0 0.5454 0 -2.0 1e-06 
0.0 0.5455 0 -2.0 1e-06 
0.0 0.5456 0 -2.0 1e-06 
0.0 0.5457 0 -2.0 1e-06 
0.0 0.5458 0 -2.0 1e-06 
0.0 0.5459 0 -2.0 1e-06 
0.0 0.546 0 -2.0 1e-06 
0.0 0.5461 0 -2.0 1e-06 
0.0 0.5462 0 -2.0 1e-06 
0.0 0.5463 0 -2.0 1e-06 
0.0 0.5464 0 -2.0 1e-06 
0.0 0.5465 0 -2.0 1e-06 
0.0 0.5466 0 -2.0 1e-06 
0.0 0.5467 0 -2.0 1e-06 
0.0 0.5468 0 -2.0 1e-06 
0.0 0.5469 0 -2.0 1e-06 
0.0 0.547 0 -2.0 1e-06 
0.0 0.5471 0 -2.0 1e-06 
0.0 0.5472 0 -2.0 1e-06 
0.0 0.5473 0 -2.0 1e-06 
0.0 0.5474 0 -2.0 1e-06 
0.0 0.5475 0 -2.0 1e-06 
0.0 0.5476 0 -2.0 1e-06 
0.0 0.5477 0 -2.0 1e-06 
0.0 0.5478 0 -2.0 1e-06 
0.0 0.5479 0 -2.0 1e-06 
0.0 0.548 0 -2.0 1e-06 
0.0 0.5481 0 -2.0 1e-06 
0.0 0.5482 0 -2.0 1e-06 
0.0 0.5483 0 -2.0 1e-06 
0.0 0.5484 0 -2.0 1e-06 
0.0 0.5485 0 -2.0 1e-06 
0.0 0.5486 0 -2.0 1e-06 
0.0 0.5487 0 -2.0 1e-06 
0.0 0.5488 0 -2.0 1e-06 
0.0 0.5489 0 -2.0 1e-06 
0.0 0.549 0 -2.0 1e-06 
0.0 0.5491 0 -2.0 1e-06 
0.0 0.5492 0 -2.0 1e-06 
0.0 0.5493 0 -2.0 1e-06 
0.0 0.5494 0 -2.0 1e-06 
0.0 0.5495 0 -2.0 1e-06 
0.0 0.5496 0 -2.0 1e-06 
0.0 0.5497 0 -2.0 1e-06 
0.0 0.5498 0 -2.0 1e-06 
0.0 0.5499 0 -2.0 1e-06 
0.0 0.55 0 -2.0 1e-06 
0.0 0.5501 0 -2.0 1e-06 
0.0 0.5502 0 -2.0 1e-06 
0.0 0.5503 0 -2.0 1e-06 
0.0 0.5504 0 -2.0 1e-06 
0.0 0.5505 0 -2.0 1e-06 
0.0 0.5506 0 -2.0 1e-06 
0.0 0.5507 0 -2.0 1e-06 
0.0 0.5508 0 -2.0 1e-06 
0.0 0.5509 0 -2.0 1e-06 
0.0 0.551 0 -2.0 1e-06 
0.0 0.5511 0 -2.0 1e-06 
0.0 0.5512 0 -2.0 1e-06 
0.0 0.5513 0 -2.0 1e-06 
0.0 0.5514 0 -2.0 1e-06 
0.0 0.5515 0 -2.0 1e-06 
0.0 0.5516 0 -2.0 1e-06 
0.0 0.5517 0 -2.0 1e-06 
0.0 0.5518 0 -2.0 1e-06 
0.0 0.5519 0 -2.0 1e-06 
0.0 0.552 0 -2.0 1e-06 
0.0 0.5521 0 -2.0 1e-06 
0.0 0.5522 0 -2.0 1e-06 
0.0 0.5523 0 -2.0 1e-06 
0.0 0.5524 0 -2.0 1e-06 
0.0 0.5525 0 -2.0 1e-06 
0.0 0.5526 0 -2.0 1e-06 
0.0 0.5527 0 -2.0 1e-06 
0.0 0.5528 0 -2.0 1e-06 
0.0 0.5529 0 -2.0 1e-06 
0.0 0.553 0 -2.0 1e-06 
0.0 0.5531 0 -2.0 1e-06 
0.0 0.5532 0 -2.0 1e-06 
0.0 0.5533 0 -2.0 1e-06 
0.0 0.5534 0 -2.0 1e-06 
0.0 0.5535 0 -2.0 1e-06 
0.0 0.5536 0 -2.0 1e-06 
0.0 0.5537 0 -2.0 1e-06 
0.0 0.5538 0 -2.0 1e-06 
0.0 0.5539 0 -2.0 1e-06 
0.0 0.554 0 -2.0 1e-06 
0.0 0.5541 0 -2.0 1e-06 
0.0 0.5542 0 -2.0 1e-06 
0.0 0.5543 0 -2.0 1e-06 
0.0 0.5544 0 -2.0 1e-06 
0.0 0.5545 0 -2.0 1e-06 
0.0 0.5546 0 -2.0 1e-06 
0.0 0.5547 0 -2.0 1e-06 
0.0 0.5548 0 -2.0 1e-06 
0.0 0.5549 0 -2.0 1e-06 
0.0 0.555 0 -2.0 1e-06 
0.0 0.5551 0 -2.0 1e-06 
0.0 0.5552 0 -2.0 1e-06 
0.0 0.5553 0 -2.0 1e-06 
0.0 0.5554 0 -2.0 1e-06 
0.0 0.5555 0 -2.0 1e-06 
0.0 0.5556 0 -2.0 1e-06 
0.0 0.5557 0 -2.0 1e-06 
0.0 0.5558 0 -2.0 1e-06 
0.0 0.5559 0 -2.0 1e-06 
0.0 0.556 0 -2.0 1e-06 
0.0 0.5561 0 -2.0 1e-06 
0.0 0.5562 0 -2.0 1e-06 
0.0 0.5563 0 -2.0 1e-06 
0.0 0.5564 0 -2.0 1e-06 
0.0 0.5565 0 -2.0 1e-06 
0.0 0.5566 0 -2.0 1e-06 
0.0 0.5567 0 -2.0 1e-06 
0.0 0.5568 0 -2.0 1e-06 
0.0 0.5569 0 -2.0 1e-06 
0.0 0.557 0 -2.0 1e-06 
0.0 0.5571 0 -2.0 1e-06 
0.0 0.5572 0 -2.0 1e-06 
0.0 0.5573 0 -2.0 1e-06 
0.0 0.5574 0 -2.0 1e-06 
0.0 0.5575 0 -2.0 1e-06 
0.0 0.5576 0 -2.0 1e-06 
0.0 0.5577 0 -2.0 1e-06 
0.0 0.5578 0 -2.0 1e-06 
0.0 0.5579 0 -2.0 1e-06 
0.0 0.558 0 -2.0 1e-06 
0.0 0.5581 0 -2.0 1e-06 
0.0 0.5582 0 -2.0 1e-06 
0.0 0.5583 0 -2.0 1e-06 
0.0 0.5584 0 -2.0 1e-06 
0.0 0.5585 0 -2.0 1e-06 
0.0 0.5586 0 -2.0 1e-06 
0.0 0.5587 0 -2.0 1e-06 
0.0 0.5588 0 -2.0 1e-06 
0.0 0.5589 0 -2.0 1e-06 
0.0 0.559 0 -2.0 1e-06 
0.0 0.5591 0 -2.0 1e-06 
0.0 0.5592 0 -2.0 1e-06 
0.0 0.5593 0 -2.0 1e-06 
0.0 0.5594 0 -2.0 1e-06 
0.0 0.5595 0 -2.0 1e-06 
0.0 0.5596 0 -2.0 1e-06 
0.0 0.5597 0 -2.0 1e-06 
0.0 0.5598 0 -2.0 1e-06 
0.0 0.5599 0 -2.0 1e-06 
0.0 0.56 0 -2.0 1e-06 
0.0 0.5601 0 -2.0 1e-06 
0.0 0.5602 0 -2.0 1e-06 
0.0 0.5603 0 -2.0 1e-06 
0.0 0.5604 0 -2.0 1e-06 
0.0 0.5605 0 -2.0 1e-06 
0.0 0.5606 0 -2.0 1e-06 
0.0 0.5607 0 -2.0 1e-06 
0.0 0.5608 0 -2.0 1e-06 
0.0 0.5609 0 -2.0 1e-06 
0.0 0.561 0 -2.0 1e-06 
0.0 0.5611 0 -2.0 1e-06 
0.0 0.5612 0 -2.0 1e-06 
0.0 0.5613 0 -2.0 1e-06 
0.0 0.5614 0 -2.0 1e-06 
0.0 0.5615 0 -2.0 1e-06 
0.0 0.5616 0 -2.0 1e-06 
0.0 0.5617 0 -2.0 1e-06 
0.0 0.5618 0 -2.0 1e-06 
0.0 0.5619 0 -2.0 1e-06 
0.0 0.562 0 -2.0 1e-06 
0.0 0.5621 0 -2.0 1e-06 
0.0 0.5622 0 -2.0 1e-06 
0.0 0.5623 0 -2.0 1e-06 
0.0 0.5624 0 -2.0 1e-06 
0.0 0.5625 0 -2.0 1e-06 
0.0 0.5626 0 -2.0 1e-06 
0.0 0.5627 0 -2.0 1e-06 
0.0 0.5628 0 -2.0 1e-06 
0.0 0.5629 0 -2.0 1e-06 
0.0 0.563 0 -2.0 1e-06 
0.0 0.5631 0 -2.0 1e-06 
0.0 0.5632 0 -2.0 1e-06 
0.0 0.5633 0 -2.0 1e-06 
0.0 0.5634 0 -2.0 1e-06 
0.0 0.5635 0 -2.0 1e-06 
0.0 0.5636 0 -2.0 1e-06 
0.0 0.5637 0 -2.0 1e-06 
0.0 0.5638 0 -2.0 1e-06 
0.0 0.5639 0 -2.0 1e-06 
0.0 0.564 0 -2.0 1e-06 
0.0 0.5641 0 -2.0 1e-06 
0.0 0.5642 0 -2.0 1e-06 
0.0 0.5643 0 -2.0 1e-06 
0.0 0.5644 0 -2.0 1e-06 
0.0 0.5645 0 -2.0 1e-06 
0.0 0.5646 0 -2.0 1e-06 
0.0 0.5647 0 -2.0 1e-06 
0.0 0.5648 0 -2.0 1e-06 
0.0 0.5649 0 -2.0 1e-06 
0.0 0.565 0 -2.0 1e-06 
0.0 0.5651 0 -2.0 1e-06 
0.0 0.5652 0 -2.0 1e-06 
0.0 0.5653 0 -2.0 1e-06 
0.0 0.5654 0 -2.0 1e-06 
0.0 0.5655 0 -2.0 1e-06 
0.0 0.5656 0 -2.0 1e-06 
0.0 0.5657 0 -2.0 1e-06 
0.0 0.5658 0 -2.0 1e-06 
0.0 0.5659 0 -2.0 1e-06 
0.0 0.566 0 -2.0 1e-06 
0.0 0.5661 0 -2.0 1e-06 
0.0 0.5662 0 -2.0 1e-06 
0.0 0.5663 0 -2.0 1e-06 
0.0 0.5664 0 -2.0 1e-06 
0.0 0.5665 0 -2.0 1e-06 
0.0 0.5666 0 -2.0 1e-06 
0.0 0.5667 0 -2.0 1e-06 
0.0 0.5668 0 -2.0 1e-06 
0.0 0.5669 0 -2.0 1e-06 
0.0 0.567 0 -2.0 1e-06 
0.0 0.5671 0 -2.0 1e-06 
0.0 0.5672 0 -2.0 1e-06 
0.0 0.5673 0 -2.0 1e-06 
0.0 0.5674 0 -2.0 1e-06 
0.0 0.5675 0 -2.0 1e-06 
0.0 0.5676 0 -2.0 1e-06 
0.0 0.5677 0 -2.0 1e-06 
0.0 0.5678 0 -2.0 1e-06 
0.0 0.5679 0 -2.0 1e-06 
0.0 0.568 0 -2.0 1e-06 
0.0 0.5681 0 -2.0 1e-06 
0.0 0.5682 0 -2.0 1e-06 
0.0 0.5683 0 -2.0 1e-06 
0.0 0.5684 0 -2.0 1e-06 
0.0 0.5685 0 -2.0 1e-06 
0.0 0.5686 0 -2.0 1e-06 
0.0 0.5687 0 -2.0 1e-06 
0.0 0.5688 0 -2.0 1e-06 
0.0 0.5689 0 -2.0 1e-06 
0.0 0.569 0 -2.0 1e-06 
0.0 0.5691 0 -2.0 1e-06 
0.0 0.5692 0 -2.0 1e-06 
0.0 0.5693 0 -2.0 1e-06 
0.0 0.5694 0 -2.0 1e-06 
0.0 0.5695 0 -2.0 1e-06 
0.0 0.5696 0 -2.0 1e-06 
0.0 0.5697 0 -2.0 1e-06 
0.0 0.5698 0 -2.0 1e-06 
0.0 0.5699 0 -2.0 1e-06 
0.0 0.57 0 -2.0 1e-06 
0.0 0.5701 0 -2.0 1e-06 
0.0 0.5702 0 -2.0 1e-06 
0.0 0.5703 0 -2.0 1e-06 
0.0 0.5704 0 -2.0 1e-06 
0.0 0.5705 0 -2.0 1e-06 
0.0 0.5706 0 -2.0 1e-06 
0.0 0.5707 0 -2.0 1e-06 
0.0 0.5708 0 -2.0 1e-06 
0.0 0.5709 0 -2.0 1e-06 
0.0 0.571 0 -2.0 1e-06 
0.0 0.5711 0 -2.0 1e-06 
0.0 0.5712 0 -2.0 1e-06 
0.0 0.5713 0 -2.0 1e-06 
0.0 0.5714 0 -2.0 1e-06 
0.0 0.5715 0 -2.0 1e-06 
0.0 0.5716 0 -2.0 1e-06 
0.0 0.5717 0 -2.0 1e-06 
0.0 0.5718 0 -2.0 1e-06 
0.0 0.5719 0 -2.0 1e-06 
0.0 0.572 0 -2.0 1e-06 
0.0 0.5721 0 -2.0 1e-06 
0.0 0.5722 0 -2.0 1e-06 
0.0 0.5723 0 -2.0 1e-06 
0.0 0.5724 0 -2.0 1e-06 
0.0 0.5725 0 -2.0 1e-06 
0.0 0.5726 0 -2.0 1e-06 
0.0 0.5727 0 -2.0 1e-06 
0.0 0.5728 0 -2.0 1e-06 
0.0 0.5729 0 -2.0 1e-06 
0.0 0.573 0 -2.0 1e-06 
0.0 0.5731 0 -2.0 1e-06 
0.0 0.5732 0 -2.0 1e-06 
0.0 0.5733 0 -2.0 1e-06 
0.0 0.5734 0 -2.0 1e-06 
0.0 0.5735 0 -2.0 1e-06 
0.0 0.5736 0 -2.0 1e-06 
0.0 0.5737 0 -2.0 1e-06 
0.0 0.5738 0 -2.0 1e-06 
0.0 0.5739 0 -2.0 1e-06 
0.0 0.574 0 -2.0 1e-06 
0.0 0.5741 0 -2.0 1e-06 
0.0 0.5742 0 -2.0 1e-06 
0.0 0.5743 0 -2.0 1e-06 
0.0 0.5744 0 -2.0 1e-06 
0.0 0.5745 0 -2.0 1e-06 
0.0 0.5746 0 -2.0 1e-06 
0.0 0.5747 0 -2.0 1e-06 
0.0 0.5748 0 -2.0 1e-06 
0.0 0.5749 0 -2.0 1e-06 
0.0 0.575 0 -2.0 1e-06 
0.0 0.5751 0 -2.0 1e-06 
0.0 0.5752 0 -2.0 1e-06 
0.0 0.5753 0 -2.0 1e-06 
0.0 0.5754 0 -2.0 1e-06 
0.0 0.5755 0 -2.0 1e-06 
0.0 0.5756 0 -2.0 1e-06 
0.0 0.5757 0 -2.0 1e-06 
0.0 0.5758 0 -2.0 1e-06 
0.0 0.5759 0 -2.0 1e-06 
0.0 0.576 0 -2.0 1e-06 
0.0 0.5761 0 -2.0 1e-06 
0.0 0.5762 0 -2.0 1e-06 
0.0 0.5763 0 -2.0 1e-06 
0.0 0.5764 0 -2.0 1e-06 
0.0 0.5765 0 -2.0 1e-06 
0.0 0.5766 0 -2.0 1e-06 
0.0 0.5767 0 -2.0 1e-06 
0.0 0.5768 0 -2.0 1e-06 
0.0 0.5769 0 -2.0 1e-06 
0.0 0.577 0 -2.0 1e-06 
0.0 0.5771 0 -2.0 1e-06 
0.0 0.5772 0 -2.0 1e-06 
0.0 0.5773 0 -2.0 1e-06 
0.0 0.5774 0 -2.0 1e-06 
0.0 0.5775 0 -2.0 1e-06 
0.0 0.5776 0 -2.0 1e-06 
0.0 0.5777 0 -2.0 1e-06 
0.0 0.5778 0 -2.0 1e-06 
0.0 0.5779 0 -2.0 1e-06 
0.0 0.578 0 -2.0 1e-06 
0.0 0.5781 0 -2.0 1e-06 
0.0 0.5782 0 -2.0 1e-06 
0.0 0.5783 0 -2.0 1e-06 
0.0 0.5784 0 -2.0 1e-06 
0.0 0.5785 0 -2.0 1e-06 
0.0 0.5786 0 -2.0 1e-06 
0.0 0.5787 0 -2.0 1e-06 
0.0 0.5788 0 -2.0 1e-06 
0.0 0.5789 0 -2.0 1e-06 
0.0 0.579 0 -2.0 1e-06 
0.0 0.5791 0 -2.0 1e-06 
0.0 0.5792 0 -2.0 1e-06 
0.0 0.5793 0 -2.0 1e-06 
0.0 0.5794 0 -2.0 1e-06 
0.0 0.5795 0 -2.0 1e-06 
0.0 0.5796 0 -2.0 1e-06 
0.0 0.5797 0 -2.0 1e-06 
0.0 0.5798 0 -2.0 1e-06 
0.0 0.5799 0 -2.0 1e-06 
0.0 0.58 0 -2.0 1e-06 
0.0 0.5801 0 -2.0 1e-06 
0.0 0.5802 0 -2.0 1e-06 
0.0 0.5803 0 -2.0 1e-06 
0.0 0.5804 0 -2.0 1e-06 
0.0 0.5805 0 -2.0 1e-06 
0.0 0.5806 0 -2.0 1e-06 
0.0 0.5807 0 -2.0 1e-06 
0.0 0.5808 0 -2.0 1e-06 
0.0 0.5809 0 -2.0 1e-06 
0.0 0.581 0 -2.0 1e-06 
0.0 0.5811 0 -2.0 1e-06 
0.0 0.5812 0 -2.0 1e-06 
0.0 0.5813 0 -2.0 1e-06 
0.0 0.5814 0 -2.0 1e-06 
0.0 0.5815 0 -2.0 1e-06 
0.0 0.5816 0 -2.0 1e-06 
0.0 0.5817 0 -2.0 1e-06 
0.0 0.5818 0 -2.0 1e-06 
0.0 0.5819 0 -2.0 1e-06 
0.0 0.582 0 -2.0 1e-06 
0.0 0.5821 0 -2.0 1e-06 
0.0 0.5822 0 -2.0 1e-06 
0.0 0.5823 0 -2.0 1e-06 
0.0 0.5824 0 -2.0 1e-06 
0.0 0.5825 0 -2.0 1e-06 
0.0 0.5826 0 -2.0 1e-06 
0.0 0.5827 0 -2.0 1e-06 
0.0 0.5828 0 -2.0 1e-06 
0.0 0.5829 0 -2.0 1e-06 
0.0 0.583 0 -2.0 1e-06 
0.0 0.5831 0 -2.0 1e-06 
0.0 0.5832 0 -2.0 1e-06 
0.0 0.5833 0 -2.0 1e-06 
0.0 0.5834 0 -2.0 1e-06 
0.0 0.5835 0 -2.0 1e-06 
0.0 0.5836 0 -2.0 1e-06 
0.0 0.5837 0 -2.0 1e-06 
0.0 0.5838 0 -2.0 1e-06 
0.0 0.5839 0 -2.0 1e-06 
0.0 0.584 0 -2.0 1e-06 
0.0 0.5841 0 -2.0 1e-06 
0.0 0.5842 0 -2.0 1e-06 
0.0 0.5843 0 -2.0 1e-06 
0.0 0.5844 0 -2.0 1e-06 
0.0 0.5845 0 -2.0 1e-06 
0.0 0.5846 0 -2.0 1e-06 
0.0 0.5847 0 -2.0 1e-06 
0.0 0.5848 0 -2.0 1e-06 
0.0 0.5849 0 -2.0 1e-06 
0.0 0.585 0 -2.0 1e-06 
0.0 0.5851 0 -2.0 1e-06 
0.0 0.5852 0 -2.0 1e-06 
0.0 0.5853 0 -2.0 1e-06 
0.0 0.5854 0 -2.0 1e-06 
0.0 0.5855 0 -2.0 1e-06 
0.0 0.5856 0 -2.0 1e-06 
0.0 0.5857 0 -2.0 1e-06 
0.0 0.5858 0 -2.0 1e-06 
0.0 0.5859 0 -2.0 1e-06 
0.0 0.586 0 -2.0 1e-06 
0.0 0.5861 0 -2.0 1e-06 
0.0 0.5862 0 -2.0 1e-06 
0.0 0.5863 0 -2.0 1e-06 
0.0 0.5864 0 -2.0 1e-06 
0.0 0.5865 0 -2.0 1e-06 
0.0 0.5866 0 -2.0 1e-06 
0.0 0.5867 0 -2.0 1e-06 
0.0 0.5868 0 -2.0 1e-06 
0.0 0.5869 0 -2.0 1e-06 
0.0 0.587 0 -2.0 1e-06 
0.0 0.5871 0 -2.0 1e-06 
0.0 0.5872 0 -2.0 1e-06 
0.0 0.5873 0 -2.0 1e-06 
0.0 0.5874 0 -2.0 1e-06 
0.0 0.5875 0 -2.0 1e-06 
0.0 0.5876 0 -2.0 1e-06 
0.0 0.5877 0 -2.0 1e-06 
0.0 0.5878 0 -2.0 1e-06 
0.0 0.5879 0 -2.0 1e-06 
0.0 0.588 0 -2.0 1e-06 
0.0 0.5881 0 -2.0 1e-06 
0.0 0.5882 0 -2.0 1e-06 
0.0 0.5883 0 -2.0 1e-06 
0.0 0.5884 0 -2.0 1e-06 
0.0 0.5885 0 -2.0 1e-06 
0.0 0.5886 0 -2.0 1e-06 
0.0 0.5887 0 -2.0 1e-06 
0.0 0.5888 0 -2.0 1e-06 
0.0 0.5889 0 -2.0 1e-06 
0.0 0.589 0 -2.0 1e-06 
0.0 0.5891 0 -2.0 1e-06 
0.0 0.5892 0 -2.0 1e-06 
0.0 0.5893 0 -2.0 1e-06 
0.0 0.5894 0 -2.0 1e-06 
0.0 0.5895 0 -2.0 1e-06 
0.0 0.5896 0 -2.0 1e-06 
0.0 0.5897 0 -2.0 1e-06 
0.0 0.5898 0 -2.0 1e-06 
0.0 0.5899 0 -2.0 1e-06 
0.0 0.59 0 -2.0 1e-06 
0.0 0.5901 0 -2.0 1e-06 
0.0 0.5902 0 -2.0 1e-06 
0.0 0.5903 0 -2.0 1e-06 
0.0 0.5904 0 -2.0 1e-06 
0.0 0.5905 0 -2.0 1e-06 
0.0 0.5906 0 -2.0 1e-06 
0.0 0.5907 0 -2.0 1e-06 
0.0 0.5908 0 -2.0 1e-06 
0.0 0.5909 0 -2.0 1e-06 
0.0 0.591 0 -2.0 1e-06 
0.0 0.5911 0 -2.0 1e-06 
0.0 0.5912 0 -2.0 1e-06 
0.0 0.5913 0 -2.0 1e-06 
0.0 0.5914 0 -2.0 1e-06 
0.0 0.5915 0 -2.0 1e-06 
0.0 0.5916 0 -2.0 1e-06 
0.0 0.5917 0 -2.0 1e-06 
0.0 0.5918 0 -2.0 1e-06 
0.0 0.5919 0 -2.0 1e-06 
0.0 0.592 0 -2.0 1e-06 
0.0 0.5921 0 -2.0 1e-06 
0.0 0.5922 0 -2.0 1e-06 
0.0 0.5923 0 -2.0 1e-06 
0.0 0.5924 0 -2.0 1e-06 
0.0 0.5925 0 -2.0 1e-06 
0.0 0.5926 0 -2.0 1e-06 
0.0 0.5927 0 -2.0 1e-06 
0.0 0.5928 0 -2.0 1e-06 
0.0 0.5929 0 -2.0 1e-06 
0.0 0.593 0 -2.0 1e-06 
0.0 0.5931 0 -2.0 1e-06 
0.0 0.5932 0 -2.0 1e-06 
0.0 0.5933 0 -2.0 1e-06 
0.0 0.5934 0 -2.0 1e-06 
0.0 0.5935 0 -2.0 1e-06 
0.0 0.5936 0 -2.0 1e-06 
0.0 0.5937 0 -2.0 1e-06 
0.0 0.5938 0 -2.0 1e-06 
0.0 0.5939 0 -2.0 1e-06 
0.0 0.594 0 -2.0 1e-06 
0.0 0.5941 0 -2.0 1e-06 
0.0 0.5942 0 -2.0 1e-06 
0.0 0.5943 0 -2.0 1e-06 
0.0 0.5944 0 -2.0 1e-06 
0.0 0.5945 0 -2.0 1e-06 
0.0 0.5946 0 -2.0 1e-06 
0.0 0.5947 0 -2.0 1e-06 
0.0 0.5948 0 -2.0 1e-06 
0.0 0.5949 0 -2.0 1e-06 
0.0 0.595 0 -2.0 1e-06 
0.0 0.5951 0 -2.0 1e-06 
0.0 0.5952 0 -2.0 1e-06 
0.0 0.5953 0 -2.0 1e-06 
0.0 0.5954 0 -2.0 1e-06 
0.0 0.5955 0 -2.0 1e-06 
0.0 0.5956 0 -2.0 1e-06 
0.0 0.5957 0 -2.0 1e-06 
0.0 0.5958 0 -2.0 1e-06 
0.0 0.5959 0 -2.0 1e-06 
0.0 0.596 0 -2.0 1e-06 
0.0 0.5961 0 -2.0 1e-06 
0.0 0.5962 0 -2.0 1e-06 
0.0 0.5963 0 -2.0 1e-06 
0.0 0.5964 0 -2.0 1e-06 
0.0 0.5965 0 -2.0 1e-06 
0.0 0.5966 0 -2.0 1e-06 
0.0 0.5967 0 -2.0 1e-06 
0.0 0.5968 0 -2.0 1e-06 
0.0 0.5969 0 -2.0 1e-06 
0.0 0.597 0 -2.0 1e-06 
0.0 0.5971 0 -2.0 1e-06 
0.0 0.5972 0 -2.0 1e-06 
0.0 0.5973 0 -2.0 1e-06 
0.0 0.5974 0 -2.0 1e-06 
0.0 0.5975 0 -2.0 1e-06 
0.0 0.5976 0 -2.0 1e-06 
0.0 0.5977 0 -2.0 1e-06 
0.0 0.5978 0 -2.0 1e-06 
0.0 0.5979 0 -2.0 1e-06 
0.0 0.598 0 -2.0 1e-06 
0.0 0.5981 0 -2.0 1e-06 
0.0 0.5982 0 -2.0 1e-06 
0.0 0.5983 0 -2.0 1e-06 
0.0 0.5984 0 -2.0 1e-06 
0.0 0.5985 0 -2.0 1e-06 
0.0 0.5986 0 -2.0 1e-06 
0.0 0.5987 0 -2.0 1e-06 
0.0 0.5988 0 -2.0 1e-06 
0.0 0.5989 0 -2.0 1e-06 
0.0 0.599 0 -2.0 1e-06 
0.0 0.5991 0 -2.0 1e-06 
0.0 0.5992 0 -2.0 1e-06 
0.0 0.5993 0 -2.0 1e-06 
0.0 0.5994 0 -2.0 1e-06 
0.0 0.5995 0 -2.0 1e-06 
0.0 0.5996 0 -2.0 1e-06 
0.0 0.5997 0 -2.0 1e-06 
0.0 0.5998 0 -2.0 1e-06 
0.0 0.5999 0 -2.0 1e-06 
0.0 0.6 0 -2.0 1e-06 
0.0 0.6001 0 -2.0 1e-06 
0.0 0.6002 0 -2.0 1e-06 
0.0 0.6003 0 -2.0 1e-06 
0.0 0.6004 0 -2.0 1e-06 
0.0 0.6005 0 -2.0 1e-06 
0.0 0.6006 0 -2.0 1e-06 
0.0 0.6007 0 -2.0 1e-06 
0.0 0.6008 0 -2.0 1e-06 
0.0 0.6009 0 -2.0 1e-06 
0.0 0.601 0 -2.0 1e-06 
0.0 0.6011 0 -2.0 1e-06 
0.0 0.6012 0 -2.0 1e-06 
0.0 0.6013 0 -2.0 1e-06 
0.0 0.6014 0 -2.0 1e-06 
0.0 0.6015 0 -2.0 1e-06 
0.0 0.6016 0 -2.0 1e-06 
0.0 0.6017 0 -2.0 1e-06 
0.0 0.6018 0 -2.0 1e-06 
0.0 0.6019 0 -2.0 1e-06 
0.0 0.602 0 -2.0 1e-06 
0.0 0.6021 0 -2.0 1e-06 
0.0 0.6022 0 -2.0 1e-06 
0.0 0.6023 0 -2.0 1e-06 
0.0 0.6024 0 -2.0 1e-06 
0.0 0.6025 0 -2.0 1e-06 
0.0 0.6026 0 -2.0 1e-06 
0.0 0.6027 0 -2.0 1e-06 
0.0 0.6028 0 -2.0 1e-06 
0.0 0.6029 0 -2.0 1e-06 
0.0 0.603 0 -2.0 1e-06 
0.0 0.6031 0 -2.0 1e-06 
0.0 0.6032 0 -2.0 1e-06 
0.0 0.6033 0 -2.0 1e-06 
0.0 0.6034 0 -2.0 1e-06 
0.0 0.6035 0 -2.0 1e-06 
0.0 0.6036 0 -2.0 1e-06 
0.0 0.6037 0 -2.0 1e-06 
0.0 0.6038 0 -2.0 1e-06 
0.0 0.6039 0 -2.0 1e-06 
0.0 0.604 0 -2.0 1e-06 
0.0 0.6041 0 -2.0 1e-06 
0.0 0.6042 0 -2.0 1e-06 
0.0 0.6043 0 -2.0 1e-06 
0.0 0.6044 0 -2.0 1e-06 
0.0 0.6045 0 -2.0 1e-06 
0.0 0.6046 0 -2.0 1e-06 
0.0 0.6047 0 -2.0 1e-06 
0.0 0.6048 0 -2.0 1e-06 
0.0 0.6049 0 -2.0 1e-06 
0.0 0.605 0 -2.0 1e-06 
0.0 0.6051 0 -2.0 1e-06 
0.0 0.6052 0 -2.0 1e-06 
0.0 0.6053 0 -2.0 1e-06 
0.0 0.6054 0 -2.0 1e-06 
0.0 0.6055 0 -2.0 1e-06 
0.0 0.6056 0 -2.0 1e-06 
0.0 0.6057 0 -2.0 1e-06 
0.0 0.6058 0 -2.0 1e-06 
0.0 0.6059 0 -2.0 1e-06 
0.0 0.606 0 -2.0 1e-06 
0.0 0.6061 0 -2.0 1e-06 
0.0 0.6062 0 -2.0 1e-06 
0.0 0.6063 0 -2.0 1e-06 
0.0 0.6064 0 -2.0 1e-06 
0.0 0.6065 0 -2.0 1e-06 
0.0 0.6066 0 -2.0 1e-06 
0.0 0.6067 0 -2.0 1e-06 
0.0 0.6068 0 -2.0 1e-06 
0.0 0.6069 0 -2.0 1e-06 
0.0 0.607 0 -2.0 1e-06 
0.0 0.6071 0 -2.0 1e-06 
0.0 0.6072 0 -2.0 1e-06 
0.0 0.6073 0 -2.0 1e-06 
0.0 0.6074 0 -2.0 1e-06 
0.0 0.6075 0 -2.0 1e-06 
0.0 0.6076 0 -2.0 1e-06 
0.0 0.6077 0 -2.0 1e-06 
0.0 0.6078 0 -2.0 1e-06 
0.0 0.6079 0 -2.0 1e-06 
0.0 0.608 0 -2.0 1e-06 
0.0 0.6081 0 -2.0 1e-06 
0.0 0.6082 0 -2.0 1e-06 
0.0 0.6083 0 -2.0 1e-06 
0.0 0.6084 0 -2.0 1e-06 
0.0 0.6085 0 -2.0 1e-06 
0.0 0.6086 0 -2.0 1e-06 
0.0 0.6087 0 -2.0 1e-06 
0.0 0.6088 0 -2.0 1e-06 
0.0 0.6089 0 -2.0 1e-06 
0.0 0.609 0 -2.0 1e-06 
0.0 0.6091 0 -2.0 1e-06 
0.0 0.6092 0 -2.0 1e-06 
0.0 0.6093 0 -2.0 1e-06 
0.0 0.6094 0 -2.0 1e-06 
0.0 0.6095 0 -2.0 1e-06 
0.0 0.6096 0 -2.0 1e-06 
0.0 0.6097 0 -2.0 1e-06 
0.0 0.6098 0 -2.0 1e-06 
0.0 0.6099 0 -2.0 1e-06 
0.0 0.61 0 -2.0 1e-06 
0.0 0.6101 0 -2.0 1e-06 
0.0 0.6102 0 -2.0 1e-06 
0.0 0.6103 0 -2.0 1e-06 
0.0 0.6104 0 -2.0 1e-06 
0.0 0.6105 0 -2.0 1e-06 
0.0 0.6106 0 -2.0 1e-06 
0.0 0.6107 0 -2.0 1e-06 
0.0 0.6108 0 -2.0 1e-06 
0.0 0.6109 0 -2.0 1e-06 
0.0 0.611 0 -2.0 1e-06 
0.0 0.6111 0 -2.0 1e-06 
0.0 0.6112 0 -2.0 1e-06 
0.0 0.6113 0 -2.0 1e-06 
0.0 0.6114 0 -2.0 1e-06 
0.0 0.6115 0 -2.0 1e-06 
0.0 0.6116 0 -2.0 1e-06 
0.0 0.6117 0 -2.0 1e-06 
0.0 0.6118 0 -2.0 1e-06 
0.0 0.6119 0 -2.0 1e-06 
0.0 0.612 0 -2.0 1e-06 
0.0 0.6121 0 -2.0 1e-06 
0.0 0.6122 0 -2.0 1e-06 
0.0 0.6123 0 -2.0 1e-06 
0.0 0.6124 0 -2.0 1e-06 
0.0 0.6125 0 -2.0 1e-06 
0.0 0.6126 0 -2.0 1e-06 
0.0 0.6127 0 -2.0 1e-06 
0.0 0.6128 0 -2.0 1e-06 
0.0 0.6129 0 -2.0 1e-06 
0.0 0.613 0 -2.0 1e-06 
0.0 0.6131 0 -2.0 1e-06 
0.0 0.6132 0 -2.0 1e-06 
0.0 0.6133 0 -2.0 1e-06 
0.0 0.6134 0 -2.0 1e-06 
0.0 0.6135 0 -2.0 1e-06 
0.0 0.6136 0 -2.0 1e-06 
0.0 0.6137 0 -2.0 1e-06 
0.0 0.6138 0 -2.0 1e-06 
0.0 0.6139 0 -2.0 1e-06 
0.0 0.614 0 -2.0 1e-06 
0.0 0.6141 0 -2.0 1e-06 
0.0 0.6142 0 -2.0 1e-06 
0.0 0.6143 0 -2.0 1e-06 
0.0 0.6144 0 -2.0 1e-06 
0.0 0.6145 0 -2.0 1e-06 
0.0 0.6146 0 -2.0 1e-06 
0.0 0.6147 0 -2.0 1e-06 
0.0 0.6148 0 -2.0 1e-06 
0.0 0.6149 0 -2.0 1e-06 
0.0 0.615 0 -2.0 1e-06 
0.0 0.6151 0 -2.0 1e-06 
0.0 0.6152 0 -2.0 1e-06 
0.0 0.6153 0 -2.0 1e-06 
0.0 0.6154 0 -2.0 1e-06 
0.0 0.6155 0 -2.0 1e-06 
0.0 0.6156 0 -2.0 1e-06 
0.0 0.6157 0 -2.0 1e-06 
0.0 0.6158 0 -2.0 1e-06 
0.0 0.6159 0 -2.0 1e-06 
0.0 0.616 0 -2.0 1e-06 
0.0 0.6161 0 -2.0 1e-06 
0.0 0.6162 0 -2.0 1e-06 
0.0 0.6163 0 -2.0 1e-06 
0.0 0.6164 0 -2.0 1e-06 
0.0 0.6165 0 -2.0 1e-06 
0.0 0.6166 0 -2.0 1e-06 
0.0 0.6167 0 -2.0 1e-06 
0.0 0.6168 0 -2.0 1e-06 
0.0 0.6169 0 -2.0 1e-06 
0.0 0.617 0 -2.0 1e-06 
0.0 0.6171 0 -2.0 1e-06 
0.0 0.6172 0 -2.0 1e-06 
0.0 0.6173 0 -2.0 1e-06 
0.0 0.6174 0 -2.0 1e-06 
0.0 0.6175 0 -2.0 1e-06 
0.0 0.6176 0 -2.0 1e-06 
0.0 0.6177 0 -2.0 1e-06 
0.0 0.6178 0 -2.0 1e-06 
0.0 0.6179 0 -2.0 1e-06 
0.0 0.618 0 -2.0 1e-06 
0.0 0.6181 0 -2.0 1e-06 
0.0 0.6182 0 -2.0 1e-06 
0.0 0.6183 0 -2.0 1e-06 
0.0 0.6184 0 -2.0 1e-06 
0.0 0.6185 0 -2.0 1e-06 
0.0 0.6186 0 -2.0 1e-06 
0.0 0.6187 0 -2.0 1e-06 
0.0 0.6188 0 -2.0 1e-06 
0.0 0.6189 0 -2.0 1e-06 
0.0 0.619 0 -2.0 1e-06 
0.0 0.6191 0 -2.0 1e-06 
0.0 0.6192 0 -2.0 1e-06 
0.0 0.6193 0 -2.0 1e-06 
0.0 0.6194 0 -2.0 1e-06 
0.0 0.6195 0 -2.0 1e-06 
0.0 0.6196 0 -2.0 1e-06 
0.0 0.6197 0 -2.0 1e-06 
0.0 0.6198 0 -2.0 1e-06 
0.0 0.6199 0 -2.0 1e-06 
0.0 0.62 0 -2.0 1e-06 
0.0 0.6201 0 -2.0 1e-06 
0.0 0.6202 0 -2.0 1e-06 
0.0 0.6203 0 -2.0 1e-06 
0.0 0.6204 0 -2.0 1e-06 
0.0 0.6205 0 -2.0 1e-06 
0.0 0.6206 0 -2.0 1e-06 
0.0 0.6207 0 -2.0 1e-06 
0.0 0.6208 0 -2.0 1e-06 
0.0 0.6209 0 -2.0 1e-06 
0.0 0.621 0 -2.0 1e-06 
0.0 0.6211 0 -2.0 1e-06 
0.0 0.6212 0 -2.0 1e-06 
0.0 0.6213 0 -2.0 1e-06 
0.0 0.6214 0 -2.0 1e-06 
0.0 0.6215 0 -2.0 1e-06 
0.0 0.6216 0 -2.0 1e-06 
0.0 0.6217 0 -2.0 1e-06 
0.0 0.6218 0 -2.0 1e-06 
0.0 0.6219 0 -2.0 1e-06 
0.0 0.622 0 -2.0 1e-06 
0.0 0.6221 0 -2.0 1e-06 
0.0 0.6222 0 -2.0 1e-06 
0.0 0.6223 0 -2.0 1e-06 
0.0 0.6224 0 -2.0 1e-06 
0.0 0.6225 0 -2.0 1e-06 
0.0 0.6226 0 -2.0 1e-06 
0.0 0.6227 0 -2.0 1e-06 
0.0 0.6228 0 -2.0 1e-06 
0.0 0.6229 0 -2.0 1e-06 
0.0 0.623 0 -2.0 1e-06 
0.0 0.6231 0 -2.0 1e-06 
0.0 0.6232 0 -2.0 1e-06 
0.0 0.6233 0 -2.0 1e-06 
0.0 0.6234 0 -2.0 1e-06 
0.0 0.6235 0 -2.0 1e-06 
0.0 0.6236 0 -2.0 1e-06 
0.0 0.6237 0 -2.0 1e-06 
0.0 0.6238 0 -2.0 1e-06 
0.0 0.6239 0 -2.0 1e-06 
0.0 0.624 0 -2.0 1e-06 
0.0 0.6241 0 -2.0 1e-06 
0.0 0.6242 0 -2.0 1e-06 
0.0 0.6243 0 -2.0 1e-06 
0.0 0.6244 0 -2.0 1e-06 
0.0 0.6245 0 -2.0 1e-06 
0.0 0.6246 0 -2.0 1e-06 
0.0 0.6247 0 -2.0 1e-06 
0.0 0.6248 0 -2.0 1e-06 
0.0 0.6249 0 -2.0 1e-06 
0.0 0.625 0 -2.0 1e-06 
0.0 0.6251 0 -2.0 1e-06 
0.0 0.6252 0 -2.0 1e-06 
0.0 0.6253 0 -2.0 1e-06 
0.0 0.6254 0 -2.0 1e-06 
0.0 0.6255 0 -2.0 1e-06 
0.0 0.6256 0 -2.0 1e-06 
0.0 0.6257 0 -2.0 1e-06 
0.0 0.6258 0 -2.0 1e-06 
0.0 0.6259 0 -2.0 1e-06 
0.0 0.626 0 -2.0 1e-06 
0.0 0.6261 0 -2.0 1e-06 
0.0 0.6262 0 -2.0 1e-06 
0.0 0.6263 0 -2.0 1e-06 
0.0 0.6264 0 -2.0 1e-06 
0.0 0.6265 0 -2.0 1e-06 
0.0 0.6266 0 -2.0 1e-06 
0.0 0.6267 0 -2.0 1e-06 
0.0 0.6268 0 -2.0 1e-06 
0.0 0.6269 0 -2.0 1e-06 
0.0 0.627 0 -2.0 1e-06 
0.0 0.6271 0 -2.0 1e-06 
0.0 0.6272 0 -2.0 1e-06 
0.0 0.6273 0 -2.0 1e-06 
0.0 0.6274 0 -2.0 1e-06 
0.0 0.6275 0 -2.0 1e-06 
0.0 0.6276 0 -2.0 1e-06 
0.0 0.6277 0 -2.0 1e-06 
0.0 0.6278 0 -2.0 1e-06 
0.0 0.6279 0 -2.0 1e-06 
0.0 0.628 0 -2.0 1e-06 
0.0 0.6281 0 -2.0 1e-06 
0.0 0.6282 0 -2.0 1e-06 
0.0 0.6283 0 -2.0 1e-06 
0.0 0.6284 0 -2.0 1e-06 
0.0 0.6285 0 -2.0 1e-06 
0.0 0.6286 0 -2.0 1e-06 
0.0 0.6287 0 -2.0 1e-06 
0.0 0.6288 0 -2.0 1e-06 
0.0 0.6289 0 -2.0 1e-06 
0.0 0.629 0 -2.0 1e-06 
0.0 0.6291 0 -2.0 1e-06 
0.0 0.6292 0 -2.0 1e-06 
0.0 0.6293 0 -2.0 1e-06 
0.0 0.6294 0 -2.0 1e-06 
0.0 0.6295 0 -2.0 1e-06 
0.0 0.6296 0 -2.0 1e-06 
0.0 0.6297 0 -2.0 1e-06 
0.0 0.6298 0 -2.0 1e-06 
0.0 0.6299 0 -2.0 1e-06 
0.0 0.63 0 -2.0 1e-06 
0.0 0.6301 0 -2.0 1e-06 
0.0 0.6302 0 -2.0 1e-06 
0.0 0.6303 0 -2.0 1e-06 
0.0 0.6304 0 -2.0 1e-06 
0.0 0.6305 0 -2.0 1e-06 
0.0 0.6306 0 -2.0 1e-06 
0.0 0.6307 0 -2.0 1e-06 
0.0 0.6308 0 -2.0 1e-06 
0.0 0.6309 0 -2.0 1e-06 
0.0 0.631 0 -2.0 1e-06 
0.0 0.6311 0 -2.0 1e-06 
0.0 0.6312 0 -2.0 1e-06 
0.0 0.6313 0 -2.0 1e-06 
0.0 0.6314 0 -2.0 1e-06 
0.0 0.6315 0 -2.0 1e-06 
0.0 0.6316 0 -2.0 1e-06 
0.0 0.6317 0 -2.0 1e-06 
0.0 0.6318 0 -2.0 1e-06 
0.0 0.6319 0 -2.0 1e-06 
0.0 0.632 0 -2.0 1e-06 
0.0 0.6321 0 -2.0 1e-06 
0.0 0.6322 0 -2.0 1e-06 
0.0 0.6323 0 -2.0 1e-06 
0.0 0.6324 0 -2.0 1e-06 
0.0 0.6325 0 -2.0 1e-06 
0.0 0.6326 0 -2.0 1e-06 
0.0 0.6327 0 -2.0 1e-06 
0.0 0.6328 0 -2.0 1e-06 
0.0 0.6329 0 -2.0 1e-06 
0.0 0.633 0 -2.0 1e-06 
0.0 0.6331 0 -2.0 1e-06 
0.0 0.6332 0 -2.0 1e-06 
0.0 0.6333 0 -2.0 1e-06 
0.0 0.6334 0 -2.0 1e-06 
0.0 0.6335 0 -2.0 1e-06 
0.0 0.6336 0 -2.0 1e-06 
0.0 0.6337 0 -2.0 1e-06 
0.0 0.6338 0 -2.0 1e-06 
0.0 0.6339 0 -2.0 1e-06 
0.0 0.634 0 -2.0 1e-06 
0.0 0.6341 0 -2.0 1e-06 
0.0 0.6342 0 -2.0 1e-06 
0.0 0.6343 0 -2.0 1e-06 
0.0 0.6344 0 -2.0 1e-06 
0.0 0.6345 0 -2.0 1e-06 
0.0 0.6346 0 -2.0 1e-06 
0.0 0.6347 0 -2.0 1e-06 
0.0 0.6348 0 -2.0 1e-06 
0.0 0.6349 0 -2.0 1e-06 
0.0 0.635 0 -2.0 1e-06 
0.0 0.6351 0 -2.0 1e-06 
0.0 0.6352 0 -2.0 1e-06 
0.0 0.6353 0 -2.0 1e-06 
0.0 0.6354 0 -2.0 1e-06 
0.0 0.6355 0 -2.0 1e-06 
0.0 0.6356 0 -2.0 1e-06 
0.0 0.6357 0 -2.0 1e-06 
0.0 0.6358 0 -2.0 1e-06 
0.0 0.6359 0 -2.0 1e-06 
0.0 0.636 0 -2.0 1e-06 
0.0 0.6361 0 -2.0 1e-06 
0.0 0.6362 0 -2.0 1e-06 
0.0 0.6363 0 -2.0 1e-06 
0.0 0.6364 0 -2.0 1e-06 
0.0 0.6365 0 -2.0 1e-06 
0.0 0.6366 0 -2.0 1e-06 
0.0 0.6367 0 -2.0 1e-06 
0.0 0.6368 0 -2.0 1e-06 
0.0 0.6369 0 -2.0 1e-06 
0.0 0.637 0 -2.0 1e-06 
0.0 0.6371 0 -2.0 1e-06 
0.0 0.6372 0 -2.0 1e-06 
0.0 0.6373 0 -2.0 1e-06 
0.0 0.6374 0 -2.0 1e-06 
0.0 0.6375 0 -2.0 1e-06 
0.0 0.6376 0 -2.0 1e-06 
0.0 0.6377 0 -2.0 1e-06 
0.0 0.6378 0 -2.0 1e-06 
0.0 0.6379 0 -2.0 1e-06 
0.0 0.638 0 -2.0 1e-06 
0.0 0.6381 0 -2.0 1e-06 
0.0 0.6382 0 -2.0 1e-06 
0.0 0.6383 0 -2.0 1e-06 
0.0 0.6384 0 -2.0 1e-06 
0.0 0.6385 0 -2.0 1e-06 
0.0 0.6386 0 -2.0 1e-06 
0.0 0.6387 0 -2.0 1e-06 
0.0 0.6388 0 -2.0 1e-06 
0.0 0.6389 0 -2.0 1e-06 
0.0 0.639 0 -2.0 1e-06 
0.0 0.6391 0 -2.0 1e-06 
0.0 0.6392 0 -2.0 1e-06 
0.0 0.6393 0 -2.0 1e-06 
0.0 0.6394 0 -2.0 1e-06 
0.0 0.6395 0 -2.0 1e-06 
0.0 0.6396 0 -2.0 1e-06 
0.0 0.6397 0 -2.0 1e-06 
0.0 0.6398 0 -2.0 1e-06 
0.0 0.6399 0 -2.0 1e-06 
0.0 0.64 0 -2.0 1e-06 
0.0 0.6401 0 -2.0 1e-06 
0.0 0.6402 0 -2.0 1e-06 
0.0 0.6403 0 -2.0 1e-06 
0.0 0.6404 0 -2.0 1e-06 
0.0 0.6405 0 -2.0 1e-06 
0.0 0.6406 0 -2.0 1e-06 
0.0 0.6407 0 -2.0 1e-06 
0.0 0.6408 0 -2.0 1e-06 
0.0 0.6409 0 -2.0 1e-06 
0.0 0.641 0 -2.0 1e-06 
0.0 0.6411 0 -2.0 1e-06 
0.0 0.6412 0 -2.0 1e-06 
0.0 0.6413 0 -2.0 1e-06 
0.0 0.6414 0 -2.0 1e-06 
0.0 0.6415 0 -2.0 1e-06 
0.0 0.6416 0 -2.0 1e-06 
0.0 0.6417 0 -2.0 1e-06 
0.0 0.6418 0 -2.0 1e-06 
0.0 0.6419 0 -2.0 1e-06 
0.0 0.642 0 -2.0 1e-06 
0.0 0.6421 0 -2.0 1e-06 
0.0 0.6422 0 -2.0 1e-06 
0.0 0.6423 0 -2.0 1e-06 
0.0 0.6424 0 -2.0 1e-06 
0.0 0.6425 0 -2.0 1e-06 
0.0 0.6426 0 -2.0 1e-06 
0.0 0.6427 0 -2.0 1e-06 
0.0 0.6428 0 -2.0 1e-06 
0.0 0.6429 0 -2.0 1e-06 
0.0 0.643 0 -2.0 1e-06 
0.0 0.6431 0 -2.0 1e-06 
0.0 0.6432 0 -2.0 1e-06 
0.0 0.6433 0 -2.0 1e-06 
0.0 0.6434 0 -2.0 1e-06 
0.0 0.6435 0 -2.0 1e-06 
0.0 0.6436 0 -2.0 1e-06 
0.0 0.6437 0 -2.0 1e-06 
0.0 0.6438 0 -2.0 1e-06 
0.0 0.6439 0 -2.0 1e-06 
0.0 0.644 0 -2.0 1e-06 
0.0 0.6441 0 -2.0 1e-06 
0.0 0.6442 0 -2.0 1e-06 
0.0 0.6443 0 -2.0 1e-06 
0.0 0.6444 0 -2.0 1e-06 
0.0 0.6445 0 -2.0 1e-06 
0.0 0.6446 0 -2.0 1e-06 
0.0 0.6447 0 -2.0 1e-06 
0.0 0.6448 0 -2.0 1e-06 
0.0 0.6449 0 -2.0 1e-06 
0.0 0.645 0 -2.0 1e-06 
0.0 0.6451 0 -2.0 1e-06 
0.0 0.6452 0 -2.0 1e-06 
0.0 0.6453 0 -2.0 1e-06 
0.0 0.6454 0 -2.0 1e-06 
0.0 0.6455 0 -2.0 1e-06 
0.0 0.6456 0 -2.0 1e-06 
0.0 0.6457 0 -2.0 1e-06 
0.0 0.6458 0 -2.0 1e-06 
0.0 0.6459 0 -2.0 1e-06 
0.0 0.646 0 -2.0 1e-06 
0.0 0.6461 0 -2.0 1e-06 
0.0 0.6462 0 -2.0 1e-06 
0.0 0.6463 0 -2.0 1e-06 
0.0 0.6464 0 -2.0 1e-06 
0.0 0.6465 0 -2.0 1e-06 
0.0 0.6466 0 -2.0 1e-06 
0.0 0.6467 0 -2.0 1e-06 
0.0 0.6468 0 -2.0 1e-06 
0.0 0.6469 0 -2.0 1e-06 
0.0 0.647 0 -2.0 1e-06 
0.0 0.6471 0 -2.0 1e-06 
0.0 0.6472 0 -2.0 1e-06 
0.0 0.6473 0 -2.0 1e-06 
0.0 0.6474 0 -2.0 1e-06 
0.0 0.6475 0 -2.0 1e-06 
0.0 0.6476 0 -2.0 1e-06 
0.0 0.6477 0 -2.0 1e-06 
0.0 0.6478 0 -2.0 1e-06 
0.0 0.6479 0 -2.0 1e-06 
0.0 0.648 0 -2.0 1e-06 
0.0 0.6481 0 -2.0 1e-06 
0.0 0.6482 0 -2.0 1e-06 
0.0 0.6483 0 -2.0 1e-06 
0.0 0.6484 0 -2.0 1e-06 
0.0 0.6485 0 -2.0 1e-06 
0.0 0.6486 0 -2.0 1e-06 
0.0 0.6487 0 -2.0 1e-06 
0.0 0.6488 0 -2.0 1e-06 
0.0 0.6489 0 -2.0 1e-06 
0.0 0.649 0 -2.0 1e-06 
0.0 0.6491 0 -2.0 1e-06 
0.0 0.6492 0 -2.0 1e-06 
0.0 0.6493 0 -2.0 1e-06 
0.0 0.6494 0 -2.0 1e-06 
0.0 0.6495 0 -2.0 1e-06 
0.0 0.6496 0 -2.0 1e-06 
0.0 0.6497 0 -2.0 1e-06 
0.0 0.6498 0 -2.0 1e-06 
0.0 0.6499 0 -2.0 1e-06 
0.0 0.65 0 -2.0 1e-06 
0.0 0.6501 0 -2.0 1e-06 
0.0 0.6502 0 -2.0 1e-06 
0.0 0.6503 0 -2.0 1e-06 
0.0 0.6504 0 -2.0 1e-06 
0.0 0.6505 0 -2.0 1e-06 
0.0 0.6506 0 -2.0 1e-06 
0.0 0.6507 0 -2.0 1e-06 
0.0 0.6508 0 -2.0 1e-06 
0.0 0.6509 0 -2.0 1e-06 
0.0 0.651 0 -2.0 1e-06 
0.0 0.6511 0 -2.0 1e-06 
0.0 0.6512 0 -2.0 1e-06 
0.0 0.6513 0 -2.0 1e-06 
0.0 0.6514 0 -2.0 1e-06 
0.0 0.6515 0 -2.0 1e-06 
0.0 0.6516 0 -2.0 1e-06 
0.0 0.6517 0 -2.0 1e-06 
0.0 0.6518 0 -2.0 1e-06 
0.0 0.6519 0 -2.0 1e-06 
0.0 0.652 0 -2.0 1e-06 
0.0 0.6521 0 -2.0 1e-06 
0.0 0.6522 0 -2.0 1e-06 
0.0 0.6523 0 -2.0 1e-06 
0.0 0.6524 0 -2.0 1e-06 
0.0 0.6525 0 -2.0 1e-06 
0.0 0.6526 0 -2.0 1e-06 
0.0 0.6527 0 -2.0 1e-06 
0.0 0.6528 0 -2.0 1e-06 
0.0 0.6529 0 -2.0 1e-06 
0.0 0.653 0 -2.0 1e-06 
0.0 0.6531 0 -2.0 1e-06 
0.0 0.6532 0 -2.0 1e-06 
0.0 0.6533 0 -2.0 1e-06 
0.0 0.6534 0 -2.0 1e-06 
0.0 0.6535 0 -2.0 1e-06 
0.0 0.6536 0 -2.0 1e-06 
0.0 0.6537 0 -2.0 1e-06 
0.0 0.6538 0 -2.0 1e-06 
0.0 0.6539 0 -2.0 1e-06 
0.0 0.654 0 -2.0 1e-06 
0.0 0.6541 0 -2.0 1e-06 
0.0 0.6542 0 -2.0 1e-06 
0.0 0.6543 0 -2.0 1e-06 
0.0 0.6544 0 -2.0 1e-06 
0.0 0.6545 0 -2.0 1e-06 
0.0 0.6546 0 -2.0 1e-06 
0.0 0.6547 0 -2.0 1e-06 
0.0 0.6548 0 -2.0 1e-06 
0.0 0.6549 0 -2.0 1e-06 
0.0 0.655 0 -2.0 1e-06 
0.0 0.6551 0 -2.0 1e-06 
0.0 0.6552 0 -2.0 1e-06 
0.0 0.6553 0 -2.0 1e-06 
0.0 0.6554 0 -2.0 1e-06 
0.0 0.6555 0 -2.0 1e-06 
0.0 0.6556 0 -2.0 1e-06 
0.0 0.6557 0 -2.0 1e-06 
0.0 0.6558 0 -2.0 1e-06 
0.0 0.6559 0 -2.0 1e-06 
0.0 0.656 0 -2.0 1e-06 
0.0 0.6561 0 -2.0 1e-06 
0.0 0.6562 0 -2.0 1e-06 
0.0 0.6563 0 -2.0 1e-06 
0.0 0.6564 0 -2.0 1e-06 
0.0 0.6565 0 -2.0 1e-06 
0.0 0.6566 0 -2.0 1e-06 
0.0 0.6567 0 -2.0 1e-06 
0.0 0.6568 0 -2.0 1e-06 
0.0 0.6569 0 -2.0 1e-06 
0.0 0.657 0 -2.0 1e-06 
0.0 0.6571 0 -2.0 1e-06 
0.0 0.6572 0 -2.0 1e-06 
0.0 0.6573 0 -2.0 1e-06 
0.0 0.6574 0 -2.0 1e-06 
0.0 0.6575 0 -2.0 1e-06 
0.0 0.6576 0 -2.0 1e-06 
0.0 0.6577 0 -2.0 1e-06 
0.0 0.6578 0 -2.0 1e-06 
0.0 0.6579 0 -2.0 1e-06 
0.0 0.658 0 -2.0 1e-06 
0.0 0.6581 0 -2.0 1e-06 
0.0 0.6582 0 -2.0 1e-06 
0.0 0.6583 0 -2.0 1e-06 
0.0 0.6584 0 -2.0 1e-06 
0.0 0.6585 0 -2.0 1e-06 
0.0 0.6586 0 -2.0 1e-06 
0.0 0.6587 0 -2.0 1e-06 
0.0 0.6588 0 -2.0 1e-06 
0.0 0.6589 0 -2.0 1e-06 
0.0 0.659 0 -2.0 1e-06 
0.0 0.6591 0 -2.0 1e-06 
0.0 0.6592 0 -2.0 1e-06 
0.0 0.6593 0 -2.0 1e-06 
0.0 0.6594 0 -2.0 1e-06 
0.0 0.6595 0 -2.0 1e-06 
0.0 0.6596 0 -2.0 1e-06 
0.0 0.6597 0 -2.0 1e-06 
0.0 0.6598 0 -2.0 1e-06 
0.0 0.6599 0 -2.0 1e-06 
0.0 0.66 0 -2.0 1e-06 
0.0 0.6601 0 -2.0 1e-06 
0.0 0.6602 0 -2.0 1e-06 
0.0 0.6603 0 -2.0 1e-06 
0.0 0.6604 0 -2.0 1e-06 
0.0 0.6605 0 -2.0 1e-06 
0.0 0.6606 0 -2.0 1e-06 
0.0 0.6607 0 -2.0 1e-06 
0.0 0.6608 0 -2.0 1e-06 
0.0 0.6609 0 -2.0 1e-06 
0.0 0.661 0 -2.0 1e-06 
0.0 0.6611 0 -2.0 1e-06 
0.0 0.6612 0 -2.0 1e-06 
0.0 0.6613 0 -2.0 1e-06 
0.0 0.6614 0 -2.0 1e-06 
0.0 0.6615 0 -2.0 1e-06 
0.0 0.6616 0 -2.0 1e-06 
0.0 0.6617 0 -2.0 1e-06 
0.0 0.6618 0 -2.0 1e-06 
0.0 0.6619 0 -2.0 1e-06 
0.0 0.662 0 -2.0 1e-06 
0.0 0.6621 0 -2.0 1e-06 
0.0 0.6622 0 -2.0 1e-06 
0.0 0.6623 0 -2.0 1e-06 
0.0 0.6624 0 -2.0 1e-06 
0.0 0.6625 0 -2.0 1e-06 
0.0 0.6626 0 -2.0 1e-06 
0.0 0.6627 0 -2.0 1e-06 
0.0 0.6628 0 -2.0 1e-06 
0.0 0.6629 0 -2.0 1e-06 
0.0 0.663 0 -2.0 1e-06 
0.0 0.6631 0 -2.0 1e-06 
0.0 0.6632 0 -2.0 1e-06 
0.0 0.6633 0 -2.0 1e-06 
0.0 0.6634 0 -2.0 1e-06 
0.0 0.6635 0 -2.0 1e-06 
0.0 0.6636 0 -2.0 1e-06 
0.0 0.6637 0 -2.0 1e-06 
0.0 0.6638 0 -2.0 1e-06 
0.0 0.6639 0 -2.0 1e-06 
0.0 0.664 0 -2.0 1e-06 
0.0 0.6641 0 -2.0 1e-06 
0.0 0.6642 0 -2.0 1e-06 
0.0 0.6643 0 -2.0 1e-06 
0.0 0.6644 0 -2.0 1e-06 
0.0 0.6645 0 -2.0 1e-06 
0.0 0.6646 0 -2.0 1e-06 
0.0 0.6647 0 -2.0 1e-06 
0.0 0.6648 0 -2.0 1e-06 
0.0 0.6649 0 -2.0 1e-06 
0.0 0.665 0 -2.0 1e-06 
0.0 0.6651 0 -2.0 1e-06 
0.0 0.6652 0 -2.0 1e-06 
0.0 0.6653 0 -2.0 1e-06 
0.0 0.6654 0 -2.0 1e-06 
0.0 0.6655 0 -2.0 1e-06 
0.0 0.6656 0 -2.0 1e-06 
0.0 0.6657 0 -2.0 1e-06 
0.0 0.6658 0 -2.0 1e-06 
0.0 0.6659 0 -2.0 1e-06 
0.0 0.666 0 -2.0 1e-06 
0.0 0.6661 0 -2.0 1e-06 
0.0 0.6662 0 -2.0 1e-06 
0.0 0.6663 0 -2.0 1e-06 
0.0 0.6664 0 -2.0 1e-06 
0.0 0.6665 0 -2.0 1e-06 
0.0 0.6666 0 -2.0 1e-06 
0.0 0.6667 0 -2.0 1e-06 
0.0 0.6668 0 -2.0 1e-06 
0.0 0.6669 0 -2.0 1e-06 
0.0 0.667 0 -2.0 1e-06 
0.0 0.6671 0 -2.0 1e-06 
0.0 0.6672 0 -2.0 1e-06 
0.0 0.6673 0 -2.0 1e-06 
0.0 0.6674 0 -2.0 1e-06 
0.0 0.6675 0 -2.0 1e-06 
0.0 0.6676 0 -2.0 1e-06 
0.0 0.6677 0 -2.0 1e-06 
0.0 0.6678 0 -2.0 1e-06 
0.0 0.6679 0 -2.0 1e-06 
0.0 0.668 0 -2.0 1e-06 
0.0 0.6681 0 -2.0 1e-06 
0.0 0.6682 0 -2.0 1e-06 
0.0 0.6683 0 -2.0 1e-06 
0.0 0.6684 0 -2.0 1e-06 
0.0 0.6685 0 -2.0 1e-06 
0.0 0.6686 0 -2.0 1e-06 
0.0 0.6687 0 -2.0 1e-06 
0.0 0.6688 0 -2.0 1e-06 
0.0 0.6689 0 -2.0 1e-06 
0.0 0.669 0 -2.0 1e-06 
0.0 0.6691 0 -2.0 1e-06 
0.0 0.6692 0 -2.0 1e-06 
0.0 0.6693 0 -2.0 1e-06 
0.0 0.6694 0 -2.0 1e-06 
0.0 0.6695 0 -2.0 1e-06 
0.0 0.6696 0 -2.0 1e-06 
0.0 0.6697 0 -2.0 1e-06 
0.0 0.6698 0 -2.0 1e-06 
0.0 0.6699 0 -2.0 1e-06 
0.0 0.67 0 -2.0 1e-06 
0.0 0.6701 0 -2.0 1e-06 
0.0 0.6702 0 -2.0 1e-06 
0.0 0.6703 0 -2.0 1e-06 
0.0 0.6704 0 -2.0 1e-06 
0.0 0.6705 0 -2.0 1e-06 
0.0 0.6706 0 -2.0 1e-06 
0.0 0.6707 0 -2.0 1e-06 
0.0 0.6708 0 -2.0 1e-06 
0.0 0.6709 0 -2.0 1e-06 
0.0 0.671 0 -2.0 1e-06 
0.0 0.6711 0 -2.0 1e-06 
0.0 0.6712 0 -2.0 1e-06 
0.0 0.6713 0 -2.0 1e-06 
0.0 0.6714 0 -2.0 1e-06 
0.0 0.6715 0 -2.0 1e-06 
0.0 0.6716 0 -2.0 1e-06 
0.0 0.6717 0 -2.0 1e-06 
0.0 0.6718 0 -2.0 1e-06 
0.0 0.6719 0 -2.0 1e-06 
0.0 0.672 0 -2.0 1e-06 
0.0 0.6721 0 -2.0 1e-06 
0.0 0.6722 0 -2.0 1e-06 
0.0 0.6723 0 -2.0 1e-06 
0.0 0.6724 0 -2.0 1e-06 
0.0 0.6725 0 -2.0 1e-06 
0.0 0.6726 0 -2.0 1e-06 
0.0 0.6727 0 -2.0 1e-06 
0.0 0.6728 0 -2.0 1e-06 
0.0 0.6729 0 -2.0 1e-06 
0.0 0.673 0 -2.0 1e-06 
0.0 0.6731 0 -2.0 1e-06 
0.0 0.6732 0 -2.0 1e-06 
0.0 0.6733 0 -2.0 1e-06 
0.0 0.6734 0 -2.0 1e-06 
0.0 0.6735 0 -2.0 1e-06 
0.0 0.6736 0 -2.0 1e-06 
0.0 0.6737 0 -2.0 1e-06 
0.0 0.6738 0 -2.0 1e-06 
0.0 0.6739 0 -2.0 1e-06 
0.0 0.674 0 -2.0 1e-06 
0.0 0.6741 0 -2.0 1e-06 
0.0 0.6742 0 -2.0 1e-06 
0.0 0.6743 0 -2.0 1e-06 
0.0 0.6744 0 -2.0 1e-06 
0.0 0.6745 0 -2.0 1e-06 
0.0 0.6746 0 -2.0 1e-06 
0.0 0.6747 0 -2.0 1e-06 
0.0 0.6748 0 -2.0 1e-06 
0.0 0.6749 0 -2.0 1e-06 
0.0 0.675 0 -2.0 1e-06 
0.0 0.6751 0 -2.0 1e-06 
0.0 0.6752 0 -2.0 1e-06 
0.0 0.6753 0 -2.0 1e-06 
0.0 0.6754 0 -2.0 1e-06 
0.0 0.6755 0 -2.0 1e-06 
0.0 0.6756 0 -2.0 1e-06 
0.0 0.6757 0 -2.0 1e-06 
0.0 0.6758 0 -2.0 1e-06 
0.0 0.6759 0 -2.0 1e-06 
0.0 0.676 0 -2.0 1e-06 
0.0 0.6761 0 -2.0 1e-06 
0.0 0.6762 0 -2.0 1e-06 
0.0 0.6763 0 -2.0 1e-06 
0.0 0.6764 0 -2.0 1e-06 
0.0 0.6765 0 -2.0 1e-06 
0.0 0.6766 0 -2.0 1e-06 
0.0 0.6767 0 -2.0 1e-06 
0.0 0.6768 0 -2.0 1e-06 
0.0 0.6769 0 -2.0 1e-06 
0.0 0.677 0 -2.0 1e-06 
0.0 0.6771 0 -2.0 1e-06 
0.0 0.6772 0 -2.0 1e-06 
0.0 0.6773 0 -2.0 1e-06 
0.0 0.6774 0 -2.0 1e-06 
0.0 0.6775 0 -2.0 1e-06 
0.0 0.6776 0 -2.0 1e-06 
0.0 0.6777 0 -2.0 1e-06 
0.0 0.6778 0 -2.0 1e-06 
0.0 0.6779 0 -2.0 1e-06 
0.0 0.678 0 -2.0 1e-06 
0.0 0.6781 0 -2.0 1e-06 
0.0 0.6782 0 -2.0 1e-06 
0.0 0.6783 0 -2.0 1e-06 
0.0 0.6784 0 -2.0 1e-06 
0.0 0.6785 0 -2.0 1e-06 
0.0 0.6786 0 -2.0 1e-06 
0.0 0.6787 0 -2.0 1e-06 
0.0 0.6788 0 -2.0 1e-06 
0.0 0.6789 0 -2.0 1e-06 
0.0 0.679 0 -2.0 1e-06 
0.0 0.6791 0 -2.0 1e-06 
0.0 0.6792 0 -2.0 1e-06 
0.0 0.6793 0 -2.0 1e-06 
0.0 0.6794 0 -2.0 1e-06 
0.0 0.6795 0 -2.0 1e-06 
0.0 0.6796 0 -2.0 1e-06 
0.0 0.6797 0 -2.0 1e-06 
0.0 0.6798 0 -2.0 1e-06 
0.0 0.6799 0 -2.0 1e-06 
0.0 0.68 0 -2.0 1e-06 
0.0 0.6801 0 -2.0 1e-06 
0.0 0.6802 0 -2.0 1e-06 
0.0 0.6803 0 -2.0 1e-06 
0.0 0.6804 0 -2.0 1e-06 
0.0 0.6805 0 -2.0 1e-06 
0.0 0.6806 0 -2.0 1e-06 
0.0 0.6807 0 -2.0 1e-06 
0.0 0.6808 0 -2.0 1e-06 
0.0 0.6809 0 -2.0 1e-06 
0.0 0.681 0 -2.0 1e-06 
0.0 0.6811 0 -2.0 1e-06 
0.0 0.6812 0 -2.0 1e-06 
0.0 0.6813 0 -2.0 1e-06 
0.0 0.6814 0 -2.0 1e-06 
0.0 0.6815 0 -2.0 1e-06 
0.0 0.6816 0 -2.0 1e-06 
0.0 0.6817 0 -2.0 1e-06 
0.0 0.6818 0 -2.0 1e-06 
0.0 0.6819 0 -2.0 1e-06 
0.0 0.682 0 -2.0 1e-06 
0.0 0.6821 0 -2.0 1e-06 
0.0 0.6822 0 -2.0 1e-06 
0.0 0.6823 0 -2.0 1e-06 
0.0 0.6824 0 -2.0 1e-06 
0.0 0.6825 0 -2.0 1e-06 
0.0 0.6826 0 -2.0 1e-06 
0.0 0.6827 0 -2.0 1e-06 
0.0 0.6828 0 -2.0 1e-06 
0.0 0.6829 0 -2.0 1e-06 
0.0 0.683 0 -2.0 1e-06 
0.0 0.6831 0 -2.0 1e-06 
0.0 0.6832 0 -2.0 1e-06 
0.0 0.6833 0 -2.0 1e-06 
0.0 0.6834 0 -2.0 1e-06 
0.0 0.6835 0 -2.0 1e-06 
0.0 0.6836 0 -2.0 1e-06 
0.0 0.6837 0 -2.0 1e-06 
0.0 0.6838 0 -2.0 1e-06 
0.0 0.6839 0 -2.0 1e-06 
0.0 0.684 0 -2.0 1e-06 
0.0 0.6841 0 -2.0 1e-06 
0.0 0.6842 0 -2.0 1e-06 
0.0 0.6843 0 -2.0 1e-06 
0.0 0.6844 0 -2.0 1e-06 
0.0 0.6845 0 -2.0 1e-06 
0.0 0.6846 0 -2.0 1e-06 
0.0 0.6847 0 -2.0 1e-06 
0.0 0.6848 0 -2.0 1e-06 
0.0 0.6849 0 -2.0 1e-06 
0.0 0.685 0 -2.0 1e-06 
0.0 0.6851 0 -2.0 1e-06 
0.0 0.6852 0 -2.0 1e-06 
0.0 0.6853 0 -2.0 1e-06 
0.0 0.6854 0 -2.0 1e-06 
0.0 0.6855 0 -2.0 1e-06 
0.0 0.6856 0 -2.0 1e-06 
0.0 0.6857 0 -2.0 1e-06 
0.0 0.6858 0 -2.0 1e-06 
0.0 0.6859 0 -2.0 1e-06 
0.0 0.686 0 -2.0 1e-06 
0.0 0.6861 0 -2.0 1e-06 
0.0 0.6862 0 -2.0 1e-06 
0.0 0.6863 0 -2.0 1e-06 
0.0 0.6864 0 -2.0 1e-06 
0.0 0.6865 0 -2.0 1e-06 
0.0 0.6866 0 -2.0 1e-06 
0.0 0.6867 0 -2.0 1e-06 
0.0 0.6868 0 -2.0 1e-06 
0.0 0.6869 0 -2.0 1e-06 
0.0 0.687 0 -2.0 1e-06 
0.0 0.6871 0 -2.0 1e-06 
0.0 0.6872 0 -2.0 1e-06 
0.0 0.6873 0 -2.0 1e-06 
0.0 0.6874 0 -2.0 1e-06 
0.0 0.6875 0 -2.0 1e-06 
0.0 0.6876 0 -2.0 1e-06 
0.0 0.6877 0 -2.0 1e-06 
0.0 0.6878 0 -2.0 1e-06 
0.0 0.6879 0 -2.0 1e-06 
0.0 0.688 0 -2.0 1e-06 
0.0 0.6881 0 -2.0 1e-06 
0.0 0.6882 0 -2.0 1e-06 
0.0 0.6883 0 -2.0 1e-06 
0.0 0.6884 0 -2.0 1e-06 
0.0 0.6885 0 -2.0 1e-06 
0.0 0.6886 0 -2.0 1e-06 
0.0 0.6887 0 -2.0 1e-06 
0.0 0.6888 0 -2.0 1e-06 
0.0 0.6889 0 -2.0 1e-06 
0.0 0.689 0 -2.0 1e-06 
0.0 0.6891 0 -2.0 1e-06 
0.0 0.6892 0 -2.0 1e-06 
0.0 0.6893 0 -2.0 1e-06 
0.0 0.6894 0 -2.0 1e-06 
0.0 0.6895 0 -2.0 1e-06 
0.0 0.6896 0 -2.0 1e-06 
0.0 0.6897 0 -2.0 1e-06 
0.0 0.6898 0 -2.0 1e-06 
0.0 0.6899 0 -2.0 1e-06 
0.0 0.69 0 -2.0 1e-06 
0.0 0.6901 0 -2.0 1e-06 
0.0 0.6902 0 -2.0 1e-06 
0.0 0.6903 0 -2.0 1e-06 
0.0 0.6904 0 -2.0 1e-06 
0.0 0.6905 0 -2.0 1e-06 
0.0 0.6906 0 -2.0 1e-06 
0.0 0.6907 0 -2.0 1e-06 
0.0 0.6908 0 -2.0 1e-06 
0.0 0.6909 0 -2.0 1e-06 
0.0 0.691 0 -2.0 1e-06 
0.0 0.6911 0 -2.0 1e-06 
0.0 0.6912 0 -2.0 1e-06 
0.0 0.6913 0 -2.0 1e-06 
0.0 0.6914 0 -2.0 1e-06 
0.0 0.6915 0 -2.0 1e-06 
0.0 0.6916 0 -2.0 1e-06 
0.0 0.6917 0 -2.0 1e-06 
0.0 0.6918 0 -2.0 1e-06 
0.0 0.6919 0 -2.0 1e-06 
0.0 0.692 0 -2.0 1e-06 
0.0 0.6921 0 -2.0 1e-06 
0.0 0.6922 0 -2.0 1e-06 
0.0 0.6923 0 -2.0 1e-06 
0.0 0.6924 0 -2.0 1e-06 
0.0 0.6925 0 -2.0 1e-06 
0.0 0.6926 0 -2.0 1e-06 
0.0 0.6927 0 -2.0 1e-06 
0.0 0.6928 0 -2.0 1e-06 
0.0 0.6929 0 -2.0 1e-06 
0.0 0.693 0 -2.0 1e-06 
0.0 0.6931 0 -2.0 1e-06 
0.0 0.6932 0 -2.0 1e-06 
0.0 0.6933 0 -2.0 1e-06 
0.0 0.6934 0 -2.0 1e-06 
0.0 0.6935 0 -2.0 1e-06 
0.0 0.6936 0 -2.0 1e-06 
0.0 0.6937 0 -2.0 1e-06 
0.0 0.6938 0 -2.0 1e-06 
0.0 0.6939 0 -2.0 1e-06 
0.0 0.694 0 -2.0 1e-06 
0.0 0.6941 0 -2.0 1e-06 
0.0 0.6942 0 -2.0 1e-06 
0.0 0.6943 0 -2.0 1e-06 
0.0 0.6944 0 -2.0 1e-06 
0.0 0.6945 0 -2.0 1e-06 
0.0 0.6946 0 -2.0 1e-06 
0.0 0.6947 0 -2.0 1e-06 
0.0 0.6948 0 -2.0 1e-06 
0.0 0.6949 0 -2.0 1e-06 
0.0 0.695 0 -2.0 1e-06 
0.0 0.6951 0 -2.0 1e-06 
0.0 0.6952 0 -2.0 1e-06 
0.0 0.6953 0 -2.0 1e-06 
0.0 0.6954 0 -2.0 1e-06 
0.0 0.6955 0 -2.0 1e-06 
0.0 0.6956 0 -2.0 1e-06 
0.0 0.6957 0 -2.0 1e-06 
0.0 0.6958 0 -2.0 1e-06 
0.0 0.6959 0 -2.0 1e-06 
0.0 0.696 0 -2.0 1e-06 
0.0 0.6961 0 -2.0 1e-06 
0.0 0.6962 0 -2.0 1e-06 
0.0 0.6963 0 -2.0 1e-06 
0.0 0.6964 0 -2.0 1e-06 
0.0 0.6965 0 -2.0 1e-06 
0.0 0.6966 0 -2.0 1e-06 
0.0 0.6967 0 -2.0 1e-06 
0.0 0.6968 0 -2.0 1e-06 
0.0 0.6969 0 -2.0 1e-06 
0.0 0.697 0 -2.0 1e-06 
0.0 0.6971 0 -2.0 1e-06 
0.0 0.6972 0 -2.0 1e-06 
0.0 0.6973 0 -2.0 1e-06 
0.0 0.6974 0 -2.0 1e-06 
0.0 0.6975 0 -2.0 1e-06 
0.0 0.6976 0 -2.0 1e-06 
0.0 0.6977 0 -2.0 1e-06 
0.0 0.6978 0 -2.0 1e-06 
0.0 0.6979 0 -2.0 1e-06 
0.0 0.698 0 -2.0 1e-06 
0.0 0.6981 0 -2.0 1e-06 
0.0 0.6982 0 -2.0 1e-06 
0.0 0.6983 0 -2.0 1e-06 
0.0 0.6984 0 -2.0 1e-06 
0.0 0.6985 0 -2.0 1e-06 
0.0 0.6986 0 -2.0 1e-06 
0.0 0.6987 0 -2.0 1e-06 
0.0 0.6988 0 -2.0 1e-06 
0.0 0.6989 0 -2.0 1e-06 
0.0 0.699 0 -2.0 1e-06 
0.0 0.6991 0 -2.0 1e-06 
0.0 0.6992 0 -2.0 1e-06 
0.0 0.6993 0 -2.0 1e-06 
0.0 0.6994 0 -2.0 1e-06 
0.0 0.6995 0 -2.0 1e-06 
0.0 0.6996 0 -2.0 1e-06 
0.0 0.6997 0 -2.0 1e-06 
0.0 0.6998 0 -2.0 1e-06 
0.0 0.6999 0 -2.0 1e-06 
0.0 0.7 0 -2.0 1e-06 
0.0 0.7001 0 -2.0 1e-06 
0.0 0.7002 0 -2.0 1e-06 
0.0 0.7003 0 -2.0 1e-06 
0.0 0.7004 0 -2.0 1e-06 
0.0 0.7005 0 -2.0 1e-06 
0.0 0.7006 0 -2.0 1e-06 
0.0 0.7007 0 -2.0 1e-06 
0.0 0.7008 0 -2.0 1e-06 
0.0 0.7009 0 -2.0 1e-06 
0.0 0.701 0 -2.0 1e-06 
0.0 0.7011 0 -2.0 1e-06 
0.0 0.7012 0 -2.0 1e-06 
0.0 0.7013 0 -2.0 1e-06 
0.0 0.7014 0 -2.0 1e-06 
0.0 0.7015 0 -2.0 1e-06 
0.0 0.7016 0 -2.0 1e-06 
0.0 0.7017 0 -2.0 1e-06 
0.0 0.7018 0 -2.0 1e-06 
0.0 0.7019 0 -2.0 1e-06 
0.0 0.702 0 -2.0 1e-06 
0.0 0.7021 0 -2.0 1e-06 
0.0 0.7022 0 -2.0 1e-06 
0.0 0.7023 0 -2.0 1e-06 
0.0 0.7024 0 -2.0 1e-06 
0.0 0.7025 0 -2.0 1e-06 
0.0 0.7026 0 -2.0 1e-06 
0.0 0.7027 0 -2.0 1e-06 
0.0 0.7028 0 -2.0 1e-06 
0.0 0.7029 0 -2.0 1e-06 
0.0 0.703 0 -2.0 1e-06 
0.0 0.7031 0 -2.0 1e-06 
0.0 0.7032 0 -2.0 1e-06 
0.0 0.7033 0 -2.0 1e-06 
0.0 0.7034 0 -2.0 1e-06 
0.0 0.7035 0 -2.0 1e-06 
0.0 0.7036 0 -2.0 1e-06 
0.0 0.7037 0 -2.0 1e-06 
0.0 0.7038 0 -2.0 1e-06 
0.0 0.7039 0 -2.0 1e-06 
0.0 0.704 0 -2.0 1e-06 
0.0 0.7041 0 -2.0 1e-06 
0.0 0.7042 0 -2.0 1e-06 
0.0 0.7043 0 -2.0 1e-06 
0.0 0.7044 0 -2.0 1e-06 
0.0 0.7045 0 -2.0 1e-06 
0.0 0.7046 0 -2.0 1e-06 
0.0 0.7047 0 -2.0 1e-06 
0.0 0.7048 0 -2.0 1e-06 
0.0 0.7049 0 -2.0 1e-06 
0.0 0.705 0 -2.0 1e-06 
0.0 0.7051 0 -2.0 1e-06 
0.0 0.7052 0 -2.0 1e-06 
0.0 0.7053 0 -2.0 1e-06 
0.0 0.7054 0 -2.0 1e-06 
0.0 0.7055 0 -2.0 1e-06 
0.0 0.7056 0 -2.0 1e-06 
0.0 0.7057 0 -2.0 1e-06 
0.0 0.7058 0 -2.0 1e-06 
0.0 0.7059 0 -2.0 1e-06 
0.0 0.706 0 -2.0 1e-06 
0.0 0.7061 0 -2.0 1e-06 
0.0 0.7062 0 -2.0 1e-06 
0.0 0.7063 0 -2.0 1e-06 
0.0 0.7064 0 -2.0 1e-06 
0.0 0.7065 0 -2.0 1e-06 
0.0 0.7066 0 -2.0 1e-06 
0.0 0.7067 0 -2.0 1e-06 
0.0 0.7068 0 -2.0 1e-06 
0.0 0.7069 0 -2.0 1e-06 
0.0 0.707 0 -2.0 1e-06 
0.0 0.7071 0 -2.0 1e-06 
0.0 0.7072 0 -2.0 1e-06 
0.0 0.7073 0 -2.0 1e-06 
0.0 0.7074 0 -2.0 1e-06 
0.0 0.7075 0 -2.0 1e-06 
0.0 0.7076 0 -2.0 1e-06 
0.0 0.7077 0 -2.0 1e-06 
0.0 0.7078 0 -2.0 1e-06 
0.0 0.7079 0 -2.0 1e-06 
0.0 0.708 0 -2.0 1e-06 
0.0 0.7081 0 -2.0 1e-06 
0.0 0.7082 0 -2.0 1e-06 
0.0 0.7083 0 -2.0 1e-06 
0.0 0.7084 0 -2.0 1e-06 
0.0 0.7085 0 -2.0 1e-06 
0.0 0.7086 0 -2.0 1e-06 
0.0 0.7087 0 -2.0 1e-06 
0.0 0.7088 0 -2.0 1e-06 
0.0 0.7089 0 -2.0 1e-06 
0.0 0.709 0 -2.0 1e-06 
0.0 0.7091 0 -2.0 1e-06 
0.0 0.7092 0 -2.0 1e-06 
0.0 0.7093 0 -2.0 1e-06 
0.0 0.7094 0 -2.0 1e-06 
0.0 0.7095 0 -2.0 1e-06 
0.0 0.7096 0 -2.0 1e-06 
0.0 0.7097 0 -2.0 1e-06 
0.0 0.7098 0 -2.0 1e-06 
0.0 0.7099 0 -2.0 1e-06 
0.0 0.71 0 -2.0 1e-06 
0.0 0.7101 0 -2.0 1e-06 
0.0 0.7102 0 -2.0 1e-06 
0.0 0.7103 0 -2.0 1e-06 
0.0 0.7104 0 -2.0 1e-06 
0.0 0.7105 0 -2.0 1e-06 
0.0 0.7106 0 -2.0 1e-06 
0.0 0.7107 0 -2.0 1e-06 
0.0 0.7108 0 -2.0 1e-06 
0.0 0.7109 0 -2.0 1e-06 
0.0 0.711 0 -2.0 1e-06 
0.0 0.7111 0 -2.0 1e-06 
0.0 0.7112 0 -2.0 1e-06 
0.0 0.7113 0 -2.0 1e-06 
0.0 0.7114 0 -2.0 1e-06 
0.0 0.7115 0 -2.0 1e-06 
0.0 0.7116 0 -2.0 1e-06 
0.0 0.7117 0 -2.0 1e-06 
0.0 0.7118 0 -2.0 1e-06 
0.0 0.7119 0 -2.0 1e-06 
0.0 0.712 0 -2.0 1e-06 
0.0 0.7121 0 -2.0 1e-06 
0.0 0.7122 0 -2.0 1e-06 
0.0 0.7123 0 -2.0 1e-06 
0.0 0.7124 0 -2.0 1e-06 
0.0 0.7125 0 -2.0 1e-06 
0.0 0.7126 0 -2.0 1e-06 
0.0 0.7127 0 -2.0 1e-06 
0.0 0.7128 0 -2.0 1e-06 
0.0 0.7129 0 -2.0 1e-06 
0.0 0.713 0 -2.0 1e-06 
0.0 0.7131 0 -2.0 1e-06 
0.0 0.7132 0 -2.0 1e-06 
0.0 0.7133 0 -2.0 1e-06 
0.0 0.7134 0 -2.0 1e-06 
0.0 0.7135 0 -2.0 1e-06 
0.0 0.7136 0 -2.0 1e-06 
0.0 0.7137 0 -2.0 1e-06 
0.0 0.7138 0 -2.0 1e-06 
0.0 0.7139 0 -2.0 1e-06 
0.0 0.714 0 -2.0 1e-06 
0.0 0.7141 0 -2.0 1e-06 
0.0 0.7142 0 -2.0 1e-06 
0.0 0.7143 0 -2.0 1e-06 
0.0 0.7144 0 -2.0 1e-06 
0.0 0.7145 0 -2.0 1e-06 
0.0 0.7146 0 -2.0 1e-06 
0.0 0.7147 0 -2.0 1e-06 
0.0 0.7148 0 -2.0 1e-06 
0.0 0.7149 0 -2.0 1e-06 
0.0 0.715 0 -2.0 1e-06 
0.0 0.7151 0 -2.0 1e-06 
0.0 0.7152 0 -2.0 1e-06 
0.0 0.7153 0 -2.0 1e-06 
0.0 0.7154 0 -2.0 1e-06 
0.0 0.7155 0 -2.0 1e-06 
0.0 0.7156 0 -2.0 1e-06 
0.0 0.7157 0 -2.0 1e-06 
0.0 0.7158 0 -2.0 1e-06 
0.0 0.7159 0 -2.0 1e-06 
0.0 0.716 0 -2.0 1e-06 
0.0 0.7161 0 -2.0 1e-06 
0.0 0.7162 0 -2.0 1e-06 
0.0 0.7163 0 -2.0 1e-06 
0.0 0.7164 0 -2.0 1e-06 
0.0 0.7165 0 -2.0 1e-06 
0.0 0.7166 0 -2.0 1e-06 
0.0 0.7167 0 -2.0 1e-06 
0.0 0.7168 0 -2.0 1e-06 
0.0 0.7169 0 -2.0 1e-06 
0.0 0.717 0 -2.0 1e-06 
0.0 0.7171 0 -2.0 1e-06 
0.0 0.7172 0 -2.0 1e-06 
0.0 0.7173 0 -2.0 1e-06 
0.0 0.7174 0 -2.0 1e-06 
0.0 0.7175 0 -2.0 1e-06 
0.0 0.7176 0 -2.0 1e-06 
0.0 0.7177 0 -2.0 1e-06 
0.0 0.7178 0 -2.0 1e-06 
0.0 0.7179 0 -2.0 1e-06 
0.0 0.718 0 -2.0 1e-06 
0.0 0.7181 0 -2.0 1e-06 
0.0 0.7182 0 -2.0 1e-06 
0.0 0.7183 0 -2.0 1e-06 
0.0 0.7184 0 -2.0 1e-06 
0.0 0.7185 0 -2.0 1e-06 
0.0 0.7186 0 -2.0 1e-06 
0.0 0.7187 0 -2.0 1e-06 
0.0 0.7188 0 -2.0 1e-06 
0.0 0.7189 0 -2.0 1e-06 
0.0 0.719 0 -2.0 1e-06 
0.0 0.7191 0 -2.0 1e-06 
0.0 0.7192 0 -2.0 1e-06 
0.0 0.7193 0 -2.0 1e-06 
0.0 0.7194 0 -2.0 1e-06 
0.0 0.7195 0 -2.0 1e-06 
0.0 0.7196 0 -2.0 1e-06 
0.0 0.7197 0 -2.0 1e-06 
0.0 0.7198 0 -2.0 1e-06 
0.0 0.7199 0 -2.0 1e-06 
0.0 0.72 0 -2.0 1e-06 
0.0 0.7201 0 -2.0 1e-06 
0.0 0.7202 0 -2.0 1e-06 
0.0 0.7203 0 -2.0 1e-06 
0.0 0.7204 0 -2.0 1e-06 
0.0 0.7205 0 -2.0 1e-06 
0.0 0.7206 0 -2.0 1e-06 
0.0 0.7207 0 -2.0 1e-06 
0.0 0.7208 0 -2.0 1e-06 
0.0 0.7209 0 -2.0 1e-06 
0.0 0.721 0 -2.0 1e-06 
0.0 0.7211 0 -2.0 1e-06 
0.0 0.7212 0 -2.0 1e-06 
0.0 0.7213 0 -2.0 1e-06 
0.0 0.7214 0 -2.0 1e-06 
0.0 0.7215 0 -2.0 1e-06 
0.0 0.7216 0 -2.0 1e-06 
0.0 0.7217 0 -2.0 1e-06 
0.0 0.7218 0 -2.0 1e-06 
0.0 0.7219 0 -2.0 1e-06 
0.0 0.722 0 -2.0 1e-06 
0.0 0.7221 0 -2.0 1e-06 
0.0 0.7222 0 -2.0 1e-06 
0.0 0.7223 0 -2.0 1e-06 
0.0 0.7224 0 -2.0 1e-06 
0.0 0.7225 0 -2.0 1e-06 
0.0 0.7226 0 -2.0 1e-06 
0.0 0.7227 0 -2.0 1e-06 
0.0 0.7228 0 -2.0 1e-06 
0.0 0.7229 0 -2.0 1e-06 
0.0 0.723 0 -2.0 1e-06 
0.0 0.7231 0 -2.0 1e-06 
0.0 0.7232 0 -2.0 1e-06 
0.0 0.7233 0 -2.0 1e-06 
0.0 0.7234 0 -2.0 1e-06 
0.0 0.7235 0 -2.0 1e-06 
0.0 0.7236 0 -2.0 1e-06 
0.0 0.7237 0 -2.0 1e-06 
0.0 0.7238 0 -2.0 1e-06 
0.0 0.7239 0 -2.0 1e-06 
0.0 0.724 0 -2.0 1e-06 
0.0 0.7241 0 -2.0 1e-06 
0.0 0.7242 0 -2.0 1e-06 
0.0 0.7243 0 -2.0 1e-06 
0.0 0.7244 0 -2.0 1e-06 
0.0 0.7245 0 -2.0 1e-06 
0.0 0.7246 0 -2.0 1e-06 
0.0 0.7247 0 -2.0 1e-06 
0.0 0.7248 0 -2.0 1e-06 
0.0 0.7249 0 -2.0 1e-06 
0.0 0.725 0 -2.0 1e-06 
0.0 0.7251 0 -2.0 1e-06 
0.0 0.7252 0 -2.0 1e-06 
0.0 0.7253 0 -2.0 1e-06 
0.0 0.7254 0 -2.0 1e-06 
0.0 0.7255 0 -2.0 1e-06 
0.0 0.7256 0 -2.0 1e-06 
0.0 0.7257 0 -2.0 1e-06 
0.0 0.7258 0 -2.0 1e-06 
0.0 0.7259 0 -2.0 1e-06 
0.0 0.726 0 -2.0 1e-06 
0.0 0.7261 0 -2.0 1e-06 
0.0 0.7262 0 -2.0 1e-06 
0.0 0.7263 0 -2.0 1e-06 
0.0 0.7264 0 -2.0 1e-06 
0.0 0.7265 0 -2.0 1e-06 
0.0 0.7266 0 -2.0 1e-06 
0.0 0.7267 0 -2.0 1e-06 
0.0 0.7268 0 -2.0 1e-06 
0.0 0.7269 0 -2.0 1e-06 
0.0 0.727 0 -2.0 1e-06 
0.0 0.7271 0 -2.0 1e-06 
0.0 0.7272 0 -2.0 1e-06 
0.0 0.7273 0 -2.0 1e-06 
0.0 0.7274 0 -2.0 1e-06 
0.0 0.7275 0 -2.0 1e-06 
0.0 0.7276 0 -2.0 1e-06 
0.0 0.7277 0 -2.0 1e-06 
0.0 0.7278 0 -2.0 1e-06 
0.0 0.7279 0 -2.0 1e-06 
0.0 0.728 0 -2.0 1e-06 
0.0 0.7281 0 -2.0 1e-06 
0.0 0.7282 0 -2.0 1e-06 
0.0 0.7283 0 -2.0 1e-06 
0.0 0.7284 0 -2.0 1e-06 
0.0 0.7285 0 -2.0 1e-06 
0.0 0.7286 0 -2.0 1e-06 
0.0 0.7287 0 -2.0 1e-06 
0.0 0.7288 0 -2.0 1e-06 
0.0 0.7289 0 -2.0 1e-06 
0.0 0.729 0 -2.0 1e-06 
0.0 0.7291 0 -2.0 1e-06 
0.0 0.7292 0 -2.0 1e-06 
0.0 0.7293 0 -2.0 1e-06 
0.0 0.7294 0 -2.0 1e-06 
0.0 0.7295 0 -2.0 1e-06 
0.0 0.7296 0 -2.0 1e-06 
0.0 0.7297 0 -2.0 1e-06 
0.0 0.7298 0 -2.0 1e-06 
0.0 0.7299 0 -2.0 1e-06 
0.0 0.73 0 -2.0 1e-06 
0.0 0.7301 0 -2.0 1e-06 
0.0 0.7302 0 -2.0 1e-06 
0.0 0.7303 0 -2.0 1e-06 
0.0 0.7304 0 -2.0 1e-06 
0.0 0.7305 0 -2.0 1e-06 
0.0 0.7306 0 -2.0 1e-06 
0.0 0.7307 0 -2.0 1e-06 
0.0 0.7308 0 -2.0 1e-06 
0.0 0.7309 0 -2.0 1e-06 
0.0 0.731 0 -2.0 1e-06 
0.0 0.7311 0 -2.0 1e-06 
0.0 0.7312 0 -2.0 1e-06 
0.0 0.7313 0 -2.0 1e-06 
0.0 0.7314 0 -2.0 1e-06 
0.0 0.7315 0 -2.0 1e-06 
0.0 0.7316 0 -2.0 1e-06 
0.0 0.7317 0 -2.0 1e-06 
0.0 0.7318 0 -2.0 1e-06 
0.0 0.7319 0 -2.0 1e-06 
0.0 0.732 0 -2.0 1e-06 
0.0 0.7321 0 -2.0 1e-06 
0.0 0.7322 0 -2.0 1e-06 
0.0 0.7323 0 -2.0 1e-06 
0.0 0.7324 0 -2.0 1e-06 
0.0 0.7325 0 -2.0 1e-06 
0.0 0.7326 0 -2.0 1e-06 
0.0 0.7327 0 -2.0 1e-06 
0.0 0.7328 0 -2.0 1e-06 
0.0 0.7329 0 -2.0 1e-06 
0.0 0.733 0 -2.0 1e-06 
0.0 0.7331 0 -2.0 1e-06 
0.0 0.7332 0 -2.0 1e-06 
0.0 0.7333 0 -2.0 1e-06 
0.0 0.7334 0 -2.0 1e-06 
0.0 0.7335 0 -2.0 1e-06 
0.0 0.7336 0 -2.0 1e-06 
0.0 0.7337 0 -2.0 1e-06 
0.0 0.7338 0 -2.0 1e-06 
0.0 0.7339 0 -2.0 1e-06 
0.0 0.734 0 -2.0 1e-06 
0.0 0.7341 0 -2.0 1e-06 
0.0 0.7342 0 -2.0 1e-06 
0.0 0.7343 0 -2.0 1e-06 
0.0 0.7344 0 -2.0 1e-06 
0.0 0.7345 0 -2.0 1e-06 
0.0 0.7346 0 -2.0 1e-06 
0.0 0.7347 0 -2.0 1e-06 
0.0 0.7348 0 -2.0 1e-06 
0.0 0.7349 0 -2.0 1e-06 
0.0 0.735 0 -2.0 1e-06 
0.0 0.7351 0 -2.0 1e-06 
0.0 0.7352 0 -2.0 1e-06 
0.0 0.7353 0 -2.0 1e-06 
0.0 0.7354 0 -2.0 1e-06 
0.0 0.7355 0 -2.0 1e-06 
0.0 0.7356 0 -2.0 1e-06 
0.0 0.7357 0 -2.0 1e-06 
0.0 0.7358 0 -2.0 1e-06 
0.0 0.7359 0 -2.0 1e-06 
0.0 0.736 0 -2.0 1e-06 
0.0 0.7361 0 -2.0 1e-06 
0.0 0.7362 0 -2.0 1e-06 
0.0 0.7363 0 -2.0 1e-06 
0.0 0.7364 0 -2.0 1e-06 
0.0 0.7365 0 -2.0 1e-06 
0.0 0.7366 0 -2.0 1e-06 
0.0 0.7367 0 -2.0 1e-06 
0.0 0.7368 0 -2.0 1e-06 
0.0 0.7369 0 -2.0 1e-06 
0.0 0.737 0 -2.0 1e-06 
0.0 0.7371 0 -2.0 1e-06 
0.0 0.7372 0 -2.0 1e-06 
0.0 0.7373 0 -2.0 1e-06 
0.0 0.7374 0 -2.0 1e-06 
0.0 0.7375 0 -2.0 1e-06 
0.0 0.7376 0 -2.0 1e-06 
0.0 0.7377 0 -2.0 1e-06 
0.0 0.7378 0 -2.0 1e-06 
0.0 0.7379 0 -2.0 1e-06 
0.0 0.738 0 -2.0 1e-06 
0.0 0.7381 0 -2.0 1e-06 
0.0 0.7382 0 -2.0 1e-06 
0.0 0.7383 0 -2.0 1e-06 
0.0 0.7384 0 -2.0 1e-06 
0.0 0.7385 0 -2.0 1e-06 
0.0 0.7386 0 -2.0 1e-06 
0.0 0.7387 0 -2.0 1e-06 
0.0 0.7388 0 -2.0 1e-06 
0.0 0.7389 0 -2.0 1e-06 
0.0 0.739 0 -2.0 1e-06 
0.0 0.7391 0 -2.0 1e-06 
0.0 0.7392 0 -2.0 1e-06 
0.0 0.7393 0 -2.0 1e-06 
0.0 0.7394 0 -2.0 1e-06 
0.0 0.7395 0 -2.0 1e-06 
0.0 0.7396 0 -2.0 1e-06 
0.0 0.7397 0 -2.0 1e-06 
0.0 0.7398 0 -2.0 1e-06 
0.0 0.7399 0 -2.0 1e-06 
0.0 0.74 0 -2.0 1e-06 
0.0 0.7401 0 -2.0 1e-06 
0.0 0.7402 0 -2.0 1e-06 
0.0 0.7403 0 -2.0 1e-06 
0.0 0.7404 0 -2.0 1e-06 
0.0 0.7405 0 -2.0 1e-06 
0.0 0.7406 0 -2.0 1e-06 
0.0 0.7407 0 -2.0 1e-06 
0.0 0.7408 0 -2.0 1e-06 
0.0 0.7409 0 -2.0 1e-06 
0.0 0.741 0 -2.0 1e-06 
0.0 0.7411 0 -2.0 1e-06 
0.0 0.7412 0 -2.0 1e-06 
0.0 0.7413 0 -2.0 1e-06 
0.0 0.7414 0 -2.0 1e-06 
0.0 0.7415 0 -2.0 1e-06 
0.0 0.7416 0 -2.0 1e-06 
0.0 0.7417 0 -2.0 1e-06 
0.0 0.7418 0 -2.0 1e-06 
0.0 0.7419 0 -2.0 1e-06 
0.0 0.742 0 -2.0 1e-06 
0.0 0.7421 0 -2.0 1e-06 
0.0 0.7422 0 -2.0 1e-06 
0.0 0.7423 0 -2.0 1e-06 
0.0 0.7424 0 -2.0 1e-06 
0.0 0.7425 0 -2.0 1e-06 
0.0 0.7426 0 -2.0 1e-06 
0.0 0.7427 0 -2.0 1e-06 
0.0 0.7428 0 -2.0 1e-06 
0.0 0.7429 0 -2.0 1e-06 
0.0 0.743 0 -2.0 1e-06 
0.0 0.7431 0 -2.0 1e-06 
0.0 0.7432 0 -2.0 1e-06 
0.0 0.7433 0 -2.0 1e-06 
0.0 0.7434 0 -2.0 1e-06 
0.0 0.7435 0 -2.0 1e-06 
0.0 0.7436 0 -2.0 1e-06 
0.0 0.7437 0 -2.0 1e-06 
0.0 0.7438 0 -2.0 1e-06 
0.0 0.7439 0 -2.0 1e-06 
0.0 0.744 0 -2.0 1e-06 
0.0 0.7441 0 -2.0 1e-06 
0.0 0.7442 0 -2.0 1e-06 
0.0 0.7443 0 -2.0 1e-06 
0.0 0.7444 0 -2.0 1e-06 
0.0 0.7445 0 -2.0 1e-06 
0.0 0.7446 0 -2.0 1e-06 
0.0 0.7447 0 -2.0 1e-06 
0.0 0.7448 0 -2.0 1e-06 
0.0 0.7449 0 -2.0 1e-06 
0.0 0.745 0 -2.0 1e-06 
0.0 0.7451 0 -2.0 1e-06 
0.0 0.7452 0 -2.0 1e-06 
0.0 0.7453 0 -2.0 1e-06 
0.0 0.7454 0 -2.0 1e-06 
0.0 0.7455 0 -2.0 1e-06 
0.0 0.7456 0 -2.0 1e-06 
0.0 0.7457 0 -2.0 1e-06 
0.0 0.7458 0 -2.0 1e-06 
0.0 0.7459 0 -2.0 1e-06 
0.0 0.746 0 -2.0 1e-06 
0.0 0.7461 0 -2.0 1e-06 
0.0 0.7462 0 -2.0 1e-06 
0.0 0.7463 0 -2.0 1e-06 
0.0 0.7464 0 -2.0 1e-06 
0.0 0.7465 0 -2.0 1e-06 
0.0 0.7466 0 -2.0 1e-06 
0.0 0.7467 0 -2.0 1e-06 
0.0 0.7468 0 -2.0 1e-06 
0.0 0.7469 0 -2.0 1e-06 
0.0 0.747 0 -2.0 1e-06 
0.0 0.7471 0 -2.0 1e-06 
0.0 0.7472 0 -2.0 1e-06 
0.0 0.7473 0 -2.0 1e-06 
0.0 0.7474 0 -2.0 1e-06 
0.0 0.7475 0 -2.0 1e-06 
0.0 0.7476 0 -2.0 1e-06 
0.0 0.7477 0 -2.0 1e-06 
0.0 0.7478 0 -2.0 1e-06 
0.0 0.7479 0 -2.0 1e-06 
0.0 0.748 0 -2.0 1e-06 
0.0 0.7481 0 -2.0 1e-06 
0.0 0.7482 0 -2.0 1e-06 
0.0 0.7483 0 -2.0 1e-06 
0.0 0.7484 0 -2.0 1e-06 
0.0 0.7485 0 -2.0 1e-06 
0.0 0.7486 0 -2.0 1e-06 
0.0 0.7487 0 -2.0 1e-06 
0.0 0.7488 0 -2.0 1e-06 
0.0 0.7489 0 -2.0 1e-06 
0.0 0.749 0 -2.0 1e-06 
0.0 0.7491 0 -2.0 1e-06 
0.0 0.7492 0 -2.0 1e-06 
0.0 0.7493 0 -2.0 1e-06 
0.0 0.7494 0 -2.0 1e-06 
0.0 0.7495 0 -2.0 1e-06 
0.0 0.7496 0 -2.0 1e-06 
0.0 0.7497 0 -2.0 1e-06 
0.0 0.7498 0 -2.0 1e-06 
0.0 0.7499 0 -2.0 1e-06 
0.0 0.75 0 -2.0 1e-06 
0.0 0.7501 0 -2.0 1e-06 
0.0 0.7502 0 -2.0 1e-06 
0.0 0.7503 0 -2.0 1e-06 
0.0 0.7504 0 -2.0 1e-06 
0.0 0.7505 0 -2.0 1e-06 
0.0 0.7506 0 -2.0 1e-06 
0.0 0.7507 0 -2.0 1e-06 
0.0 0.7508 0 -2.0 1e-06 
0.0 0.7509 0 -2.0 1e-06 
0.0 0.751 0 -2.0 1e-06 
0.0 0.7511 0 -2.0 1e-06 
0.0 0.7512 0 -2.0 1e-06 
0.0 0.7513 0 -2.0 1e-06 
0.0 0.7514 0 -2.0 1e-06 
0.0 0.7515 0 -2.0 1e-06 
0.0 0.7516 0 -2.0 1e-06 
0.0 0.7517 0 -2.0 1e-06 
0.0 0.7518 0 -2.0 1e-06 
0.0 0.7519 0 -2.0 1e-06 
0.0 0.752 0 -2.0 1e-06 
0.0 0.7521 0 -2.0 1e-06 
0.0 0.7522 0 -2.0 1e-06 
0.0 0.7523 0 -2.0 1e-06 
0.0 0.7524 0 -2.0 1e-06 
0.0 0.7525 0 -2.0 1e-06 
0.0 0.7526 0 -2.0 1e-06 
0.0 0.7527 0 -2.0 1e-06 
0.0 0.7528 0 -2.0 1e-06 
0.0 0.7529 0 -2.0 1e-06 
0.0 0.753 0 -2.0 1e-06 
0.0 0.7531 0 -2.0 1e-06 
0.0 0.7532 0 -2.0 1e-06 
0.0 0.7533 0 -2.0 1e-06 
0.0 0.7534 0 -2.0 1e-06 
0.0 0.7535 0 -2.0 1e-06 
0.0 0.7536 0 -2.0 1e-06 
0.0 0.7537 0 -2.0 1e-06 
0.0 0.7538 0 -2.0 1e-06 
0.0 0.7539 0 -2.0 1e-06 
0.0 0.754 0 -2.0 1e-06 
0.0 0.7541 0 -2.0 1e-06 
0.0 0.7542 0 -2.0 1e-06 
0.0 0.7543 0 -2.0 1e-06 
0.0 0.7544 0 -2.0 1e-06 
0.0 0.7545 0 -2.0 1e-06 
0.0 0.7546 0 -2.0 1e-06 
0.0 0.7547 0 -2.0 1e-06 
0.0 0.7548 0 -2.0 1e-06 
0.0 0.7549 0 -2.0 1e-06 
0.0 0.755 0 -2.0 1e-06 
0.0 0.7551 0 -2.0 1e-06 
0.0 0.7552 0 -2.0 1e-06 
0.0 0.7553 0 -2.0 1e-06 
0.0 0.7554 0 -2.0 1e-06 
0.0 0.7555 0 -2.0 1e-06 
0.0 0.7556 0 -2.0 1e-06 
0.0 0.7557 0 -2.0 1e-06 
0.0 0.7558 0 -2.0 1e-06 
0.0 0.7559 0 -2.0 1e-06 
0.0 0.756 0 -2.0 1e-06 
0.0 0.7561 0 -2.0 1e-06 
0.0 0.7562 0 -2.0 1e-06 
0.0 0.7563 0 -2.0 1e-06 
0.0 0.7564 0 -2.0 1e-06 
0.0 0.7565 0 -2.0 1e-06 
0.0 0.7566 0 -2.0 1e-06 
0.0 0.7567 0 -2.0 1e-06 
0.0 0.7568 0 -2.0 1e-06 
0.0 0.7569 0 -2.0 1e-06 
0.0 0.757 0 -2.0 1e-06 
0.0 0.7571 0 -2.0 1e-06 
0.0 0.7572 0 -2.0 1e-06 
0.0 0.7573 0 -2.0 1e-06 
0.0 0.7574 0 -2.0 1e-06 
0.0 0.7575 0 -2.0 1e-06 
0.0 0.7576 0 -2.0 1e-06 
0.0 0.7577 0 -2.0 1e-06 
0.0 0.7578 0 -2.0 1e-06 
0.0 0.7579 0 -2.0 1e-06 
0.0 0.758 0 -2.0 1e-06 
0.0 0.7581 0 -2.0 1e-06 
0.0 0.7582 0 -2.0 1e-06 
0.0 0.7583 0 -2.0 1e-06 
0.0 0.7584 0 -2.0 1e-06 
0.0 0.7585 0 -2.0 1e-06 
0.0 0.7586 0 -2.0 1e-06 
0.0 0.7587 0 -2.0 1e-06 
0.0 0.7588 0 -2.0 1e-06 
0.0 0.7589 0 -2.0 1e-06 
0.0 0.759 0 -2.0 1e-06 
0.0 0.7591 0 -2.0 1e-06 
0.0 0.7592 0 -2.0 1e-06 
0.0 0.7593 0 -2.0 1e-06 
0.0 0.7594 0 -2.0 1e-06 
0.0 0.7595 0 -2.0 1e-06 
0.0 0.7596 0 -2.0 1e-06 
0.0 0.7597 0 -2.0 1e-06 
0.0 0.7598 0 -2.0 1e-06 
0.0 0.7599 0 -2.0 1e-06 
0.0 0.76 0 -2.0 1e-06 
0.0 0.7601 0 -2.0 1e-06 
0.0 0.7602 0 -2.0 1e-06 
0.0 0.7603 0 -2.0 1e-06 
0.0 0.7604 0 -2.0 1e-06 
0.0 0.7605 0 -2.0 1e-06 
0.0 0.7606 0 -2.0 1e-06 
0.0 0.7607 0 -2.0 1e-06 
0.0 0.7608 0 -2.0 1e-06 
0.0 0.7609 0 -2.0 1e-06 
0.0 0.761 0 -2.0 1e-06 
0.0 0.7611 0 -2.0 1e-06 
0.0 0.7612 0 -2.0 1e-06 
0.0 0.7613 0 -2.0 1e-06 
0.0 0.7614 0 -2.0 1e-06 
0.0 0.7615 0 -2.0 1e-06 
0.0 0.7616 0 -2.0 1e-06 
0.0 0.7617 0 -2.0 1e-06 
0.0 0.7618 0 -2.0 1e-06 
0.0 0.7619 0 -2.0 1e-06 
0.0 0.762 0 -2.0 1e-06 
0.0 0.7621 0 -2.0 1e-06 
0.0 0.7622 0 -2.0 1e-06 
0.0 0.7623 0 -2.0 1e-06 
0.0 0.7624 0 -2.0 1e-06 
0.0 0.7625 0 -2.0 1e-06 
0.0 0.7626 0 -2.0 1e-06 
0.0 0.7627 0 -2.0 1e-06 
0.0 0.7628 0 -2.0 1e-06 
0.0 0.7629 0 -2.0 1e-06 
0.0 0.763 0 -2.0 1e-06 
0.0 0.7631 0 -2.0 1e-06 
0.0 0.7632 0 -2.0 1e-06 
0.0 0.7633 0 -2.0 1e-06 
0.0 0.7634 0 -2.0 1e-06 
0.0 0.7635 0 -2.0 1e-06 
0.0 0.7636 0 -2.0 1e-06 
0.0 0.7637 0 -2.0 1e-06 
0.0 0.7638 0 -2.0 1e-06 
0.0 0.7639 0 -2.0 1e-06 
0.0 0.764 0 -2.0 1e-06 
0.0 0.7641 0 -2.0 1e-06 
0.0 0.7642 0 -2.0 1e-06 
0.0 0.7643 0 -2.0 1e-06 
0.0 0.7644 0 -2.0 1e-06 
0.0 0.7645 0 -2.0 1e-06 
0.0 0.7646 0 -2.0 1e-06 
0.0 0.7647 0 -2.0 1e-06 
0.0 0.7648 0 -2.0 1e-06 
0.0 0.7649 0 -2.0 1e-06 
0.0 0.765 0 -2.0 1e-06 
0.0 0.7651 0 -2.0 1e-06 
0.0 0.7652 0 -2.0 1e-06 
0.0 0.7653 0 -2.0 1e-06 
0.0 0.7654 0 -2.0 1e-06 
0.0 0.7655 0 -2.0 1e-06 
0.0 0.7656 0 -2.0 1e-06 
0.0 0.7657 0 -2.0 1e-06 
0.0 0.7658 0 -2.0 1e-06 
0.0 0.7659 0 -2.0 1e-06 
0.0 0.766 0 -2.0 1e-06 
0.0 0.7661 0 -2.0 1e-06 
0.0 0.7662 0 -2.0 1e-06 
0.0 0.7663 0 -2.0 1e-06 
0.0 0.7664 0 -2.0 1e-06 
0.0 0.7665 0 -2.0 1e-06 
0.0 0.7666 0 -2.0 1e-06 
0.0 0.7667 0 -2.0 1e-06 
0.0 0.7668 0 -2.0 1e-06 
0.0 0.7669 0 -2.0 1e-06 
0.0 0.767 0 -2.0 1e-06 
0.0 0.7671 0 -2.0 1e-06 
0.0 0.7672 0 -2.0 1e-06 
0.0 0.7673 0 -2.0 1e-06 
0.0 0.7674 0 -2.0 1e-06 
0.0 0.7675 0 -2.0 1e-06 
0.0 0.7676 0 -2.0 1e-06 
0.0 0.7677 0 -2.0 1e-06 
0.0 0.7678 0 -2.0 1e-06 
0.0 0.7679 0 -2.0 1e-06 
0.0 0.768 0 -2.0 1e-06 
0.0 0.7681 0 -2.0 1e-06 
0.0 0.7682 0 -2.0 1e-06 
0.0 0.7683 0 -2.0 1e-06 
0.0 0.7684 0 -2.0 1e-06 
0.0 0.7685 0 -2.0 1e-06 
0.0 0.7686 0 -2.0 1e-06 
0.0 0.7687 0 -2.0 1e-06 
0.0 0.7688 0 -2.0 1e-06 
0.0 0.7689 0 -2.0 1e-06 
0.0 0.769 0 -2.0 1e-06 
0.0 0.7691 0 -2.0 1e-06 
0.0 0.7692 0 -2.0 1e-06 
0.0 0.7693 0 -2.0 1e-06 
0.0 0.7694 0 -2.0 1e-06 
0.0 0.7695 0 -2.0 1e-06 
0.0 0.7696 0 -2.0 1e-06 
0.0 0.7697 0 -2.0 1e-06 
0.0 0.7698 0 -2.0 1e-06 
0.0 0.7699 0 -2.0 1e-06 
0.0 0.77 0 -2.0 1e-06 
0.0 0.7701 0 -2.0 1e-06 
0.0 0.7702 0 -2.0 1e-06 
0.0 0.7703 0 -2.0 1e-06 
0.0 0.7704 0 -2.0 1e-06 
0.0 0.7705 0 -2.0 1e-06 
0.0 0.7706 0 -2.0 1e-06 
0.0 0.7707 0 -2.0 1e-06 
0.0 0.7708 0 -2.0 1e-06 
0.0 0.7709 0 -2.0 1e-06 
0.0 0.771 0 -2.0 1e-06 
0.0 0.7711 0 -2.0 1e-06 
0.0 0.7712 0 -2.0 1e-06 
0.0 0.7713 0 -2.0 1e-06 
0.0 0.7714 0 -2.0 1e-06 
0.0 0.7715 0 -2.0 1e-06 
0.0 0.7716 0 -2.0 1e-06 
0.0 0.7717 0 -2.0 1e-06 
0.0 0.7718 0 -2.0 1e-06 
0.0 0.7719 0 -2.0 1e-06 
0.0 0.772 0 -2.0 1e-06 
0.0 0.7721 0 -2.0 1e-06 
0.0 0.7722 0 -2.0 1e-06 
0.0 0.7723 0 -2.0 1e-06 
0.0 0.7724 0 -2.0 1e-06 
0.0 0.7725 0 -2.0 1e-06 
0.0 0.7726 0 -2.0 1e-06 
0.0 0.7727 0 -2.0 1e-06 
0.0 0.7728 0 -2.0 1e-06 
0.0 0.7729 0 -2.0 1e-06 
0.0 0.773 0 -2.0 1e-06 
0.0 0.7731 0 -2.0 1e-06 
0.0 0.7732 0 -2.0 1e-06 
0.0 0.7733 0 -2.0 1e-06 
0.0 0.7734 0 -2.0 1e-06 
0.0 0.7735 0 -2.0 1e-06 
0.0 0.7736 0 -2.0 1e-06 
0.0 0.7737 0 -2.0 1e-06 
0.0 0.7738 0 -2.0 1e-06 
0.0 0.7739 0 -2.0 1e-06 
0.0 0.774 0 -2.0 1e-06 
0.0 0.7741 0 -2.0 1e-06 
0.0 0.7742 0 -2.0 1e-06 
0.0 0.7743 0 -2.0 1e-06 
0.0 0.7744 0 -2.0 1e-06 
0.0 0.7745 0 -2.0 1e-06 
0.0 0.7746 0 -2.0 1e-06 
0.0 0.7747 0 -2.0 1e-06 
0.0 0.7748 0 -2.0 1e-06 
0.0 0.7749 0 -2.0 1e-06 
0.0 0.775 0 -2.0 1e-06 
0.0 0.7751 0 -2.0 1e-06 
0.0 0.7752 0 -2.0 1e-06 
0.0 0.7753 0 -2.0 1e-06 
0.0 0.7754 0 -2.0 1e-06 
0.0 0.7755 0 -2.0 1e-06 
0.0 0.7756 0 -2.0 1e-06 
0.0 0.7757 0 -2.0 1e-06 
0.0 0.7758 0 -2.0 1e-06 
0.0 0.7759 0 -2.0 1e-06 
0.0 0.776 0 -2.0 1e-06 
0.0 0.7761 0 -2.0 1e-06 
0.0 0.7762 0 -2.0 1e-06 
0.0 0.7763 0 -2.0 1e-06 
0.0 0.7764 0 -2.0 1e-06 
0.0 0.7765 0 -2.0 1e-06 
0.0 0.7766 0 -2.0 1e-06 
0.0 0.7767 0 -2.0 1e-06 
0.0 0.7768 0 -2.0 1e-06 
0.0 0.7769 0 -2.0 1e-06 
0.0 0.777 0 -2.0 1e-06 
0.0 0.7771 0 -2.0 1e-06 
0.0 0.7772 0 -2.0 1e-06 
0.0 0.7773 0 -2.0 1e-06 
0.0 0.7774 0 -2.0 1e-06 
0.0 0.7775 0 -2.0 1e-06 
0.0 0.7776 0 -2.0 1e-06 
0.0 0.7777 0 -2.0 1e-06 
0.0 0.7778 0 -2.0 1e-06 
0.0 0.7779 0 -2.0 1e-06 
0.0 0.778 0 -2.0 1e-06 
0.0 0.7781 0 -2.0 1e-06 
0.0 0.7782 0 -2.0 1e-06 
0.0 0.7783 0 -2.0 1e-06 
0.0 0.7784 0 -2.0 1e-06 
0.0 0.7785 0 -2.0 1e-06 
0.0 0.7786 0 -2.0 1e-06 
0.0 0.7787 0 -2.0 1e-06 
0.0 0.7788 0 -2.0 1e-06 
0.0 0.7789 0 -2.0 1e-06 
0.0 0.779 0 -2.0 1e-06 
0.0 0.7791 0 -2.0 1e-06 
0.0 0.7792 0 -2.0 1e-06 
0.0 0.7793 0 -2.0 1e-06 
0.0 0.7794 0 -2.0 1e-06 
0.0 0.7795 0 -2.0 1e-06 
0.0 0.7796 0 -2.0 1e-06 
0.0 0.7797 0 -2.0 1e-06 
0.0 0.7798 0 -2.0 1e-06 
0.0 0.7799 0 -2.0 1e-06 
0.0 0.78 0 -2.0 1e-06 
0.0 0.7801 0 -2.0 1e-06 
0.0 0.7802 0 -2.0 1e-06 
0.0 0.7803 0 -2.0 1e-06 
0.0 0.7804 0 -2.0 1e-06 
0.0 0.7805 0 -2.0 1e-06 
0.0 0.7806 0 -2.0 1e-06 
0.0 0.7807 0 -2.0 1e-06 
0.0 0.7808 0 -2.0 1e-06 
0.0 0.7809 0 -2.0 1e-06 
0.0 0.781 0 -2.0 1e-06 
0.0 0.7811 0 -2.0 1e-06 
0.0 0.7812 0 -2.0 1e-06 
0.0 0.7813 0 -2.0 1e-06 
0.0 0.7814 0 -2.0 1e-06 
0.0 0.7815 0 -2.0 1e-06 
0.0 0.7816 0 -2.0 1e-06 
0.0 0.7817 0 -2.0 1e-06 
0.0 0.7818 0 -2.0 1e-06 
0.0 0.7819 0 -2.0 1e-06 
0.0 0.782 0 -2.0 1e-06 
0.0 0.7821 0 -2.0 1e-06 
0.0 0.7822 0 -2.0 1e-06 
0.0 0.7823 0 -2.0 1e-06 
0.0 0.7824 0 -2.0 1e-06 
0.0 0.7825 0 -2.0 1e-06 
0.0 0.7826 0 -2.0 1e-06 
0.0 0.7827 0 -2.0 1e-06 
0.0 0.7828 0 -2.0 1e-06 
0.0 0.7829 0 -2.0 1e-06 
0.0 0.783 0 -2.0 1e-06 
0.0 0.7831 0 -2.0 1e-06 
0.0 0.7832 0 -2.0 1e-06 
0.0 0.7833 0 -2.0 1e-06 
0.0 0.7834 0 -2.0 1e-06 
0.0 0.7835 0 -2.0 1e-06 
0.0 0.7836 0 -2.0 1e-06 
0.0 0.7837 0 -2.0 1e-06 
0.0 0.7838 0 -2.0 1e-06 
0.0 0.7839 0 -2.0 1e-06 
0.0 0.784 0 -2.0 1e-06 
0.0 0.7841 0 -2.0 1e-06 
0.0 0.7842 0 -2.0 1e-06 
0.0 0.7843 0 -2.0 1e-06 
0.0 0.7844 0 -2.0 1e-06 
0.0 0.7845 0 -2.0 1e-06 
0.0 0.7846 0 -2.0 1e-06 
0.0 0.7847 0 -2.0 1e-06 
0.0 0.7848 0 -2.0 1e-06 
0.0 0.7849 0 -2.0 1e-06 
0.0 0.785 0 -2.0 1e-06 
0.0 0.7851 0 -2.0 1e-06 
0.0 0.7852 0 -2.0 1e-06 
0.0 0.7853 0 -2.0 1e-06 
0.0 0.7854 0 -2.0 1e-06 
0.0 0.7855 0 -2.0 1e-06 
0.0 0.7856 0 -2.0 1e-06 
0.0 0.7857 0 -2.0 1e-06 
0.0 0.7858 0 -2.0 1e-06 
0.0 0.7859 0 -2.0 1e-06 
0.0 0.786 0 -2.0 1e-06 
0.0 0.7861 0 -2.0 1e-06 
0.0 0.7862 0 -2.0 1e-06 
0.0 0.7863 0 -2.0 1e-06 
0.0 0.7864 0 -2.0 1e-06 
0.0 0.7865 0 -2.0 1e-06 
0.0 0.7866 0 -2.0 1e-06 
0.0 0.7867 0 -2.0 1e-06 
0.0 0.7868 0 -2.0 1e-06 
0.0 0.7869 0 -2.0 1e-06 
0.0 0.787 0 -2.0 1e-06 
0.0 0.7871 0 -2.0 1e-06 
0.0 0.7872 0 -2.0 1e-06 
0.0 0.7873 0 -2.0 1e-06 
0.0 0.7874 0 -2.0 1e-06 
0.0 0.7875 0 -2.0 1e-06 
0.0 0.7876 0 -2.0 1e-06 
0.0 0.7877 0 -2.0 1e-06 
0.0 0.7878 0 -2.0 1e-06 
0.0 0.7879 0 -2.0 1e-06 
0.0 0.788 0 -2.0 1e-06 
0.0 0.7881 0 -2.0 1e-06 
0.0 0.7882 0 -2.0 1e-06 
0.0 0.7883 0 -2.0 1e-06 
0.0 0.7884 0 -2.0 1e-06 
0.0 0.7885 0 -2.0 1e-06 
0.0 0.7886 0 -2.0 1e-06 
0.0 0.7887 0 -2.0 1e-06 
0.0 0.7888 0 -2.0 1e-06 
0.0 0.7889 0 -2.0 1e-06 
0.0 0.789 0 -2.0 1e-06 
0.0 0.7891 0 -2.0 1e-06 
0.0 0.7892 0 -2.0 1e-06 
0.0 0.7893 0 -2.0 1e-06 
0.0 0.7894 0 -2.0 1e-06 
0.0 0.7895 0 -2.0 1e-06 
0.0 0.7896 0 -2.0 1e-06 
0.0 0.7897 0 -2.0 1e-06 
0.0 0.7898 0 -2.0 1e-06 
0.0 0.7899 0 -2.0 1e-06 
0.0 0.79 0 -2.0 1e-06 
0.0 0.7901 0 -2.0 1e-06 
0.0 0.7902 0 -2.0 1e-06 
0.0 0.7903 0 -2.0 1e-06 
0.0 0.7904 0 -2.0 1e-06 
0.0 0.7905 0 -2.0 1e-06 
0.0 0.7906 0 -2.0 1e-06 
0.0 0.7907 0 -2.0 1e-06 
0.0 0.7908 0 -2.0 1e-06 
0.0 0.7909 0 -2.0 1e-06 
0.0 0.791 0 -2.0 1e-06 
0.0 0.7911 0 -2.0 1e-06 
0.0 0.7912 0 -2.0 1e-06 
0.0 0.7913 0 -2.0 1e-06 
0.0 0.7914 0 -2.0 1e-06 
0.0 0.7915 0 -2.0 1e-06 
0.0 0.7916 0 -2.0 1e-06 
0.0 0.7917 0 -2.0 1e-06 
0.0 0.7918 0 -2.0 1e-06 
0.0 0.7919 0 -2.0 1e-06 
0.0 0.792 0 -2.0 1e-06 
0.0 0.7921 0 -2.0 1e-06 
0.0 0.7922 0 -2.0 1e-06 
0.0 0.7923 0 -2.0 1e-06 
0.0 0.7924 0 -2.0 1e-06 
0.0 0.7925 0 -2.0 1e-06 
0.0 0.7926 0 -2.0 1e-06 
0.0 0.7927 0 -2.0 1e-06 
0.0 0.7928 0 -2.0 1e-06 
0.0 0.7929 0 -2.0 1e-06 
0.0 0.793 0 -2.0 1e-06 
0.0 0.7931 0 -2.0 1e-06 
0.0 0.7932 0 -2.0 1e-06 
0.0 0.7933 0 -2.0 1e-06 
0.0 0.7934 0 -2.0 1e-06 
0.0 0.7935 0 -2.0 1e-06 
0.0 0.7936 0 -2.0 1e-06 
0.0 0.7937 0 -2.0 1e-06 
0.0 0.7938 0 -2.0 1e-06 
0.0 0.7939 0 -2.0 1e-06 
0.0 0.794 0 -2.0 1e-06 
0.0 0.7941 0 -2.0 1e-06 
0.0 0.7942 0 -2.0 1e-06 
0.0 0.7943 0 -2.0 1e-06 
0.0 0.7944 0 -2.0 1e-06 
0.0 0.7945 0 -2.0 1e-06 
0.0 0.7946 0 -2.0 1e-06 
0.0 0.7947 0 -2.0 1e-06 
0.0 0.7948 0 -2.0 1e-06 
0.0 0.7949 0 -2.0 1e-06 
0.0 0.795 0 -2.0 1e-06 
0.0 0.7951 0 -2.0 1e-06 
0.0 0.7952 0 -2.0 1e-06 
0.0 0.7953 0 -2.0 1e-06 
0.0 0.7954 0 -2.0 1e-06 
0.0 0.7955 0 -2.0 1e-06 
0.0 0.7956 0 -2.0 1e-06 
0.0 0.7957 0 -2.0 1e-06 
0.0 0.7958 0 -2.0 1e-06 
0.0 0.7959 0 -2.0 1e-06 
0.0 0.796 0 -2.0 1e-06 
0.0 0.7961 0 -2.0 1e-06 
0.0 0.7962 0 -2.0 1e-06 
0.0 0.7963 0 -2.0 1e-06 
0.0 0.7964 0 -2.0 1e-06 
0.0 0.7965 0 -2.0 1e-06 
0.0 0.7966 0 -2.0 1e-06 
0.0 0.7967 0 -2.0 1e-06 
0.0 0.7968 0 -2.0 1e-06 
0.0 0.7969 0 -2.0 1e-06 
0.0 0.797 0 -2.0 1e-06 
0.0 0.7971 0 -2.0 1e-06 
0.0 0.7972 0 -2.0 1e-06 
0.0 0.7973 0 -2.0 1e-06 
0.0 0.7974 0 -2.0 1e-06 
0.0 0.7975 0 -2.0 1e-06 
0.0 0.7976 0 -2.0 1e-06 
0.0 0.7977 0 -2.0 1e-06 
0.0 0.7978 0 -2.0 1e-06 
0.0 0.7979 0 -2.0 1e-06 
0.0 0.798 0 -2.0 1e-06 
0.0 0.7981 0 -2.0 1e-06 
0.0 0.7982 0 -2.0 1e-06 
0.0 0.7983 0 -2.0 1e-06 
0.0 0.7984 0 -2.0 1e-06 
0.0 0.7985 0 -2.0 1e-06 
0.0 0.7986 0 -2.0 1e-06 
0.0 0.7987 0 -2.0 1e-06 
0.0 0.7988 0 -2.0 1e-06 
0.0 0.7989 0 -2.0 1e-06 
0.0 0.799 0 -2.0 1e-06 
0.0 0.7991 0 -2.0 1e-06 
0.0 0.7992 0 -2.0 1e-06 
0.0 0.7993 0 -2.0 1e-06 
0.0 0.7994 0 -2.0 1e-06 
0.0 0.7995 0 -2.0 1e-06 
0.0 0.7996 0 -2.0 1e-06 
0.0 0.7997 0 -2.0 1e-06 
0.0 0.7998 0 -2.0 1e-06 
0.0 0.7999 0 -2.0 1e-06 
0.0 0.8 0 -2.0 1e-06 
0.0 0.8001 0 -2.0 1e-06 
0.0 0.8002 0 -2.0 1e-06 
0.0 0.8003 0 -2.0 1e-06 
0.0 0.8004 0 -2.0 1e-06 
0.0 0.8005 0 -2.0 1e-06 
0.0 0.8006 0 -2.0 1e-06 
0.0 0.8007 0 -2.0 1e-06 
0.0 0.8008 0 -2.0 1e-06 
0.0 0.8009 0 -2.0 1e-06 
0.0 0.801 0 -2.0 1e-06 
0.0 0.8011 0 -2.0 1e-06 
0.0 0.8012 0 -2.0 1e-06 
0.0 0.8013 0 -2.0 1e-06 
0.0 0.8014 0 -2.0 1e-06 
0.0 0.8015 0 -2.0 1e-06 
0.0 0.8016 0 -2.0 1e-06 
0.0 0.8017 0 -2.0 1e-06 
0.0 0.8018 0 -2.0 1e-06 
0.0 0.8019 0 -2.0 1e-06 
0.0 0.802 0 -2.0 1e-06 
0.0 0.8021 0 -2.0 1e-06 
0.0 0.8022 0 -2.0 1e-06 
0.0 0.8023 0 -2.0 1e-06 
0.0 0.8024 0 -2.0 1e-06 
0.0 0.8025 0 -2.0 1e-06 
0.0 0.8026 0 -2.0 1e-06 
0.0 0.8027 0 -2.0 1e-06 
0.0 0.8028 0 -2.0 1e-06 
0.0 0.8029 0 -2.0 1e-06 
0.0 0.803 0 -2.0 1e-06 
0.0 0.8031 0 -2.0 1e-06 
0.0 0.8032 0 -2.0 1e-06 
0.0 0.8033 0 -2.0 1e-06 
0.0 0.8034 0 -2.0 1e-06 
0.0 0.8035 0 -2.0 1e-06 
0.0 0.8036 0 -2.0 1e-06 
0.0 0.8037 0 -2.0 1e-06 
0.0 0.8038 0 -2.0 1e-06 
0.0 0.8039 0 -2.0 1e-06 
0.0 0.804 0 -2.0 1e-06 
0.0 0.8041 0 -2.0 1e-06 
0.0 0.8042 0 -2.0 1e-06 
0.0 0.8043 0 -2.0 1e-06 
0.0 0.8044 0 -2.0 1e-06 
0.0 0.8045 0 -2.0 1e-06 
0.0 0.8046 0 -2.0 1e-06 
0.0 0.8047 0 -2.0 1e-06 
0.0 0.8048 0 -2.0 1e-06 
0.0 0.8049 0 -2.0 1e-06 
0.0 0.805 0 -2.0 1e-06 
0.0 0.8051 0 -2.0 1e-06 
0.0 0.8052 0 -2.0 1e-06 
0.0 0.8053 0 -2.0 1e-06 
0.0 0.8054 0 -2.0 1e-06 
0.0 0.8055 0 -2.0 1e-06 
0.0 0.8056 0 -2.0 1e-06 
0.0 0.8057 0 -2.0 1e-06 
0.0 0.8058 0 -2.0 1e-06 
0.0 0.8059 0 -2.0 1e-06 
0.0 0.806 0 -2.0 1e-06 
0.0 0.8061 0 -2.0 1e-06 
0.0 0.8062 0 -2.0 1e-06 
0.0 0.8063 0 -2.0 1e-06 
0.0 0.8064 0 -2.0 1e-06 
0.0 0.8065 0 -2.0 1e-06 
0.0 0.8066 0 -2.0 1e-06 
0.0 0.8067 0 -2.0 1e-06 
0.0 0.8068 0 -2.0 1e-06 
0.0 0.8069 0 -2.0 1e-06 
0.0 0.807 0 -2.0 1e-06 
0.0 0.8071 0 -2.0 1e-06 
0.0 0.8072 0 -2.0 1e-06 
0.0 0.8073 0 -2.0 1e-06 
0.0 0.8074 0 -2.0 1e-06 
0.0 0.8075 0 -2.0 1e-06 
0.0 0.8076 0 -2.0 1e-06 
0.0 0.8077 0 -2.0 1e-06 
0.0 0.8078 0 -2.0 1e-06 
0.0 0.8079 0 -2.0 1e-06 
0.0 0.808 0 -2.0 1e-06 
0.0 0.8081 0 -2.0 1e-06 
0.0 0.8082 0 -2.0 1e-06 
0.0 0.8083 0 -2.0 1e-06 
0.0 0.8084 0 -2.0 1e-06 
0.0 0.8085 0 -2.0 1e-06 
0.0 0.8086 0 -2.0 1e-06 
0.0 0.8087 0 -2.0 1e-06 
0.0 0.8088 0 -2.0 1e-06 
0.0 0.8089 0 -2.0 1e-06 
0.0 0.809 0 -2.0 1e-06 
0.0 0.8091 0 -2.0 1e-06 
0.0 0.8092 0 -2.0 1e-06 
0.0 0.8093 0 -2.0 1e-06 
0.0 0.8094 0 -2.0 1e-06 
0.0 0.8095 0 -2.0 1e-06 
0.0 0.8096 0 -2.0 1e-06 
0.0 0.8097 0 -2.0 1e-06 
0.0 0.8098 0 -2.0 1e-06 
0.0 0.8099 0 -2.0 1e-06 
0.0 0.81 0 -2.0 1e-06 
0.0 0.8101 0 -2.0 1e-06 
0.0 0.8102 0 -2.0 1e-06 
0.0 0.8103 0 -2.0 1e-06 
0.0 0.8104 0 -2.0 1e-06 
0.0 0.8105 0 -2.0 1e-06 
0.0 0.8106 0 -2.0 1e-06 
0.0 0.8107 0 -2.0 1e-06 
0.0 0.8108 0 -2.0 1e-06 
0.0 0.8109 0 -2.0 1e-06 
0.0 0.811 0 -2.0 1e-06 
0.0 0.8111 0 -2.0 1e-06 
0.0 0.8112 0 -2.0 1e-06 
0.0 0.8113 0 -2.0 1e-06 
0.0 0.8114 0 -2.0 1e-06 
0.0 0.8115 0 -2.0 1e-06 
0.0 0.8116 0 -2.0 1e-06 
0.0 0.8117 0 -2.0 1e-06 
0.0 0.8118 0 -2.0 1e-06 
0.0 0.8119 0 -2.0 1e-06 
0.0 0.812 0 -2.0 1e-06 
0.0 0.8121 0 -2.0 1e-06 
0.0 0.8122 0 -2.0 1e-06 
0.0 0.8123 0 -2.0 1e-06 
0.0 0.8124 0 -2.0 1e-06 
0.0 0.8125 0 -2.0 1e-06 
0.0 0.8126 0 -2.0 1e-06 
0.0 0.8127 0 -2.0 1e-06 
0.0 0.8128 0 -2.0 1e-06 
0.0 0.8129 0 -2.0 1e-06 
0.0 0.813 0 -2.0 1e-06 
0.0 0.8131 0 -2.0 1e-06 
0.0 0.8132 0 -2.0 1e-06 
0.0 0.8133 0 -2.0 1e-06 
0.0 0.8134 0 -2.0 1e-06 
0.0 0.8135 0 -2.0 1e-06 
0.0 0.8136 0 -2.0 1e-06 
0.0 0.8137 0 -2.0 1e-06 
0.0 0.8138 0 -2.0 1e-06 
0.0 0.8139 0 -2.0 1e-06 
0.0 0.814 0 -2.0 1e-06 
0.0 0.8141 0 -2.0 1e-06 
0.0 0.8142 0 -2.0 1e-06 
0.0 0.8143 0 -2.0 1e-06 
0.0 0.8144 0 -2.0 1e-06 
0.0 0.8145 0 -2.0 1e-06 
0.0 0.8146 0 -2.0 1e-06 
0.0 0.8147 0 -2.0 1e-06 
0.0 0.8148 0 -2.0 1e-06 
0.0 0.8149 0 -2.0 1e-06 
0.0 0.815 0 -2.0 1e-06 
0.0 0.8151 0 -2.0 1e-06 
0.0 0.8152 0 -2.0 1e-06 
0.0 0.8153 0 -2.0 1e-06 
0.0 0.8154 0 -2.0 1e-06 
0.0 0.8155 0 -2.0 1e-06 
0.0 0.8156 0 -2.0 1e-06 
0.0 0.8157 0 -2.0 1e-06 
0.0 0.8158 0 -2.0 1e-06 
0.0 0.8159 0 -2.0 1e-06 
0.0 0.816 0 -2.0 1e-06 
0.0 0.8161 0 -2.0 1e-06 
0.0 0.8162 0 -2.0 1e-06 
0.0 0.8163 0 -2.0 1e-06 
0.0 0.8164 0 -2.0 1e-06 
0.0 0.8165 0 -2.0 1e-06 
0.0 0.8166 0 -2.0 1e-06 
0.0 0.8167 0 -2.0 1e-06 
0.0 0.8168 0 -2.0 1e-06 
0.0 0.8169 0 -2.0 1e-06 
0.0 0.817 0 -2.0 1e-06 
0.0 0.8171 0 -2.0 1e-06 
0.0 0.8172 0 -2.0 1e-06 
0.0 0.8173 0 -2.0 1e-06 
0.0 0.8174 0 -2.0 1e-06 
0.0 0.8175 0 -2.0 1e-06 
0.0 0.8176 0 -2.0 1e-06 
0.0 0.8177 0 -2.0 1e-06 
0.0 0.8178 0 -2.0 1e-06 
0.0 0.8179 0 -2.0 1e-06 
0.0 0.818 0 -2.0 1e-06 
0.0 0.8181 0 -2.0 1e-06 
0.0 0.8182 0 -2.0 1e-06 
0.0 0.8183 0 -2.0 1e-06 
0.0 0.8184 0 -2.0 1e-06 
0.0 0.8185 0 -2.0 1e-06 
0.0 0.8186 0 -2.0 1e-06 
0.0 0.8187 0 -2.0 1e-06 
0.0 0.8188 0 -2.0 1e-06 
0.0 0.8189 0 -2.0 1e-06 
0.0 0.819 0 -2.0 1e-06 
0.0 0.8191 0 -2.0 1e-06 
0.0 0.8192 0 -2.0 1e-06 
0.0 0.8193 0 -2.0 1e-06 
0.0 0.8194 0 -2.0 1e-06 
0.0 0.8195 0 -2.0 1e-06 
0.0 0.8196 0 -2.0 1e-06 
0.0 0.8197 0 -2.0 1e-06 
0.0 0.8198 0 -2.0 1e-06 
0.0 0.8199 0 -2.0 1e-06 
0.0 0.82 0 -2.0 1e-06 
0.0 0.8201 0 -2.0 1e-06 
0.0 0.8202 0 -2.0 1e-06 
0.0 0.8203 0 -2.0 1e-06 
0.0 0.8204 0 -2.0 1e-06 
0.0 0.8205 0 -2.0 1e-06 
0.0 0.8206 0 -2.0 1e-06 
0.0 0.8207 0 -2.0 1e-06 
0.0 0.8208 0 -2.0 1e-06 
0.0 0.8209 0 -2.0 1e-06 
0.0 0.821 0 -2.0 1e-06 
0.0 0.8211 0 -2.0 1e-06 
0.0 0.8212 0 -2.0 1e-06 
0.0 0.8213 0 -2.0 1e-06 
0.0 0.8214 0 -2.0 1e-06 
0.0 0.8215 0 -2.0 1e-06 
0.0 0.8216 0 -2.0 1e-06 
0.0 0.8217 0 -2.0 1e-06 
0.0 0.8218 0 -2.0 1e-06 
0.0 0.8219 0 -2.0 1e-06 
0.0 0.822 0 -2.0 1e-06 
0.0 0.8221 0 -2.0 1e-06 
0.0 0.8222 0 -2.0 1e-06 
0.0 0.8223 0 -2.0 1e-06 
0.0 0.8224 0 -2.0 1e-06 
0.0 0.8225 0 -2.0 1e-06 
0.0 0.8226 0 -2.0 1e-06 
0.0 0.8227 0 -2.0 1e-06 
0.0 0.8228 0 -2.0 1e-06 
0.0 0.8229 0 -2.0 1e-06 
0.0 0.823 0 -2.0 1e-06 
0.0 0.8231 0 -2.0 1e-06 
0.0 0.8232 0 -2.0 1e-06 
0.0 0.8233 0 -2.0 1e-06 
0.0 0.8234 0 -2.0 1e-06 
0.0 0.8235 0 -2.0 1e-06 
0.0 0.8236 0 -2.0 1e-06 
0.0 0.8237 0 -2.0 1e-06 
0.0 0.8238 0 -2.0 1e-06 
0.0 0.8239 0 -2.0 1e-06 
0.0 0.824 0 -2.0 1e-06 
0.0 0.8241 0 -2.0 1e-06 
0.0 0.8242 0 -2.0 1e-06 
0.0 0.8243 0 -2.0 1e-06 
0.0 0.8244 0 -2.0 1e-06 
0.0 0.8245 0 -2.0 1e-06 
0.0 0.8246 0 -2.0 1e-06 
0.0 0.8247 0 -2.0 1e-06 
0.0 0.8248 0 -2.0 1e-06 
0.0 0.8249 0 -2.0 1e-06 
0.0 0.825 0 -2.0 1e-06 
0.0 0.8251 0 -2.0 1e-06 
0.0 0.8252 0 -2.0 1e-06 
0.0 0.8253 0 -2.0 1e-06 
0.0 0.8254 0 -2.0 1e-06 
0.0 0.8255 0 -2.0 1e-06 
0.0 0.8256 0 -2.0 1e-06 
0.0 0.8257 0 -2.0 1e-06 
0.0 0.8258 0 -2.0 1e-06 
0.0 0.8259 0 -2.0 1e-06 
0.0 0.826 0 -2.0 1e-06 
0.0 0.8261 0 -2.0 1e-06 
0.0 0.8262 0 -2.0 1e-06 
0.0 0.8263 0 -2.0 1e-06 
0.0 0.8264 0 -2.0 1e-06 
0.0 0.8265 0 -2.0 1e-06 
0.0 0.8266 0 -2.0 1e-06 
0.0 0.8267 0 -2.0 1e-06 
0.0 0.8268 0 -2.0 1e-06 
0.0 0.8269 0 -2.0 1e-06 
0.0 0.827 0 -2.0 1e-06 
0.0 0.8271 0 -2.0 1e-06 
0.0 0.8272 0 -2.0 1e-06 
0.0 0.8273 0 -2.0 1e-06 
0.0 0.8274 0 -2.0 1e-06 
0.0 0.8275 0 -2.0 1e-06 
0.0 0.8276 0 -2.0 1e-06 
0.0 0.8277 0 -2.0 1e-06 
0.0 0.8278 0 -2.0 1e-06 
0.0 0.8279 0 -2.0 1e-06 
0.0 0.828 0 -2.0 1e-06 
0.0 0.8281 0 -2.0 1e-06 
0.0 0.8282 0 -2.0 1e-06 
0.0 0.8283 0 -2.0 1e-06 
0.0 0.8284 0 -2.0 1e-06 
0.0 0.8285 0 -2.0 1e-06 
0.0 0.8286 0 -2.0 1e-06 
0.0 0.8287 0 -2.0 1e-06 
0.0 0.8288 0 -2.0 1e-06 
0.0 0.8289 0 -2.0 1e-06 
0.0 0.829 0 -2.0 1e-06 
0.0 0.8291 0 -2.0 1e-06 
0.0 0.8292 0 -2.0 1e-06 
0.0 0.8293 0 -2.0 1e-06 
0.0 0.8294 0 -2.0 1e-06 
0.0 0.8295 0 -2.0 1e-06 
0.0 0.8296 0 -2.0 1e-06 
0.0 0.8297 0 -2.0 1e-06 
0.0 0.8298 0 -2.0 1e-06 
0.0 0.8299 0 -2.0 1e-06 
0.0 0.83 0 -2.0 1e-06 
0.0 0.8301 0 -2.0 1e-06 
0.0 0.8302 0 -2.0 1e-06 
0.0 0.8303 0 -2.0 1e-06 
0.0 0.8304 0 -2.0 1e-06 
0.0 0.8305 0 -2.0 1e-06 
0.0 0.8306 0 -2.0 1e-06 
0.0 0.8307 0 -2.0 1e-06 
0.0 0.8308 0 -2.0 1e-06 
0.0 0.8309 0 -2.0 1e-06 
0.0 0.831 0 -2.0 1e-06 
0.0 0.8311 0 -2.0 1e-06 
0.0 0.8312 0 -2.0 1e-06 
0.0 0.8313 0 -2.0 1e-06 
0.0 0.8314 0 -2.0 1e-06 
0.0 0.8315 0 -2.0 1e-06 
0.0 0.8316 0 -2.0 1e-06 
0.0 0.8317 0 -2.0 1e-06 
0.0 0.8318 0 -2.0 1e-06 
0.0 0.8319 0 -2.0 1e-06 
0.0 0.832 0 -2.0 1e-06 
0.0 0.8321 0 -2.0 1e-06 
0.0 0.8322 0 -2.0 1e-06 
0.0 0.8323 0 -2.0 1e-06 
0.0 0.8324 0 -2.0 1e-06 
0.0 0.8325 0 -2.0 1e-06 
0.0 0.8326 0 -2.0 1e-06 
0.0 0.8327 0 -2.0 1e-06 
0.0 0.8328 0 -2.0 1e-06 
0.0 0.8329 0 -2.0 1e-06 
0.0 0.833 0 -2.0 1e-06 
0.0 0.8331 0 -2.0 1e-06 
0.0 0.8332 0 -2.0 1e-06 
0.0 0.8333 0 -2.0 1e-06 
0.0 0.8334 0 -2.0 1e-06 
0.0 0.8335 0 -2.0 1e-06 
0.0 0.8336 0 -2.0 1e-06 
0.0 0.8337 0 -2.0 1e-06 
0.0 0.8338 0 -2.0 1e-06 
0.0 0.8339 0 -2.0 1e-06 
0.0 0.834 0 -2.0 1e-06 
0.0 0.8341 0 -2.0 1e-06 
0.0 0.8342 0 -2.0 1e-06 
0.0 0.8343 0 -2.0 1e-06 
0.0 0.8344 0 -2.0 1e-06 
0.0 0.8345 0 -2.0 1e-06 
0.0 0.8346 0 -2.0 1e-06 
0.0 0.8347 0 -2.0 1e-06 
0.0 0.8348 0 -2.0 1e-06 
0.0 0.8349 0 -2.0 1e-06 
0.0 0.835 0 -2.0 1e-06 
0.0 0.8351 0 -2.0 1e-06 
0.0 0.8352 0 -2.0 1e-06 
0.0 0.8353 0 -2.0 1e-06 
0.0 0.8354 0 -2.0 1e-06 
0.0 0.8355 0 -2.0 1e-06 
0.0 0.8356 0 -2.0 1e-06 
0.0 0.8357 0 -2.0 1e-06 
0.0 0.8358 0 -2.0 1e-06 
0.0 0.8359 0 -2.0 1e-06 
0.0 0.836 0 -2.0 1e-06 
0.0 0.8361 0 -2.0 1e-06 
0.0 0.8362 0 -2.0 1e-06 
0.0 0.8363 0 -2.0 1e-06 
0.0 0.8364 0 -2.0 1e-06 
0.0 0.8365 0 -2.0 1e-06 
0.0 0.8366 0 -2.0 1e-06 
0.0 0.8367 0 -2.0 1e-06 
0.0 0.8368 0 -2.0 1e-06 
0.0 0.8369 0 -2.0 1e-06 
0.0 0.837 0 -2.0 1e-06 
0.0 0.8371 0 -2.0 1e-06 
0.0 0.8372 0 -2.0 1e-06 
0.0 0.8373 0 -2.0 1e-06 
0.0 0.8374 0 -2.0 1e-06 
0.0 0.8375 0 -2.0 1e-06 
0.0 0.8376 0 -2.0 1e-06 
0.0 0.8377 0 -2.0 1e-06 
0.0 0.8378 0 -2.0 1e-06 
0.0 0.8379 0 -2.0 1e-06 
0.0 0.838 0 -2.0 1e-06 
0.0 0.8381 0 -2.0 1e-06 
0.0 0.8382 0 -2.0 1e-06 
0.0 0.8383 0 -2.0 1e-06 
0.0 0.8384 0 -2.0 1e-06 
0.0 0.8385 0 -2.0 1e-06 
0.0 0.8386 0 -2.0 1e-06 
0.0 0.8387 0 -2.0 1e-06 
0.0 0.8388 0 -2.0 1e-06 
0.0 0.8389 0 -2.0 1e-06 
0.0 0.839 0 -2.0 1e-06 
0.0 0.8391 0 -2.0 1e-06 
0.0 0.8392 0 -2.0 1e-06 
0.0 0.8393 0 -2.0 1e-06 
0.0 0.8394 0 -2.0 1e-06 
0.0 0.8395 0 -2.0 1e-06 
0.0 0.8396 0 -2.0 1e-06 
0.0 0.8397 0 -2.0 1e-06 
0.0 0.8398 0 -2.0 1e-06 
0.0 0.8399 0 -2.0 1e-06 
0.0 0.84 0 -2.0 1e-06 
0.0 0.8401 0 -2.0 1e-06 
0.0 0.8402 0 -2.0 1e-06 
0.0 0.8403 0 -2.0 1e-06 
0.0 0.8404 0 -2.0 1e-06 
0.0 0.8405 0 -2.0 1e-06 
0.0 0.8406 0 -2.0 1e-06 
0.0 0.8407 0 -2.0 1e-06 
0.0 0.8408 0 -2.0 1e-06 
0.0 0.8409 0 -2.0 1e-06 
0.0 0.841 0 -2.0 1e-06 
0.0 0.8411 0 -2.0 1e-06 
0.0 0.8412 0 -2.0 1e-06 
0.0 0.8413 0 -2.0 1e-06 
0.0 0.8414 0 -2.0 1e-06 
0.0 0.8415 0 -2.0 1e-06 
0.0 0.8416 0 -2.0 1e-06 
0.0 0.8417 0 -2.0 1e-06 
0.0 0.8418 0 -2.0 1e-06 
0.0 0.8419 0 -2.0 1e-06 
0.0 0.842 0 -2.0 1e-06 
0.0 0.8421 0 -2.0 1e-06 
0.0 0.8422 0 -2.0 1e-06 
0.0 0.8423 0 -2.0 1e-06 
0.0 0.8424 0 -2.0 1e-06 
0.0 0.8425 0 -2.0 1e-06 
0.0 0.8426 0 -2.0 1e-06 
0.0 0.8427 0 -2.0 1e-06 
0.0 0.8428 0 -2.0 1e-06 
0.0 0.8429 0 -2.0 1e-06 
0.0 0.843 0 -2.0 1e-06 
0.0 0.8431 0 -2.0 1e-06 
0.0 0.8432 0 -2.0 1e-06 
0.0 0.8433 0 -2.0 1e-06 
0.0 0.8434 0 -2.0 1e-06 
0.0 0.8435 0 -2.0 1e-06 
0.0 0.8436 0 -2.0 1e-06 
0.0 0.8437 0 -2.0 1e-06 
0.0 0.8438 0 -2.0 1e-06 
0.0 0.8439 0 -2.0 1e-06 
0.0 0.844 0 -2.0 1e-06 
0.0 0.8441 0 -2.0 1e-06 
0.0 0.8442 0 -2.0 1e-06 
0.0 0.8443 0 -2.0 1e-06 
0.0 0.8444 0 -2.0 1e-06 
0.0 0.8445 0 -2.0 1e-06 
0.0 0.8446 0 -2.0 1e-06 
0.0 0.8447 0 -2.0 1e-06 
0.0 0.8448 0 -2.0 1e-06 
0.0 0.8449 0 -2.0 1e-06 
0.0 0.845 0 -2.0 1e-06 
0.0 0.8451 0 -2.0 1e-06 
0.0 0.8452 0 -2.0 1e-06 
0.0 0.8453 0 -2.0 1e-06 
0.0 0.8454 0 -2.0 1e-06 
0.0 0.8455 0 -2.0 1e-06 
0.0 0.8456 0 -2.0 1e-06 
0.0 0.8457 0 -2.0 1e-06 
0.0 0.8458 0 -2.0 1e-06 
0.0 0.8459 0 -2.0 1e-06 
0.0 0.846 0 -2.0 1e-06 
0.0 0.8461 0 -2.0 1e-06 
0.0 0.8462 0 -2.0 1e-06 
0.0 0.8463 0 -2.0 1e-06 
0.0 0.8464 0 -2.0 1e-06 
0.0 0.8465 0 -2.0 1e-06 
0.0 0.8466 0 -2.0 1e-06 
0.0 0.8467 0 -2.0 1e-06 
0.0 0.8468 0 -2.0 1e-06 
0.0 0.8469 0 -2.0 1e-06 
0.0 0.847 0 -2.0 1e-06 
0.0 0.8471 0 -2.0 1e-06 
0.0 0.8472 0 -2.0 1e-06 
0.0 0.8473 0 -2.0 1e-06 
0.0 0.8474 0 -2.0 1e-06 
0.0 0.8475 0 -2.0 1e-06 
0.0 0.8476 0 -2.0 1e-06 
0.0 0.8477 0 -2.0 1e-06 
0.0 0.8478 0 -2.0 1e-06 
0.0 0.8479 0 -2.0 1e-06 
0.0 0.848 0 -2.0 1e-06 
0.0 0.8481 0 -2.0 1e-06 
0.0 0.8482 0 -2.0 1e-06 
0.0 0.8483 0 -2.0 1e-06 
0.0 0.8484 0 -2.0 1e-06 
0.0 0.8485 0 -2.0 1e-06 
0.0 0.8486 0 -2.0 1e-06 
0.0 0.8487 0 -2.0 1e-06 
0.0 0.8488 0 -2.0 1e-06 
0.0 0.8489 0 -2.0 1e-06 
0.0 0.849 0 -2.0 1e-06 
0.0 0.8491 0 -2.0 1e-06 
0.0 0.8492 0 -2.0 1e-06 
0.0 0.8493 0 -2.0 1e-06 
0.0 0.8494 0 -2.0 1e-06 
0.0 0.8495 0 -2.0 1e-06 
0.0 0.8496 0 -2.0 1e-06 
0.0 0.8497 0 -2.0 1e-06 
0.0 0.8498 0 -2.0 1e-06 
0.0 0.8499 0 -2.0 1e-06 
0.0 0.85 0 -2.0 1e-06 
0.0 0.8501 0 -2.0 1e-06 
0.0 0.8502 0 -2.0 1e-06 
0.0 0.8503 0 -2.0 1e-06 
0.0 0.8504 0 -2.0 1e-06 
0.0 0.8505 0 -2.0 1e-06 
0.0 0.8506 0 -2.0 1e-06 
0.0 0.8507 0 -2.0 1e-06 
0.0 0.8508 0 -2.0 1e-06 
0.0 0.8509 0 -2.0 1e-06 
0.0 0.851 0 -2.0 1e-06 
0.0 0.8511 0 -2.0 1e-06 
0.0 0.8512 0 -2.0 1e-06 
0.0 0.8513 0 -2.0 1e-06 
0.0 0.8514 0 -2.0 1e-06 
0.0 0.8515 0 -2.0 1e-06 
0.0 0.8516 0 -2.0 1e-06 
0.0 0.8517 0 -2.0 1e-06 
0.0 0.8518 0 -2.0 1e-06 
0.0 0.8519 0 -2.0 1e-06 
0.0 0.852 0 -2.0 1e-06 
0.0 0.8521 0 -2.0 1e-06 
0.0 0.8522 0 -2.0 1e-06 
0.0 0.8523 0 -2.0 1e-06 
0.0 0.8524 0 -2.0 1e-06 
0.0 0.8525 0 -2.0 1e-06 
0.0 0.8526 0 -2.0 1e-06 
0.0 0.8527 0 -2.0 1e-06 
0.0 0.8528 0 -2.0 1e-06 
0.0 0.8529 0 -2.0 1e-06 
0.0 0.853 0 -2.0 1e-06 
0.0 0.8531 0 -2.0 1e-06 
0.0 0.8532 0 -2.0 1e-06 
0.0 0.8533 0 -2.0 1e-06 
0.0 0.8534 0 -2.0 1e-06 
0.0 0.8535 0 -2.0 1e-06 
0.0 0.8536 0 -2.0 1e-06 
0.0 0.8537 0 -2.0 1e-06 
0.0 0.8538 0 -2.0 1e-06 
0.0 0.8539 0 -2.0 1e-06 
0.0 0.854 0 -2.0 1e-06 
0.0 0.8541 0 -2.0 1e-06 
0.0 0.8542 0 -2.0 1e-06 
0.0 0.8543 0 -2.0 1e-06 
0.0 0.8544 0 -2.0 1e-06 
0.0 0.8545 0 -2.0 1e-06 
0.0 0.8546 0 -2.0 1e-06 
0.0 0.8547 0 -2.0 1e-06 
0.0 0.8548 0 -2.0 1e-06 
0.0 0.8549 0 -2.0 1e-06 
0.0 0.855 0 -2.0 1e-06 
0.0 0.8551 0 -2.0 1e-06 
0.0 0.8552 0 -2.0 1e-06 
0.0 0.8553 0 -2.0 1e-06 
0.0 0.8554 0 -2.0 1e-06 
0.0 0.8555 0 -2.0 1e-06 
0.0 0.8556 0 -2.0 1e-06 
0.0 0.8557 0 -2.0 1e-06 
0.0 0.8558 0 -2.0 1e-06 
0.0 0.8559 0 -2.0 1e-06 
0.0 0.856 0 -2.0 1e-06 
0.0 0.8561 0 -2.0 1e-06 
0.0 0.8562 0 -2.0 1e-06 
0.0 0.8563 0 -2.0 1e-06 
0.0 0.8564 0 -2.0 1e-06 
0.0 0.8565 0 -2.0 1e-06 
0.0 0.8566 0 -2.0 1e-06 
0.0 0.8567 0 -2.0 1e-06 
0.0 0.8568 0 -2.0 1e-06 
0.0 0.8569 0 -2.0 1e-06 
0.0 0.857 0 -2.0 1e-06 
0.0 0.8571 0 -2.0 1e-06 
0.0 0.8572 0 -2.0 1e-06 
0.0 0.8573 0 -2.0 1e-06 
0.0 0.8574 0 -2.0 1e-06 
0.0 0.8575 0 -2.0 1e-06 
0.0 0.8576 0 -2.0 1e-06 
0.0 0.8577 0 -2.0 1e-06 
0.0 0.8578 0 -2.0 1e-06 
0.0 0.8579 0 -2.0 1e-06 
0.0 0.858 0 -2.0 1e-06 
0.0 0.8581 0 -2.0 1e-06 
0.0 0.8582 0 -2.0 1e-06 
0.0 0.8583 0 -2.0 1e-06 
0.0 0.8584 0 -2.0 1e-06 
0.0 0.8585 0 -2.0 1e-06 
0.0 0.8586 0 -2.0 1e-06 
0.0 0.8587 0 -2.0 1e-06 
0.0 0.8588 0 -2.0 1e-06 
0.0 0.8589 0 -2.0 1e-06 
0.0 0.859 0 -2.0 1e-06 
0.0 0.8591 0 -2.0 1e-06 
0.0 0.8592 0 -2.0 1e-06 
0.0 0.8593 0 -2.0 1e-06 
0.0 0.8594 0 -2.0 1e-06 
0.0 0.8595 0 -2.0 1e-06 
0.0 0.8596 0 -2.0 1e-06 
0.0 0.8597 0 -2.0 1e-06 
0.0 0.8598 0 -2.0 1e-06 
0.0 0.8599 0 -2.0 1e-06 
0.0 0.86 0 -2.0 1e-06 
0.0 0.8601 0 -2.0 1e-06 
0.0 0.8602 0 -2.0 1e-06 
0.0 0.8603 0 -2.0 1e-06 
0.0 0.8604 0 -2.0 1e-06 
0.0 0.8605 0 -2.0 1e-06 
0.0 0.8606 0 -2.0 1e-06 
0.0 0.8607 0 -2.0 1e-06 
0.0 0.8608 0 -2.0 1e-06 
0.0 0.8609 0 -2.0 1e-06 
0.0 0.861 0 -2.0 1e-06 
0.0 0.8611 0 -2.0 1e-06 
0.0 0.8612 0 -2.0 1e-06 
0.0 0.8613 0 -2.0 1e-06 
0.0 0.8614 0 -2.0 1e-06 
0.0 0.8615 0 -2.0 1e-06 
0.0 0.8616 0 -2.0 1e-06 
0.0 0.8617 0 -2.0 1e-06 
0.0 0.8618 0 -2.0 1e-06 
0.0 0.8619 0 -2.0 1e-06 
0.0 0.862 0 -2.0 1e-06 
0.0 0.8621 0 -2.0 1e-06 
0.0 0.8622 0 -2.0 1e-06 
0.0 0.8623 0 -2.0 1e-06 
0.0 0.8624 0 -2.0 1e-06 
0.0 0.8625 0 -2.0 1e-06 
0.0 0.8626 0 -2.0 1e-06 
0.0 0.8627 0 -2.0 1e-06 
0.0 0.8628 0 -2.0 1e-06 
0.0 0.8629 0 -2.0 1e-06 
0.0 0.863 0 -2.0 1e-06 
0.0 0.8631 0 -2.0 1e-06 
0.0 0.8632 0 -2.0 1e-06 
0.0 0.8633 0 -2.0 1e-06 
0.0 0.8634 0 -2.0 1e-06 
0.0 0.8635 0 -2.0 1e-06 
0.0 0.8636 0 -2.0 1e-06 
0.0 0.8637 0 -2.0 1e-06 
0.0 0.8638 0 -2.0 1e-06 
0.0 0.8639 0 -2.0 1e-06 
0.0 0.864 0 -2.0 1e-06 
0.0 0.8641 0 -2.0 1e-06 
0.0 0.8642 0 -2.0 1e-06 
0.0 0.8643 0 -2.0 1e-06 
0.0 0.8644 0 -2.0 1e-06 
0.0 0.8645 0 -2.0 1e-06 
0.0 0.8646 0 -2.0 1e-06 
0.0 0.8647 0 -2.0 1e-06 
0.0 0.8648 0 -2.0 1e-06 
0.0 0.8649 0 -2.0 1e-06 
0.0 0.865 0 -2.0 1e-06 
0.0 0.8651 0 -2.0 1e-06 
0.0 0.8652 0 -2.0 1e-06 
0.0 0.8653 0 -2.0 1e-06 
0.0 0.8654 0 -2.0 1e-06 
0.0 0.8655 0 -2.0 1e-06 
0.0 0.8656 0 -2.0 1e-06 
0.0 0.8657 0 -2.0 1e-06 
0.0 0.8658 0 -2.0 1e-06 
0.0 0.8659 0 -2.0 1e-06 
0.0 0.866 0 -2.0 1e-06 
0.0 0.8661 0 -2.0 1e-06 
0.0 0.8662 0 -2.0 1e-06 
0.0 0.8663 0 -2.0 1e-06 
0.0 0.8664 0 -2.0 1e-06 
0.0 0.8665 0 -2.0 1e-06 
0.0 0.8666 0 -2.0 1e-06 
0.0 0.8667 0 -2.0 1e-06 
0.0 0.8668 0 -2.0 1e-06 
0.0 0.8669 0 -2.0 1e-06 
0.0 0.867 0 -2.0 1e-06 
0.0 0.8671 0 -2.0 1e-06 
0.0 0.8672 0 -2.0 1e-06 
0.0 0.8673 0 -2.0 1e-06 
0.0 0.8674 0 -2.0 1e-06 
0.0 0.8675 0 -2.0 1e-06 
0.0 0.8676 0 -2.0 1e-06 
0.0 0.8677 0 -2.0 1e-06 
0.0 0.8678 0 -2.0 1e-06 
0.0 0.8679 0 -2.0 1e-06 
0.0 0.868 0 -2.0 1e-06 
0.0 0.8681 0 -2.0 1e-06 
0.0 0.8682 0 -2.0 1e-06 
0.0 0.8683 0 -2.0 1e-06 
0.0 0.8684 0 -2.0 1e-06 
0.0 0.8685 0 -2.0 1e-06 
0.0 0.8686 0 -2.0 1e-06 
0.0 0.8687 0 -2.0 1e-06 
0.0 0.8688 0 -2.0 1e-06 
0.0 0.8689 0 -2.0 1e-06 
0.0 0.869 0 -2.0 1e-06 
0.0 0.8691 0 -2.0 1e-06 
0.0 0.8692 0 -2.0 1e-06 
0.0 0.8693 0 -2.0 1e-06 
0.0 0.8694 0 -2.0 1e-06 
0.0 0.8695 0 -2.0 1e-06 
0.0 0.8696 0 -2.0 1e-06 
0.0 0.8697 0 -2.0 1e-06 
0.0 0.8698 0 -2.0 1e-06 
0.0 0.8699 0 -2.0 1e-06 
0.0 0.87 0 -2.0 1e-06 
0.0 0.8701 0 -2.0 1e-06 
0.0 0.8702 0 -2.0 1e-06 
0.0 0.8703 0 -2.0 1e-06 
0.0 0.8704 0 -2.0 1e-06 
0.0 0.8705 0 -2.0 1e-06 
0.0 0.8706 0 -2.0 1e-06 
0.0 0.8707 0 -2.0 1e-06 
0.0 0.8708 0 -2.0 1e-06 
0.0 0.8709 0 -2.0 1e-06 
0.0 0.871 0 -2.0 1e-06 
0.0 0.8711 0 -2.0 1e-06 
0.0 0.8712 0 -2.0 1e-06 
0.0 0.8713 0 -2.0 1e-06 
0.0 0.8714 0 -2.0 1e-06 
0.0 0.8715 0 -2.0 1e-06 
0.0 0.8716 0 -2.0 1e-06 
0.0 0.8717 0 -2.0 1e-06 
0.0 0.8718 0 -2.0 1e-06 
0.0 0.8719 0 -2.0 1e-06 
0.0 0.872 0 -2.0 1e-06 
0.0 0.8721 0 -2.0 1e-06 
0.0 0.8722 0 -2.0 1e-06 
0.0 0.8723 0 -2.0 1e-06 
0.0 0.8724 0 -2.0 1e-06 
0.0 0.8725 0 -2.0 1e-06 
0.0 0.8726 0 -2.0 1e-06 
0.0 0.8727 0 -2.0 1e-06 
0.0 0.8728 0 -2.0 1e-06 
0.0 0.8729 0 -2.0 1e-06 
0.0 0.873 0 -2.0 1e-06 
0.0 0.8731 0 -2.0 1e-06 
0.0 0.8732 0 -2.0 1e-06 
0.0 0.8733 0 -2.0 1e-06 
0.0 0.8734 0 -2.0 1e-06 
0.0 0.8735 0 -2.0 1e-06 
0.0 0.8736 0 -2.0 1e-06 
0.0 0.8737 0 -2.0 1e-06 
0.0 0.8738 0 -2.0 1e-06 
0.0 0.8739 0 -2.0 1e-06 
0.0 0.874 0 -2.0 1e-06 
0.0 0.8741 0 -2.0 1e-06 
0.0 0.8742 0 -2.0 1e-06 
0.0 0.8743 0 -2.0 1e-06 
0.0 0.8744 0 -2.0 1e-06 
0.0 0.8745 0 -2.0 1e-06 
0.0 0.8746 0 -2.0 1e-06 
0.0 0.8747 0 -2.0 1e-06 
0.0 0.8748 0 -2.0 1e-06 
0.0 0.8749 0 -2.0 1e-06 
0.0 0.875 0 -2.0 1e-06 
0.0 0.8751 0 -2.0 1e-06 
0.0 0.8752 0 -2.0 1e-06 
0.0 0.8753 0 -2.0 1e-06 
0.0 0.8754 0 -2.0 1e-06 
0.0 0.8755 0 -2.0 1e-06 
0.0 0.8756 0 -2.0 1e-06 
0.0 0.8757 0 -2.0 1e-06 
0.0 0.8758 0 -2.0 1e-06 
0.0 0.8759 0 -2.0 1e-06 
0.0 0.876 0 -2.0 1e-06 
0.0 0.8761 0 -2.0 1e-06 
0.0 0.8762 0 -2.0 1e-06 
0.0 0.8763 0 -2.0 1e-06 
0.0 0.8764 0 -2.0 1e-06 
0.0 0.8765 0 -2.0 1e-06 
0.0 0.8766 0 -2.0 1e-06 
0.0 0.8767 0 -2.0 1e-06 
0.0 0.8768 0 -2.0 1e-06 
0.0 0.8769 0 -2.0 1e-06 
0.0 0.877 0 -2.0 1e-06 
0.0 0.8771 0 -2.0 1e-06 
0.0 0.8772 0 -2.0 1e-06 
0.0 0.8773 0 -2.0 1e-06 
0.0 0.8774 0 -2.0 1e-06 
0.0 0.8775 0 -2.0 1e-06 
0.0 0.8776 0 -2.0 1e-06 
0.0 0.8777 0 -2.0 1e-06 
0.0 0.8778 0 -2.0 1e-06 
0.0 0.8779 0 -2.0 1e-06 
0.0 0.878 0 -2.0 1e-06 
0.0 0.8781 0 -2.0 1e-06 
0.0 0.8782 0 -2.0 1e-06 
0.0 0.8783 0 -2.0 1e-06 
0.0 0.8784 0 -2.0 1e-06 
0.0 0.8785 0 -2.0 1e-06 
0.0 0.8786 0 -2.0 1e-06 
0.0 0.8787 0 -2.0 1e-06 
0.0 0.8788 0 -2.0 1e-06 
0.0 0.8789 0 -2.0 1e-06 
0.0 0.879 0 -2.0 1e-06 
0.0 0.8791 0 -2.0 1e-06 
0.0 0.8792 0 -2.0 1e-06 
0.0 0.8793 0 -2.0 1e-06 
0.0 0.8794 0 -2.0 1e-06 
0.0 0.8795 0 -2.0 1e-06 
0.0 0.8796 0 -2.0 1e-06 
0.0 0.8797 0 -2.0 1e-06 
0.0 0.8798 0 -2.0 1e-06 
0.0 0.8799 0 -2.0 1e-06 
0.0 0.88 0 -2.0 1e-06 
0.0 0.8801 0 -2.0 1e-06 
0.0 0.8802 0 -2.0 1e-06 
0.0 0.8803 0 -2.0 1e-06 
0.0 0.8804 0 -2.0 1e-06 
0.0 0.8805 0 -2.0 1e-06 
0.0 0.8806 0 -2.0 1e-06 
0.0 0.8807 0 -2.0 1e-06 
0.0 0.8808 0 -2.0 1e-06 
0.0 0.8809 0 -2.0 1e-06 
0.0 0.881 0 -2.0 1e-06 
0.0 0.8811 0 -2.0 1e-06 
0.0 0.8812 0 -2.0 1e-06 
0.0 0.8813 0 -2.0 1e-06 
0.0 0.8814 0 -2.0 1e-06 
0.0 0.8815 0 -2.0 1e-06 
0.0 0.8816 0 -2.0 1e-06 
0.0 0.8817 0 -2.0 1e-06 
0.0 0.8818 0 -2.0 1e-06 
0.0 0.8819 0 -2.0 1e-06 
0.0 0.882 0 -2.0 1e-06 
0.0 0.8821 0 -2.0 1e-06 
0.0 0.8822 0 -2.0 1e-06 
0.0 0.8823 0 -2.0 1e-06 
0.0 0.8824 0 -2.0 1e-06 
0.0 0.8825 0 -2.0 1e-06 
0.0 0.8826 0 -2.0 1e-06 
0.0 0.8827 0 -2.0 1e-06 
0.0 0.8828 0 -2.0 1e-06 
0.0 0.8829 0 -2.0 1e-06 
0.0 0.883 0 -2.0 1e-06 
0.0 0.8831 0 -2.0 1e-06 
0.0 0.8832 0 -2.0 1e-06 
0.0 0.8833 0 -2.0 1e-06 
0.0 0.8834 0 -2.0 1e-06 
0.0 0.8835 0 -2.0 1e-06 
0.0 0.8836 0 -2.0 1e-06 
0.0 0.8837 0 -2.0 1e-06 
0.0 0.8838 0 -2.0 1e-06 
0.0 0.8839 0 -2.0 1e-06 
0.0 0.884 0 -2.0 1e-06 
0.0 0.8841 0 -2.0 1e-06 
0.0 0.8842 0 -2.0 1e-06 
0.0 0.8843 0 -2.0 1e-06 
0.0 0.8844 0 -2.0 1e-06 
0.0 0.8845 0 -2.0 1e-06 
0.0 0.8846 0 -2.0 1e-06 
0.0 0.8847 0 -2.0 1e-06 
0.0 0.8848 0 -2.0 1e-06 
0.0 0.8849 0 -2.0 1e-06 
0.0 0.885 0 -2.0 1e-06 
0.0 0.8851 0 -2.0 1e-06 
0.0 0.8852 0 -2.0 1e-06 
0.0 0.8853 0 -2.0 1e-06 
0.0 0.8854 0 -2.0 1e-06 
0.0 0.8855 0 -2.0 1e-06 
0.0 0.8856 0 -2.0 1e-06 
0.0 0.8857 0 -2.0 1e-06 
0.0 0.8858 0 -2.0 1e-06 
0.0 0.8859 0 -2.0 1e-06 
0.0 0.886 0 -2.0 1e-06 
0.0 0.8861 0 -2.0 1e-06 
0.0 0.8862 0 -2.0 1e-06 
0.0 0.8863 0 -2.0 1e-06 
0.0 0.8864 0 -2.0 1e-06 
0.0 0.8865 0 -2.0 1e-06 
0.0 0.8866 0 -2.0 1e-06 
0.0 0.8867 0 -2.0 1e-06 
0.0 0.8868 0 -2.0 1e-06 
0.0 0.8869 0 -2.0 1e-06 
0.0 0.887 0 -2.0 1e-06 
0.0 0.8871 0 -2.0 1e-06 
0.0 0.8872 0 -2.0 1e-06 
0.0 0.8873 0 -2.0 1e-06 
0.0 0.8874 0 -2.0 1e-06 
0.0 0.8875 0 -2.0 1e-06 
0.0 0.8876 0 -2.0 1e-06 
0.0 0.8877 0 -2.0 1e-06 
0.0 0.8878 0 -2.0 1e-06 
0.0 0.8879 0 -2.0 1e-06 
0.0 0.888 0 -2.0 1e-06 
0.0 0.8881 0 -2.0 1e-06 
0.0 0.8882 0 -2.0 1e-06 
0.0 0.8883 0 -2.0 1e-06 
0.0 0.8884 0 -2.0 1e-06 
0.0 0.8885 0 -2.0 1e-06 
0.0 0.8886 0 -2.0 1e-06 
0.0 0.8887 0 -2.0 1e-06 
0.0 0.8888 0 -2.0 1e-06 
0.0 0.8889 0 -2.0 1e-06 
0.0 0.889 0 -2.0 1e-06 
0.0 0.8891 0 -2.0 1e-06 
0.0 0.8892 0 -2.0 1e-06 
0.0 0.8893 0 -2.0 1e-06 
0.0 0.8894 0 -2.0 1e-06 
0.0 0.8895 0 -2.0 1e-06 
0.0 0.8896 0 -2.0 1e-06 
0.0 0.8897 0 -2.0 1e-06 
0.0 0.8898 0 -2.0 1e-06 
0.0 0.8899 0 -2.0 1e-06 
0.0 0.89 0 -2.0 1e-06 
0.0 0.8901 0 -2.0 1e-06 
0.0 0.8902 0 -2.0 1e-06 
0.0 0.8903 0 -2.0 1e-06 
0.0 0.8904 0 -2.0 1e-06 
0.0 0.8905 0 -2.0 1e-06 
0.0 0.8906 0 -2.0 1e-06 
0.0 0.8907 0 -2.0 1e-06 
0.0 0.8908 0 -2.0 1e-06 
0.0 0.8909 0 -2.0 1e-06 
0.0 0.891 0 -2.0 1e-06 
0.0 0.8911 0 -2.0 1e-06 
0.0 0.8912 0 -2.0 1e-06 
0.0 0.8913 0 -2.0 1e-06 
0.0 0.8914 0 -2.0 1e-06 
0.0 0.8915 0 -2.0 1e-06 
0.0 0.8916 0 -2.0 1e-06 
0.0 0.8917 0 -2.0 1e-06 
0.0 0.8918 0 -2.0 1e-06 
0.0 0.8919 0 -2.0 1e-06 
0.0 0.892 0 -2.0 1e-06 
0.0 0.8921 0 -2.0 1e-06 
0.0 0.8922 0 -2.0 1e-06 
0.0 0.8923 0 -2.0 1e-06 
0.0 0.8924 0 -2.0 1e-06 
0.0 0.8925 0 -2.0 1e-06 
0.0 0.8926 0 -2.0 1e-06 
0.0 0.8927 0 -2.0 1e-06 
0.0 0.8928 0 -2.0 1e-06 
0.0 0.8929 0 -2.0 1e-06 
0.0 0.893 0 -2.0 1e-06 
0.0 0.8931 0 -2.0 1e-06 
0.0 0.8932 0 -2.0 1e-06 
0.0 0.8933 0 -2.0 1e-06 
0.0 0.8934 0 -2.0 1e-06 
0.0 0.8935 0 -2.0 1e-06 
0.0 0.8936 0 -2.0 1e-06 
0.0 0.8937 0 -2.0 1e-06 
0.0 0.8938 0 -2.0 1e-06 
0.0 0.8939 0 -2.0 1e-06 
0.0 0.894 0 -2.0 1e-06 
0.0 0.8941 0 -2.0 1e-06 
0.0 0.8942 0 -2.0 1e-06 
0.0 0.8943 0 -2.0 1e-06 
0.0 0.8944 0 -2.0 1e-06 
0.0 0.8945 0 -2.0 1e-06 
0.0 0.8946 0 -2.0 1e-06 
0.0 0.8947 0 -2.0 1e-06 
0.0 0.8948 0 -2.0 1e-06 
0.0 0.8949 0 -2.0 1e-06 
0.0 0.895 0 -2.0 1e-06 
0.0 0.8951 0 -2.0 1e-06 
0.0 0.8952 0 -2.0 1e-06 
0.0 0.8953 0 -2.0 1e-06 
0.0 0.8954 0 -2.0 1e-06 
0.0 0.8955 0 -2.0 1e-06 
0.0 0.8956 0 -2.0 1e-06 
0.0 0.8957 0 -2.0 1e-06 
0.0 0.8958 0 -2.0 1e-06 
0.0 0.8959 0 -2.0 1e-06 
0.0 0.896 0 -2.0 1e-06 
0.0 0.8961 0 -2.0 1e-06 
0.0 0.8962 0 -2.0 1e-06 
0.0 0.8963 0 -2.0 1e-06 
0.0 0.8964 0 -2.0 1e-06 
0.0 0.8965 0 -2.0 1e-06 
0.0 0.8966 0 -2.0 1e-06 
0.0 0.8967 0 -2.0 1e-06 
0.0 0.8968 0 -2.0 1e-06 
0.0 0.8969 0 -2.0 1e-06 
0.0 0.897 0 -2.0 1e-06 
0.0 0.8971 0 -2.0 1e-06 
0.0 0.8972 0 -2.0 1e-06 
0.0 0.8973 0 -2.0 1e-06 
0.0 0.8974 0 -2.0 1e-06 
0.0 0.8975 0 -2.0 1e-06 
0.0 0.8976 0 -2.0 1e-06 
0.0 0.8977 0 -2.0 1e-06 
0.0 0.8978 0 -2.0 1e-06 
0.0 0.8979 0 -2.0 1e-06 
0.0 0.898 0 -2.0 1e-06 
0.0 0.8981 0 -2.0 1e-06 
0.0 0.8982 0 -2.0 1e-06 
0.0 0.8983 0 -2.0 1e-06 
0.0 0.8984 0 -2.0 1e-06 
0.0 0.8985 0 -2.0 1e-06 
0.0 0.8986 0 -2.0 1e-06 
0.0 0.8987 0 -2.0 1e-06 
0.0 0.8988 0 -2.0 1e-06 
0.0 0.8989 0 -2.0 1e-06 
0.0 0.899 0 -2.0 1e-06 
0.0 0.8991 0 -2.0 1e-06 
0.0 0.8992 0 -2.0 1e-06 
0.0 0.8993 0 -2.0 1e-06 
0.0 0.8994 0 -2.0 1e-06 
0.0 0.8995 0 -2.0 1e-06 
0.0 0.8996 0 -2.0 1e-06 
0.0 0.8997 0 -2.0 1e-06 
0.0 0.8998 0 -2.0 1e-06 
0.0 0.8999 0 -2.0 1e-06 
0.0 0.9 0 -2.0 1e-06 
0.0 0.9001 0 -2.0 1e-06 
0.0 0.9002 0 -2.0 1e-06 
0.0 0.9003 0 -2.0 1e-06 
0.0 0.9004 0 -2.0 1e-06 
0.0 0.9005 0 -2.0 1e-06 
0.0 0.9006 0 -2.0 1e-06 
0.0 0.9007 0 -2.0 1e-06 
0.0 0.9008 0 -2.0 1e-06 
0.0 0.9009 0 -2.0 1e-06 
0.0 0.901 0 -2.0 1e-06 
0.0 0.9011 0 -2.0 1e-06 
0.0 0.9012 0 -2.0 1e-06 
0.0 0.9013 0 -2.0 1e-06 
0.0 0.9014 0 -2.0 1e-06 
0.0 0.9015 0 -2.0 1e-06 
0.0 0.9016 0 -2.0 1e-06 
0.0 0.9017 0 -2.0 1e-06 
0.0 0.9018 0 -2.0 1e-06 
0.0 0.9019 0 -2.0 1e-06 
0.0 0.902 0 -2.0 1e-06 
0.0 0.9021 0 -2.0 1e-06 
0.0 0.9022 0 -2.0 1e-06 
0.0 0.9023 0 -2.0 1e-06 
0.0 0.9024 0 -2.0 1e-06 
0.0 0.9025 0 -2.0 1e-06 
0.0 0.9026 0 -2.0 1e-06 
0.0 0.9027 0 -2.0 1e-06 
0.0 0.9028 0 -2.0 1e-06 
0.0 0.9029 0 -2.0 1e-06 
0.0 0.903 0 -2.0 1e-06 
0.0 0.9031 0 -2.0 1e-06 
0.0 0.9032 0 -2.0 1e-06 
0.0 0.9033 0 -2.0 1e-06 
0.0 0.9034 0 -2.0 1e-06 
0.0 0.9035 0 -2.0 1e-06 
0.0 0.9036 0 -2.0 1e-06 
0.0 0.9037 0 -2.0 1e-06 
0.0 0.9038 0 -2.0 1e-06 
0.0 0.9039 0 -2.0 1e-06 
0.0 0.904 0 -2.0 1e-06 
0.0 0.9041 0 -2.0 1e-06 
0.0 0.9042 0 -2.0 1e-06 
0.0 0.9043 0 -2.0 1e-06 
0.0 0.9044 0 -2.0 1e-06 
0.0 0.9045 0 -2.0 1e-06 
0.0 0.9046 0 -2.0 1e-06 
0.0 0.9047 0 -2.0 1e-06 
0.0 0.9048 0 -2.0 1e-06 
0.0 0.9049 0 -2.0 1e-06 
0.0 0.905 0 -2.0 1e-06 
0.0 0.9051 0 -2.0 1e-06 
0.0 0.9052 0 -2.0 1e-06 
0.0 0.9053 0 -2.0 1e-06 
0.0 0.9054 0 -2.0 1e-06 
0.0 0.9055 0 -2.0 1e-06 
0.0 0.9056 0 -2.0 1e-06 
0.0 0.9057 0 -2.0 1e-06 
0.0 0.9058 0 -2.0 1e-06 
0.0 0.9059 0 -2.0 1e-06 
0.0 0.906 0 -2.0 1e-06 
0.0 0.9061 0 -2.0 1e-06 
0.0 0.9062 0 -2.0 1e-06 
0.0 0.9063 0 -2.0 1e-06 
0.0 0.9064 0 -2.0 1e-06 
0.0 0.9065 0 -2.0 1e-06 
0.0 0.9066 0 -2.0 1e-06 
0.0 0.9067 0 -2.0 1e-06 
0.0 0.9068 0 -2.0 1e-06 
0.0 0.9069 0 -2.0 1e-06 
0.0 0.907 0 -2.0 1e-06 
0.0 0.9071 0 -2.0 1e-06 
0.0 0.9072 0 -2.0 1e-06 
0.0 0.9073 0 -2.0 1e-06 
0.0 0.9074 0 -2.0 1e-06 
0.0 0.9075 0 -2.0 1e-06 
0.0 0.9076 0 -2.0 1e-06 
0.0 0.9077 0 -2.0 1e-06 
0.0 0.9078 0 -2.0 1e-06 
0.0 0.9079 0 -2.0 1e-06 
0.0 0.908 0 -2.0 1e-06 
0.0 0.9081 0 -2.0 1e-06 
0.0 0.9082 0 -2.0 1e-06 
0.0 0.9083 0 -2.0 1e-06 
0.0 0.9084 0 -2.0 1e-06 
0.0 0.9085 0 -2.0 1e-06 
0.0 0.9086 0 -2.0 1e-06 
0.0 0.9087 0 -2.0 1e-06 
0.0 0.9088 0 -2.0 1e-06 
0.0 0.9089 0 -2.0 1e-06 
0.0 0.909 0 -2.0 1e-06 
0.0 0.9091 0 -2.0 1e-06 
0.0 0.9092 0 -2.0 1e-06 
0.0 0.9093 0 -2.0 1e-06 
0.0 0.9094 0 -2.0 1e-06 
0.0 0.9095 0 -2.0 1e-06 
0.0 0.9096 0 -2.0 1e-06 
0.0 0.9097 0 -2.0 1e-06 
0.0 0.9098 0 -2.0 1e-06 
0.0 0.9099 0 -2.0 1e-06 
0.0 0.91 0 -2.0 1e-06 
0.0 0.9101 0 -2.0 1e-06 
0.0 0.9102 0 -2.0 1e-06 
0.0 0.9103 0 -2.0 1e-06 
0.0 0.9104 0 -2.0 1e-06 
0.0 0.9105 0 -2.0 1e-06 
0.0 0.9106 0 -2.0 1e-06 
0.0 0.9107 0 -2.0 1e-06 
0.0 0.9108 0 -2.0 1e-06 
0.0 0.9109 0 -2.0 1e-06 
0.0 0.911 0 -2.0 1e-06 
0.0 0.9111 0 -2.0 1e-06 
0.0 0.9112 0 -2.0 1e-06 
0.0 0.9113 0 -2.0 1e-06 
0.0 0.9114 0 -2.0 1e-06 
0.0 0.9115 0 -2.0 1e-06 
0.0 0.9116 0 -2.0 1e-06 
0.0 0.9117 0 -2.0 1e-06 
0.0 0.9118 0 -2.0 1e-06 
0.0 0.9119 0 -2.0 1e-06 
0.0 0.912 0 -2.0 1e-06 
0.0 0.9121 0 -2.0 1e-06 
0.0 0.9122 0 -2.0 1e-06 
0.0 0.9123 0 -2.0 1e-06 
0.0 0.9124 0 -2.0 1e-06 
0.0 0.9125 0 -2.0 1e-06 
0.0 0.9126 0 -2.0 1e-06 
0.0 0.9127 0 -2.0 1e-06 
0.0 0.9128 0 -2.0 1e-06 
0.0 0.9129 0 -2.0 1e-06 
0.0 0.913 0 -2.0 1e-06 
0.0 0.9131 0 -2.0 1e-06 
0.0 0.9132 0 -2.0 1e-06 
0.0 0.9133 0 -2.0 1e-06 
0.0 0.9134 0 -2.0 1e-06 
0.0 0.9135 0 -2.0 1e-06 
0.0 0.9136 0 -2.0 1e-06 
0.0 0.9137 0 -2.0 1e-06 
0.0 0.9138 0 -2.0 1e-06 
0.0 0.9139 0 -2.0 1e-06 
0.0 0.914 0 -2.0 1e-06 
0.0 0.9141 0 -2.0 1e-06 
0.0 0.9142 0 -2.0 1e-06 
0.0 0.9143 0 -2.0 1e-06 
0.0 0.9144 0 -2.0 1e-06 
0.0 0.9145 0 -2.0 1e-06 
0.0 0.9146 0 -2.0 1e-06 
0.0 0.9147 0 -2.0 1e-06 
0.0 0.9148 0 -2.0 1e-06 
0.0 0.9149 0 -2.0 1e-06 
0.0 0.915 0 -2.0 1e-06 
0.0 0.9151 0 -2.0 1e-06 
0.0 0.9152 0 -2.0 1e-06 
0.0 0.9153 0 -2.0 1e-06 
0.0 0.9154 0 -2.0 1e-06 
0.0 0.9155 0 -2.0 1e-06 
0.0 0.9156 0 -2.0 1e-06 
0.0 0.9157 0 -2.0 1e-06 
0.0 0.9158 0 -2.0 1e-06 
0.0 0.9159 0 -2.0 1e-06 
0.0 0.916 0 -2.0 1e-06 
0.0 0.9161 0 -2.0 1e-06 
0.0 0.9162 0 -2.0 1e-06 
0.0 0.9163 0 -2.0 1e-06 
0.0 0.9164 0 -2.0 1e-06 
0.0 0.9165 0 -2.0 1e-06 
0.0 0.9166 0 -2.0 1e-06 
0.0 0.9167 0 -2.0 1e-06 
0.0 0.9168 0 -2.0 1e-06 
0.0 0.9169 0 -2.0 1e-06 
0.0 0.917 0 -2.0 1e-06 
0.0 0.9171 0 -2.0 1e-06 
0.0 0.9172 0 -2.0 1e-06 
0.0 0.9173 0 -2.0 1e-06 
0.0 0.9174 0 -2.0 1e-06 
0.0 0.9175 0 -2.0 1e-06 
0.0 0.9176 0 -2.0 1e-06 
0.0 0.9177 0 -2.0 1e-06 
0.0 0.9178 0 -2.0 1e-06 
0.0 0.9179 0 -2.0 1e-06 
0.0 0.918 0 -2.0 1e-06 
0.0 0.9181 0 -2.0 1e-06 
0.0 0.9182 0 -2.0 1e-06 
0.0 0.9183 0 -2.0 1e-06 
0.0 0.9184 0 -2.0 1e-06 
0.0 0.9185 0 -2.0 1e-06 
0.0 0.9186 0 -2.0 1e-06 
0.0 0.9187 0 -2.0 1e-06 
0.0 0.9188 0 -2.0 1e-06 
0.0 0.9189 0 -2.0 1e-06 
0.0 0.919 0 -2.0 1e-06 
0.0 0.9191 0 -2.0 1e-06 
0.0 0.9192 0 -2.0 1e-06 
0.0 0.9193 0 -2.0 1e-06 
0.0 0.9194 0 -2.0 1e-06 
0.0 0.9195 0 -2.0 1e-06 
0.0 0.9196 0 -2.0 1e-06 
0.0 0.9197 0 -2.0 1e-06 
0.0 0.9198 0 -2.0 1e-06 
0.0 0.9199 0 -2.0 1e-06 
0.0 0.92 0 -2.0 1e-06 
0.0 0.9201 0 -2.0 1e-06 
0.0 0.9202 0 -2.0 1e-06 
0.0 0.9203 0 -2.0 1e-06 
0.0 0.9204 0 -2.0 1e-06 
0.0 0.9205 0 -2.0 1e-06 
0.0 0.9206 0 -2.0 1e-06 
0.0 0.9207 0 -2.0 1e-06 
0.0 0.9208 0 -2.0 1e-06 
0.0 0.9209 0 -2.0 1e-06 
0.0 0.921 0 -2.0 1e-06 
0.0 0.9211 0 -2.0 1e-06 
0.0 0.9212 0 -2.0 1e-06 
0.0 0.9213 0 -2.0 1e-06 
0.0 0.9214 0 -2.0 1e-06 
0.0 0.9215 0 -2.0 1e-06 
0.0 0.9216 0 -2.0 1e-06 
0.0 0.9217 0 -2.0 1e-06 
0.0 0.9218 0 -2.0 1e-06 
0.0 0.9219 0 -2.0 1e-06 
0.0 0.922 0 -2.0 1e-06 
0.0 0.9221 0 -2.0 1e-06 
0.0 0.9222 0 -2.0 1e-06 
0.0 0.9223 0 -2.0 1e-06 
0.0 0.9224 0 -2.0 1e-06 
0.0 0.9225 0 -2.0 1e-06 
0.0 0.9226 0 -2.0 1e-06 
0.0 0.9227 0 -2.0 1e-06 
0.0 0.9228 0 -2.0 1e-06 
0.0 0.9229 0 -2.0 1e-06 
0.0 0.923 0 -2.0 1e-06 
0.0 0.9231 0 -2.0 1e-06 
0.0 0.9232 0 -2.0 1e-06 
0.0 0.9233 0 -2.0 1e-06 
0.0 0.9234 0 -2.0 1e-06 
0.0 0.9235 0 -2.0 1e-06 
0.0 0.9236 0 -2.0 1e-06 
0.0 0.9237 0 -2.0 1e-06 
0.0 0.9238 0 -2.0 1e-06 
0.0 0.9239 0 -2.0 1e-06 
0.0 0.924 0 -2.0 1e-06 
0.0 0.9241 0 -2.0 1e-06 
0.0 0.9242 0 -2.0 1e-06 
0.0 0.9243 0 -2.0 1e-06 
0.0 0.9244 0 -2.0 1e-06 
0.0 0.9245 0 -2.0 1e-06 
0.0 0.9246 0 -2.0 1e-06 
0.0 0.9247 0 -2.0 1e-06 
0.0 0.9248 0 -2.0 1e-06 
0.0 0.9249 0 -2.0 1e-06 
0.0 0.925 0 -2.0 1e-06 
0.0 0.9251 0 -2.0 1e-06 
0.0 0.9252 0 -2.0 1e-06 
0.0 0.9253 0 -2.0 1e-06 
0.0 0.9254 0 -2.0 1e-06 
0.0 0.9255 0 -2.0 1e-06 
0.0 0.9256 0 -2.0 1e-06 
0.0 0.9257 0 -2.0 1e-06 
0.0 0.9258 0 -2.0 1e-06 
0.0 0.9259 0 -2.0 1e-06 
0.0 0.926 0 -2.0 1e-06 
0.0 0.9261 0 -2.0 1e-06 
0.0 0.9262 0 -2.0 1e-06 
0.0 0.9263 0 -2.0 1e-06 
0.0 0.9264 0 -2.0 1e-06 
0.0 0.9265 0 -2.0 1e-06 
0.0 0.9266 0 -2.0 1e-06 
0.0 0.9267 0 -2.0 1e-06 
0.0 0.9268 0 -2.0 1e-06 
0.0 0.9269 0 -2.0 1e-06 
0.0 0.927 0 -2.0 1e-06 
0.0 0.9271 0 -2.0 1e-06 
0.0 0.9272 0 -2.0 1e-06 
0.0 0.9273 0 -2.0 1e-06 
0.0 0.9274 0 -2.0 1e-06 
0.0 0.9275 0 -2.0 1e-06 
0.0 0.9276 0 -2.0 1e-06 
0.0 0.9277 0 -2.0 1e-06 
0.0 0.9278 0 -2.0 1e-06 
0.0 0.9279 0 -2.0 1e-06 
0.0 0.928 0 -2.0 1e-06 
0.0 0.9281 0 -2.0 1e-06 
0.0 0.9282 0 -2.0 1e-06 
0.0 0.9283 0 -2.0 1e-06 
0.0 0.9284 0 -2.0 1e-06 
0.0 0.9285 0 -2.0 1e-06 
0.0 0.9286 0 -2.0 1e-06 
0.0 0.9287 0 -2.0 1e-06 
0.0 0.9288 0 -2.0 1e-06 
0.0 0.9289 0 -2.0 1e-06 
0.0 0.929 0 -2.0 1e-06 
0.0 0.9291 0 -2.0 1e-06 
0.0 0.9292 0 -2.0 1e-06 
0.0 0.9293 0 -2.0 1e-06 
0.0 0.9294 0 -2.0 1e-06 
0.0 0.9295 0 -2.0 1e-06 
0.0 0.9296 0 -2.0 1e-06 
0.0 0.9297 0 -2.0 1e-06 
0.0 0.9298 0 -2.0 1e-06 
0.0 0.9299 0 -2.0 1e-06 
0.0 0.93 0 -2.0 1e-06 
0.0 0.9301 0 -2.0 1e-06 
0.0 0.9302 0 -2.0 1e-06 
0.0 0.9303 0 -2.0 1e-06 
0.0 0.9304 0 -2.0 1e-06 
0.0 0.9305 0 -2.0 1e-06 
0.0 0.9306 0 -2.0 1e-06 
0.0 0.9307 0 -2.0 1e-06 
0.0 0.9308 0 -2.0 1e-06 
0.0 0.9309 0 -2.0 1e-06 
0.0 0.931 0 -2.0 1e-06 
0.0 0.9311 0 -2.0 1e-06 
0.0 0.9312 0 -2.0 1e-06 
0.0 0.9313 0 -2.0 1e-06 
0.0 0.9314 0 -2.0 1e-06 
0.0 0.9315 0 -2.0 1e-06 
0.0 0.9316 0 -2.0 1e-06 
0.0 0.9317 0 -2.0 1e-06 
0.0 0.9318 0 -2.0 1e-06 
0.0 0.9319 0 -2.0 1e-06 
0.0 0.932 0 -2.0 1e-06 
0.0 0.9321 0 -2.0 1e-06 
0.0 0.9322 0 -2.0 1e-06 
0.0 0.9323 0 -2.0 1e-06 
0.0 0.9324 0 -2.0 1e-06 
0.0 0.9325 0 -2.0 1e-06 
0.0 0.9326 0 -2.0 1e-06 
0.0 0.9327 0 -2.0 1e-06 
0.0 0.9328 0 -2.0 1e-06 
0.0 0.9329 0 -2.0 1e-06 
0.0 0.933 0 -2.0 1e-06 
0.0 0.9331 0 -2.0 1e-06 
0.0 0.9332 0 -2.0 1e-06 
0.0 0.9333 0 -2.0 1e-06 
0.0 0.9334 0 -2.0 1e-06 
0.0 0.9335 0 -2.0 1e-06 
0.0 0.9336 0 -2.0 1e-06 
0.0 0.9337 0 -2.0 1e-06 
0.0 0.9338 0 -2.0 1e-06 
0.0 0.9339 0 -2.0 1e-06 
0.0 0.934 0 -2.0 1e-06 
0.0 0.9341 0 -2.0 1e-06 
0.0 0.9342 0 -2.0 1e-06 
0.0 0.9343 0 -2.0 1e-06 
0.0 0.9344 0 -2.0 1e-06 
0.0 0.9345 0 -2.0 1e-06 
0.0 0.9346 0 -2.0 1e-06 
0.0 0.9347 0 -2.0 1e-06 
0.0 0.9348 0 -2.0 1e-06 
0.0 0.9349 0 -2.0 1e-06 
0.0 0.935 0 -2.0 1e-06 
0.0 0.9351 0 -2.0 1e-06 
0.0 0.9352 0 -2.0 1e-06 
0.0 0.9353 0 -2.0 1e-06 
0.0 0.9354 0 -2.0 1e-06 
0.0 0.9355 0 -2.0 1e-06 
0.0 0.9356 0 -2.0 1e-06 
0.0 0.9357 0 -2.0 1e-06 
0.0 0.9358 0 -2.0 1e-06 
0.0 0.9359 0 -2.0 1e-06 
0.0 0.936 0 -2.0 1e-06 
0.0 0.9361 0 -2.0 1e-06 
0.0 0.9362 0 -2.0 1e-06 
0.0 0.9363 0 -2.0 1e-06 
0.0 0.9364 0 -2.0 1e-06 
0.0 0.9365 0 -2.0 1e-06 
0.0 0.9366 0 -2.0 1e-06 
0.0 0.9367 0 -2.0 1e-06 
0.0 0.9368 0 -2.0 1e-06 
0.0 0.9369 0 -2.0 1e-06 
0.0 0.937 0 -2.0 1e-06 
0.0 0.9371 0 -2.0 1e-06 
0.0 0.9372 0 -2.0 1e-06 
0.0 0.9373 0 -2.0 1e-06 
0.0 0.9374 0 -2.0 1e-06 
0.0 0.9375 0 -2.0 1e-06 
0.0 0.9376 0 -2.0 1e-06 
0.0 0.9377 0 -2.0 1e-06 
0.0 0.9378 0 -2.0 1e-06 
0.0 0.9379 0 -2.0 1e-06 
0.0 0.938 0 -2.0 1e-06 
0.0 0.9381 0 -2.0 1e-06 
0.0 0.9382 0 -2.0 1e-06 
0.0 0.9383 0 -2.0 1e-06 
0.0 0.9384 0 -2.0 1e-06 
0.0 0.9385 0 -2.0 1e-06 
0.0 0.9386 0 -2.0 1e-06 
0.0 0.9387 0 -2.0 1e-06 
0.0 0.9388 0 -2.0 1e-06 
0.0 0.9389 0 -2.0 1e-06 
0.0 0.939 0 -2.0 1e-06 
0.0 0.9391 0 -2.0 1e-06 
0.0 0.9392 0 -2.0 1e-06 
0.0 0.9393 0 -2.0 1e-06 
0.0 0.9394 0 -2.0 1e-06 
0.0 0.9395 0 -2.0 1e-06 
0.0 0.9396 0 -2.0 1e-06 
0.0 0.9397 0 -2.0 1e-06 
0.0 0.9398 0 -2.0 1e-06 
0.0 0.9399 0 -2.0 1e-06 
0.0 0.94 0 -2.0 1e-06 
0.0 0.9401 0 -2.0 1e-06 
0.0 0.9402 0 -2.0 1e-06 
0.0 0.9403 0 -2.0 1e-06 
0.0 0.9404 0 -2.0 1e-06 
0.0 0.9405 0 -2.0 1e-06 
0.0 0.9406 0 -2.0 1e-06 
0.0 0.9407 0 -2.0 1e-06 
0.0 0.9408 0 -2.0 1e-06 
0.0 0.9409 0 -2.0 1e-06 
0.0 0.941 0 -2.0 1e-06 
0.0 0.9411 0 -2.0 1e-06 
0.0 0.9412 0 -2.0 1e-06 
0.0 0.9413 0 -2.0 1e-06 
0.0 0.9414 0 -2.0 1e-06 
0.0 0.9415 0 -2.0 1e-06 
0.0 0.9416 0 -2.0 1e-06 
0.0 0.9417 0 -2.0 1e-06 
0.0 0.9418 0 -2.0 1e-06 
0.0 0.9419 0 -2.0 1e-06 
0.0 0.942 0 -2.0 1e-06 
0.0 0.9421 0 -2.0 1e-06 
0.0 0.9422 0 -2.0 1e-06 
0.0 0.9423 0 -2.0 1e-06 
0.0 0.9424 0 -2.0 1e-06 
0.0 0.9425 0 -2.0 1e-06 
0.0 0.9426 0 -2.0 1e-06 
0.0 0.9427 0 -2.0 1e-06 
0.0 0.9428 0 -2.0 1e-06 
0.0 0.9429 0 -2.0 1e-06 
0.0 0.943 0 -2.0 1e-06 
0.0 0.9431 0 -2.0 1e-06 
0.0 0.9432 0 -2.0 1e-06 
0.0 0.9433 0 -2.0 1e-06 
0.0 0.9434 0 -2.0 1e-06 
0.0 0.9435 0 -2.0 1e-06 
0.0 0.9436 0 -2.0 1e-06 
0.0 0.9437 0 -2.0 1e-06 
0.0 0.9438 0 -2.0 1e-06 
0.0 0.9439 0 -2.0 1e-06 
0.0 0.944 0 -2.0 1e-06 
0.0 0.9441 0 -2.0 1e-06 
0.0 0.9442 0 -2.0 1e-06 
0.0 0.9443 0 -2.0 1e-06 
0.0 0.9444 0 -2.0 1e-06 
0.0 0.9445 0 -2.0 1e-06 
0.0 0.9446 0 -2.0 1e-06 
0.0 0.9447 0 -2.0 1e-06 
0.0 0.9448 0 -2.0 1e-06 
0.0 0.9449 0 -2.0 1e-06 
0.0 0.945 0 -2.0 1e-06 
0.0 0.9451 0 -2.0 1e-06 
0.0 0.9452 0 -2.0 1e-06 
0.0 0.9453 0 -2.0 1e-06 
0.0 0.9454 0 -2.0 1e-06 
0.0 0.9455 0 -2.0 1e-06 
0.0 0.9456 0 -2.0 1e-06 
0.0 0.9457 0 -2.0 1e-06 
0.0 0.9458 0 -2.0 1e-06 
0.0 0.9459 0 -2.0 1e-06 
0.0 0.946 0 -2.0 1e-06 
0.0 0.9461 0 -2.0 1e-06 
0.0 0.9462 0 -2.0 1e-06 
0.0 0.9463 0 -2.0 1e-06 
0.0 0.9464 0 -2.0 1e-06 
0.0 0.9465 0 -2.0 1e-06 
0.0 0.9466 0 -2.0 1e-06 
0.0 0.9467 0 -2.0 1e-06 
0.0 0.9468 0 -2.0 1e-06 
0.0 0.9469 0 -2.0 1e-06 
0.0 0.947 0 -2.0 1e-06 
0.0 0.9471 0 -2.0 1e-06 
0.0 0.9472 0 -2.0 1e-06 
0.0 0.9473 0 -2.0 1e-06 
0.0 0.9474 0 -2.0 1e-06 
0.0 0.9475 0 -2.0 1e-06 
0.0 0.9476 0 -2.0 1e-06 
0.0 0.9477 0 -2.0 1e-06 
0.0 0.9478 0 -2.0 1e-06 
0.0 0.9479 0 -2.0 1e-06 
0.0 0.948 0 -2.0 1e-06 
0.0 0.9481 0 -2.0 1e-06 
0.0 0.9482 0 -2.0 1e-06 
0.0 0.9483 0 -2.0 1e-06 
0.0 0.9484 0 -2.0 1e-06 
0.0 0.9485 0 -2.0 1e-06 
0.0 0.9486 0 -2.0 1e-06 
0.0 0.9487 0 -2.0 1e-06 
0.0 0.9488 0 -2.0 1e-06 
0.0 0.9489 0 -2.0 1e-06 
0.0 0.949 0 -2.0 1e-06 
0.0 0.9491 0 -2.0 1e-06 
0.0 0.9492 0 -2.0 1e-06 
0.0 0.9493 0 -2.0 1e-06 
0.0 0.9494 0 -2.0 1e-06 
0.0 0.9495 0 -2.0 1e-06 
0.0 0.9496 0 -2.0 1e-06 
0.0 0.9497 0 -2.0 1e-06 
0.0 0.9498 0 -2.0 1e-06 
0.0 0.9499 0 -2.0 1e-06 
0.0 0.95 0 -2.0 1e-06 
0.0 0.9501 0 -2.0 1e-06 
0.0 0.9502 0 -2.0 1e-06 
0.0 0.9503 0 -2.0 1e-06 
0.0 0.9504 0 -2.0 1e-06 
0.0 0.9505 0 -2.0 1e-06 
0.0 0.9506 0 -2.0 1e-06 
0.0 0.9507 0 -2.0 1e-06 
0.0 0.9508 0 -2.0 1e-06 
0.0 0.9509 0 -2.0 1e-06 
0.0 0.951 0 -2.0 1e-06 
0.0 0.9511 0 -2.0 1e-06 
0.0 0.9512 0 -2.0 1e-06 
0.0 0.9513 0 -2.0 1e-06 
0.0 0.9514 0 -2.0 1e-06 
0.0 0.9515 0 -2.0 1e-06 
0.0 0.9516 0 -2.0 1e-06 
0.0 0.9517 0 -2.0 1e-06 
0.0 0.9518 0 -2.0 1e-06 
0.0 0.9519 0 -2.0 1e-06 
0.0 0.952 0 -2.0 1e-06 
0.0 0.9521 0 -2.0 1e-06 
0.0 0.9522 0 -2.0 1e-06 
0.0 0.9523 0 -2.0 1e-06 
0.0 0.9524 0 -2.0 1e-06 
0.0 0.9525 0 -2.0 1e-06 
0.0 0.9526 0 -2.0 1e-06 
0.0 0.9527 0 -2.0 1e-06 
0.0 0.9528 0 -2.0 1e-06 
0.0 0.9529 0 -2.0 1e-06 
0.0 0.953 0 -2.0 1e-06 
0.0 0.9531 0 -2.0 1e-06 
0.0 0.9532 0 -2.0 1e-06 
0.0 0.9533 0 -2.0 1e-06 
0.0 0.9534 0 -2.0 1e-06 
0.0 0.9535 0 -2.0 1e-06 
0.0 0.9536 0 -2.0 1e-06 
0.0 0.9537 0 -2.0 1e-06 
0.0 0.9538 0 -2.0 1e-06 
0.0 0.9539 0 -2.0 1e-06 
0.0 0.954 0 -2.0 1e-06 
0.0 0.9541 0 -2.0 1e-06 
0.0 0.9542 0 -2.0 1e-06 
0.0 0.9543 0 -2.0 1e-06 
0.0 0.9544 0 -2.0 1e-06 
0.0 0.9545 0 -2.0 1e-06 
0.0 0.9546 0 -2.0 1e-06 
0.0 0.9547 0 -2.0 1e-06 
0.0 0.9548 0 -2.0 1e-06 
0.0 0.9549 0 -2.0 1e-06 
0.0 0.955 0 -2.0 1e-06 
0.0 0.9551 0 -2.0 1e-06 
0.0 0.9552 0 -2.0 1e-06 
0.0 0.9553 0 -2.0 1e-06 
0.0 0.9554 0 -2.0 1e-06 
0.0 0.9555 0 -2.0 1e-06 
0.0 0.9556 0 -2.0 1e-06 
0.0 0.9557 0 -2.0 1e-06 
0.0 0.9558 0 -2.0 1e-06 
0.0 0.9559 0 -2.0 1e-06 
0.0 0.956 0 -2.0 1e-06 
0.0 0.9561 0 -2.0 1e-06 
0.0 0.9562 0 -2.0 1e-06 
0.0 0.9563 0 -2.0 1e-06 
0.0 0.9564 0 -2.0 1e-06 
0.0 0.9565 0 -2.0 1e-06 
0.0 0.9566 0 -2.0 1e-06 
0.0 0.9567 0 -2.0 1e-06 
0.0 0.9568 0 -2.0 1e-06 
0.0 0.9569 0 -2.0 1e-06 
0.0 0.957 0 -2.0 1e-06 
0.0 0.9571 0 -2.0 1e-06 
0.0 0.9572 0 -2.0 1e-06 
0.0 0.9573 0 -2.0 1e-06 
0.0 0.9574 0 -2.0 1e-06 
0.0 0.9575 0 -2.0 1e-06 
0.0 0.9576 0 -2.0 1e-06 
0.0 0.9577 0 -2.0 1e-06 
0.0 0.9578 0 -2.0 1e-06 
0.0 0.9579 0 -2.0 1e-06 
0.0 0.958 0 -2.0 1e-06 
0.0 0.9581 0 -2.0 1e-06 
0.0 0.9582 0 -2.0 1e-06 
0.0 0.9583 0 -2.0 1e-06 
0.0 0.9584 0 -2.0 1e-06 
0.0 0.9585 0 -2.0 1e-06 
0.0 0.9586 0 -2.0 1e-06 
0.0 0.9587 0 -2.0 1e-06 
0.0 0.9588 0 -2.0 1e-06 
0.0 0.9589 0 -2.0 1e-06 
0.0 0.959 0 -2.0 1e-06 
0.0 0.9591 0 -2.0 1e-06 
0.0 0.9592 0 -2.0 1e-06 
0.0 0.9593 0 -2.0 1e-06 
0.0 0.9594 0 -2.0 1e-06 
0.0 0.9595 0 -2.0 1e-06 
0.0 0.9596 0 -2.0 1e-06 
0.0 0.9597 0 -2.0 1e-06 
0.0 0.9598 0 -2.0 1e-06 
0.0 0.9599 0 -2.0 1e-06 
0.0 0.96 0 -2.0 1e-06 
0.0 0.9601 0 -2.0 1e-06 
0.0 0.9602 0 -2.0 1e-06 
0.0 0.9603 0 -2.0 1e-06 
0.0 0.9604 0 -2.0 1e-06 
0.0 0.9605 0 -2.0 1e-06 
0.0 0.9606 0 -2.0 1e-06 
0.0 0.9607 0 -2.0 1e-06 
0.0 0.9608 0 -2.0 1e-06 
0.0 0.9609 0 -2.0 1e-06 
0.0 0.961 0 -2.0 1e-06 
0.0 0.9611 0 -2.0 1e-06 
0.0 0.9612 0 -2.0 1e-06 
0.0 0.9613 0 -2.0 1e-06 
0.0 0.9614 0 -2.0 1e-06 
0.0 0.9615 0 -2.0 1e-06 
0.0 0.9616 0 -2.0 1e-06 
0.0 0.9617 0 -2.0 1e-06 
0.0 0.9618 0 -2.0 1e-06 
0.0 0.9619 0 -2.0 1e-06 
0.0 0.962 0 -2.0 1e-06 
0.0 0.9621 0 -2.0 1e-06 
0.0 0.9622 0 -2.0 1e-06 
0.0 0.9623 0 -2.0 1e-06 
0.0 0.9624 0 -2.0 1e-06 
0.0 0.9625 0 -2.0 1e-06 
0.0 0.9626 0 -2.0 1e-06 
0.0 0.9627 0 -2.0 1e-06 
0.0 0.9628 0 -2.0 1e-06 
0.0 0.9629 0 -2.0 1e-06 
0.0 0.963 0 -2.0 1e-06 
0.0 0.9631 0 -2.0 1e-06 
0.0 0.9632 0 -2.0 1e-06 
0.0 0.9633 0 -2.0 1e-06 
0.0 0.9634 0 -2.0 1e-06 
0.0 0.9635 0 -2.0 1e-06 
0.0 0.9636 0 -2.0 1e-06 
0.0 0.9637 0 -2.0 1e-06 
0.0 0.9638 0 -2.0 1e-06 
0.0 0.9639 0 -2.0 1e-06 
0.0 0.964 0 -2.0 1e-06 
0.0 0.9641 0 -2.0 1e-06 
0.0 0.9642 0 -2.0 1e-06 
0.0 0.9643 0 -2.0 1e-06 
0.0 0.9644 0 -2.0 1e-06 
0.0 0.9645 0 -2.0 1e-06 
0.0 0.9646 0 -2.0 1e-06 
0.0 0.9647 0 -2.0 1e-06 
0.0 0.9648 0 -2.0 1e-06 
0.0 0.9649 0 -2.0 1e-06 
0.0 0.965 0 -2.0 1e-06 
0.0 0.9651 0 -2.0 1e-06 
0.0 0.9652 0 -2.0 1e-06 
0.0 0.9653 0 -2.0 1e-06 
0.0 0.9654 0 -2.0 1e-06 
0.0 0.9655 0 -2.0 1e-06 
0.0 0.9656 0 -2.0 1e-06 
0.0 0.9657 0 -2.0 1e-06 
0.0 0.9658 0 -2.0 1e-06 
0.0 0.9659 0 -2.0 1e-06 
0.0 0.966 0 -2.0 1e-06 
0.0 0.9661 0 -2.0 1e-06 
0.0 0.9662 0 -2.0 1e-06 
0.0 0.9663 0 -2.0 1e-06 
0.0 0.9664 0 -2.0 1e-06 
0.0 0.9665 0 -2.0 1e-06 
0.0 0.9666 0 -2.0 1e-06 
0.0 0.9667 0 -2.0 1e-06 
0.0 0.9668 0 -2.0 1e-06 
0.0 0.9669 0 -2.0 1e-06 
0.0 0.967 0 -2.0 1e-06 
0.0 0.9671 0 -2.0 1e-06 
0.0 0.9672 0 -2.0 1e-06 
0.0 0.9673 0 -2.0 1e-06 
0.0 0.9674 0 -2.0 1e-06 
0.0 0.9675 0 -2.0 1e-06 
0.0 0.9676 0 -2.0 1e-06 
0.0 0.9677 0 -2.0 1e-06 
0.0 0.9678 0 -2.0 1e-06 
0.0 0.9679 0 -2.0 1e-06 
0.0 0.968 0 -2.0 1e-06 
0.0 0.9681 0 -2.0 1e-06 
0.0 0.9682 0 -2.0 1e-06 
0.0 0.9683 0 -2.0 1e-06 
0.0 0.9684 0 -2.0 1e-06 
0.0 0.9685 0 -2.0 1e-06 
0.0 0.9686 0 -2.0 1e-06 
0.0 0.9687 0 -2.0 1e-06 
0.0 0.9688 0 -2.0 1e-06 
0.0 0.9689 0 -2.0 1e-06 
0.0 0.969 0 -2.0 1e-06 
0.0 0.9691 0 -2.0 1e-06 
0.0 0.9692 0 -2.0 1e-06 
0.0 0.9693 0 -2.0 1e-06 
0.0 0.9694 0 -2.0 1e-06 
0.0 0.9695 0 -2.0 1e-06 
0.0 0.9696 0 -2.0 1e-06 
0.0 0.9697 0 -2.0 1e-06 
0.0 0.9698 0 -2.0 1e-06 
0.0 0.9699 0 -2.0 1e-06 
0.0 0.97 0 -2.0 1e-06 
0.0 0.9701 0 -2.0 1e-06 
0.0 0.9702 0 -2.0 1e-06 
0.0 0.9703 0 -2.0 1e-06 
0.0 0.9704 0 -2.0 1e-06 
0.0 0.9705 0 -2.0 1e-06 
0.0 0.9706 0 -2.0 1e-06 
0.0 0.9707 0 -2.0 1e-06 
0.0 0.9708 0 -2.0 1e-06 
0.0 0.9709 0 -2.0 1e-06 
0.0 0.971 0 -2.0 1e-06 
0.0 0.9711 0 -2.0 1e-06 
0.0 0.9712 0 -2.0 1e-06 
0.0 0.9713 0 -2.0 1e-06 
0.0 0.9714 0 -2.0 1e-06 
0.0 0.9715 0 -2.0 1e-06 
0.0 0.9716 0 -2.0 1e-06 
0.0 0.9717 0 -2.0 1e-06 
0.0 0.9718 0 -2.0 1e-06 
0.0 0.9719 0 -2.0 1e-06 
0.0 0.972 0 -2.0 1e-06 
0.0 0.9721 0 -2.0 1e-06 
0.0 0.9722 0 -2.0 1e-06 
0.0 0.9723 0 -2.0 1e-06 
0.0 0.9724 0 -2.0 1e-06 
0.0 0.9725 0 -2.0 1e-06 
0.0 0.9726 0 -2.0 1e-06 
0.0 0.9727 0 -2.0 1e-06 
0.0 0.9728 0 -2.0 1e-06 
0.0 0.9729 0 -2.0 1e-06 
0.0 0.973 0 -2.0 1e-06 
0.0 0.9731 0 -2.0 1e-06 
0.0 0.9732 0 -2.0 1e-06 
0.0 0.9733 0 -2.0 1e-06 
0.0 0.9734 0 -2.0 1e-06 
0.0 0.9735 0 -2.0 1e-06 
0.0 0.9736 0 -2.0 1e-06 
0.0 0.9737 0 -2.0 1e-06 
0.0 0.9738 0 -2.0 1e-06 
0.0 0.9739 0 -2.0 1e-06 
0.0 0.974 0 -2.0 1e-06 
0.0 0.9741 0 -2.0 1e-06 
0.0 0.9742 0 -2.0 1e-06 
0.0 0.9743 0 -2.0 1e-06 
0.0 0.9744 0 -2.0 1e-06 
0.0 0.9745 0 -2.0 1e-06 
0.0 0.9746 0 -2.0 1e-06 
0.0 0.9747 0 -2.0 1e-06 
0.0 0.9748 0 -2.0 1e-06 
0.0 0.9749 0 -2.0 1e-06 
0.0 0.975 0 -2.0 1e-06 
0.0 0.9751 0 -2.0 1e-06 
0.0 0.9752 0 -2.0 1e-06 
0.0 0.9753 0 -2.0 1e-06 
0.0 0.9754 0 -2.0 1e-06 
0.0 0.9755 0 -2.0 1e-06 
0.0 0.9756 0 -2.0 1e-06 
0.0 0.9757 0 -2.0 1e-06 
0.0 0.9758 0 -2.0 1e-06 
0.0 0.9759 0 -2.0 1e-06 
0.0 0.976 0 -2.0 1e-06 
0.0 0.9761 0 -2.0 1e-06 
0.0 0.9762 0 -2.0 1e-06 
0.0 0.9763 0 -2.0 1e-06 
0.0 0.9764 0 -2.0 1e-06 
0.0 0.9765 0 -2.0 1e-06 
0.0 0.9766 0 -2.0 1e-06 
0.0 0.9767 0 -2.0 1e-06 
0.0 0.9768 0 -2.0 1e-06 
0.0 0.9769 0 -2.0 1e-06 
0.0 0.977 0 -2.0 1e-06 
0.0 0.9771 0 -2.0 1e-06 
0.0 0.9772 0 -2.0 1e-06 
0.0 0.9773 0 -2.0 1e-06 
0.0 0.9774 0 -2.0 1e-06 
0.0 0.9775 0 -2.0 1e-06 
0.0 0.9776 0 -2.0 1e-06 
0.0 0.9777 0 -2.0 1e-06 
0.0 0.9778 0 -2.0 1e-06 
0.0 0.9779 0 -2.0 1e-06 
0.0 0.978 0 -2.0 1e-06 
0.0 0.9781 0 -2.0 1e-06 
0.0 0.9782 0 -2.0 1e-06 
0.0 0.9783 0 -2.0 1e-06 
0.0 0.9784 0 -2.0 1e-06 
0.0 0.9785 0 -2.0 1e-06 
0.0 0.9786 0 -2.0 1e-06 
0.0 0.9787 0 -2.0 1e-06 
0.0 0.9788 0 -2.0 1e-06 
0.0 0.9789 0 -2.0 1e-06 
0.0 0.979 0 -2.0 1e-06 
0.0 0.9791 0 -2.0 1e-06 
0.0 0.9792 0 -2.0 1e-06 
0.0 0.9793 0 -2.0 1e-06 
0.0 0.9794 0 -2.0 1e-06 
0.0 0.9795 0 -2.0 1e-06 
0.0 0.9796 0 -2.0 1e-06 
0.0 0.9797 0 -2.0 1e-06 
0.0 0.9798 0 -2.0 1e-06 
0.0 0.9799 0 -2.0 1e-06 
0.0 0.98 0 -2.0 1e-06 
0.0 0.9801 0 -2.0 1e-06 
0.0 0.9802 0 -2.0 1e-06 
0.0 0.9803 0 -2.0 1e-06 
0.0 0.9804 0 -2.0 1e-06 
0.0 0.9805 0 -2.0 1e-06 
0.0 0.9806 0 -2.0 1e-06 
0.0 0.9807 0 -2.0 1e-06 
0.0 0.9808 0 -2.0 1e-06 
0.0 0.9809 0 -2.0 1e-06 
0.0 0.981 0 -2.0 1e-06 
0.0 0.9811 0 -2.0 1e-06 
0.0 0.9812 0 -2.0 1e-06 
0.0 0.9813 0 -2.0 1e-06 
0.0 0.9814 0 -2.0 1e-06 
0.0 0.9815 0 -2.0 1e-06 
0.0 0.9816 0 -2.0 1e-06 
0.0 0.9817 0 -2.0 1e-06 
0.0 0.9818 0 -2.0 1e-06 
0.0 0.9819 0 -2.0 1e-06 
0.0 0.982 0 -2.0 1e-06 
0.0 0.9821 0 -2.0 1e-06 
0.0 0.9822 0 -2.0 1e-06 
0.0 0.9823 0 -2.0 1e-06 
0.0 0.9824 0 -2.0 1e-06 
0.0 0.9825 0 -2.0 1e-06 
0.0 0.9826 0 -2.0 1e-06 
0.0 0.9827 0 -2.0 1e-06 
0.0 0.9828 0 -2.0 1e-06 
0.0 0.9829 0 -2.0 1e-06 
0.0 0.983 0 -2.0 1e-06 
0.0 0.9831 0 -2.0 1e-06 
0.0 0.9832 0 -2.0 1e-06 
0.0 0.9833 0 -2.0 1e-06 
0.0 0.9834 0 -2.0 1e-06 
0.0 0.9835 0 -2.0 1e-06 
0.0 0.9836 0 -2.0 1e-06 
0.0 0.9837 0 -2.0 1e-06 
0.0 0.9838 0 -2.0 1e-06 
0.0 0.9839 0 -2.0 1e-06 
0.0 0.984 0 -2.0 1e-06 
0.0 0.9841 0 -2.0 1e-06 
0.0 0.9842 0 -2.0 1e-06 
0.0 0.9843 0 -2.0 1e-06 
0.0 0.9844 0 -2.0 1e-06 
0.0 0.9845 0 -2.0 1e-06 
0.0 0.9846 0 -2.0 1e-06 
0.0 0.9847 0 -2.0 1e-06 
0.0 0.9848 0 -2.0 1e-06 
0.0 0.9849 0 -2.0 1e-06 
0.0 0.985 0 -2.0 1e-06 
0.0 0.9851 0 -2.0 1e-06 
0.0 0.9852 0 -2.0 1e-06 
0.0 0.9853 0 -2.0 1e-06 
0.0 0.9854 0 -2.0 1e-06 
0.0 0.9855 0 -2.0 1e-06 
0.0 0.9856 0 -2.0 1e-06 
0.0 0.9857 0 -2.0 1e-06 
0.0 0.9858 0 -2.0 1e-06 
0.0 0.9859 0 -2.0 1e-06 
0.0 0.986 0 -2.0 1e-06 
0.0 0.9861 0 -2.0 1e-06 
0.0 0.9862 0 -2.0 1e-06 
0.0 0.9863 0 -2.0 1e-06 
0.0 0.9864 0 -2.0 1e-06 
0.0 0.9865 0 -2.0 1e-06 
0.0 0.9866 0 -2.0 1e-06 
0.0 0.9867 0 -2.0 1e-06 
0.0 0.9868 0 -2.0 1e-06 
0.0 0.9869 0 -2.0 1e-06 
0.0 0.987 0 -2.0 1e-06 
0.0 0.9871 0 -2.0 1e-06 
0.0 0.9872 0 -2.0 1e-06 
0.0 0.9873 0 -2.0 1e-06 
0.0 0.9874 0 -2.0 1e-06 
0.0 0.9875 0 -2.0 1e-06 
0.0 0.9876 0 -2.0 1e-06 
0.0 0.9877 0 -2.0 1e-06 
0.0 0.9878 0 -2.0 1e-06 
0.0 0.9879 0 -2.0 1e-06 
0.0 0.988 0 -2.0 1e-06 
0.0 0.9881 0 -2.0 1e-06 
0.0 0.9882 0 -2.0 1e-06 
0.0 0.9883 0 -2.0 1e-06 
0.0 0.9884 0 -2.0 1e-06 
0.0 0.9885 0 -2.0 1e-06 
0.0 0.9886 0 -2.0 1e-06 
0.0 0.9887 0 -2.0 1e-06 
0.0 0.9888 0 -2.0 1e-06 
0.0 0.9889 0 -2.0 1e-06 
0.0 0.989 0 -2.0 1e-06 
0.0 0.9891 0 -2.0 1e-06 
0.0 0.9892 0 -2.0 1e-06 
0.0 0.9893 0 -2.0 1e-06 
0.0 0.9894 0 -2.0 1e-06 
0.0 0.9895 0 -2.0 1e-06 
0.0 0.9896 0 -2.0 1e-06 
0.0 0.9897 0 -2.0 1e-06 
0.0 0.9898 0 -2.0 1e-06 
0.0 0.9899 0 -2.0 1e-06 
0.0 0.99 0 -2.0 1e-06 
0.0 0.9901 0 -2.0 1e-06 
0.0 0.9902 0 -2.0 1e-06 
0.0 0.9903 0 -2.0 1e-06 
0.0 0.9904 0 -2.0 1e-06 
0.0 0.9905 0 -2.0 1e-06 
0.0 0.9906 0 -2.0 1e-06 
0.0 0.9907 0 -2.0 1e-06 
0.0 0.9908 0 -2.0 1e-06 
0.0 0.9909 0 -2.0 1e-06 
0.0 0.991 0 -2.0 1e-06 
0.0 0.9911 0 -2.0 1e-06 
0.0 0.9912 0 -2.0 1e-06 
0.0 0.9913 0 -2.0 1e-06 
0.0 0.9914 0 -2.0 1e-06 
0.0 0.9915 0 -2.0 1e-06 
0.0 0.9916 0 -2.0 1e-06 
0.0 0.9917 0 -2.0 1e-06 
0.0 0.9918 0 -2.0 1e-06 
0.0 0.9919 0 -2.0 1e-06 
0.0 0.992 0 -2.0 1e-06 
0.0 0.9921 0 -2.0 1e-06 
0.0 0.9922 0 -2.0 1e-06 
0.0 0.9923 0 -2.0 1e-06 
0.0 0.9924 0 -2.0 1e-06 
0.0 0.9925 0 -2.0 1e-06 
0.0 0.9926 0 -2.0 1e-06 
0.0 0.9927 0 -2.0 1e-06 
0.0 0.9928 0 -2.0 1e-06 
0.0 0.9929 0 -2.0 1e-06 
0.0 0.993 0 -2.0 1e-06 
0.0 0.9931 0 -2.0 1e-06 
0.0 0.9932 0 -2.0 1e-06 
0.0 0.9933 0 -2.0 1e-06 
0.0 0.9934 0 -2.0 1e-06 
0.0 0.9935 0 -2.0 1e-06 
0.0 0.9936 0 -2.0 1e-06 
0.0 0.9937 0 -2.0 1e-06 
0.0 0.9938 0 -2.0 1e-06 
0.0 0.9939 0 -2.0 1e-06 
0.0 0.994 0 -2.0 1e-06 
0.0 0.9941 0 -2.0 1e-06 
0.0 0.9942 0 -2.0 1e-06 
0.0 0.9943 0 -2.0 1e-06 
0.0 0.9944 0 -2.0 1e-06 
0.0 0.9945 0 -2.0 1e-06 
0.0 0.9946 0 -2.0 1e-06 
0.0 0.9947 0 -2.0 1e-06 
0.0 0.9948 0 -2.0 1e-06 
0.0 0.9949 0 -2.0 1e-06 
0.0 0.995 0 -2.0 1e-06 
0.0 0.9951 0 -2.0 1e-06 
0.0 0.9952 0 -2.0 1e-06 
0.0 0.9953 0 -2.0 1e-06 
0.0 0.9954 0 -2.0 1e-06 
0.0 0.9955 0 -2.0 1e-06 
0.0 0.9956 0 -2.0 1e-06 
0.0 0.9957 0 -2.0 1e-06 
0.0 0.9958 0 -2.0 1e-06 
0.0 0.9959 0 -2.0 1e-06 
0.0 0.996 0 -2.0 1e-06 
0.0 0.9961 0 -2.0 1e-06 
0.0 0.9962 0 -2.0 1e-06 
0.0 0.9963 0 -2.0 1e-06 
0.0 0.9964 0 -2.0 1e-06 
0.0 0.9965 0 -2.0 1e-06 
0.0 0.9966 0 -2.0 1e-06 
0.0 0.9967 0 -2.0 1e-06 
0.0 0.9968 0 -2.0 1e-06 
0.0 0.9969 0 -2.0 1e-06 
0.0 0.997 0 -2.0 1e-06 
0.0 0.9971 0 -2.0 1e-06 
0.0 0.9972 0 -2.0 1e-06 
0.0 0.9973 0 -2.0 1e-06 
0.0 0.9974 0 -2.0 1e-06 
0.0 0.9975 0 -2.0 1e-06 
0.0 0.9976 0 -2.0 1e-06 
0.0 0.9977 0 -2.0 1e-06 
0.0 0.9978 0 -2.0 1e-06 
0.0 0.9979 0 -2.0 1e-06 
0.0 0.998 0 -2.0 1e-06 
0.0 0.9981 0 -2.0 1e-06 
0.0 0.9982 0 -2.0 1e-06 
0.0 0.9983 0 -2.0 1e-06 
0.0 0.9984 0 -2.0 1e-06 
0.0 0.9985 0 -2.0 1e-06 
0.0 0.9986 0 -2.0 1e-06 
0.0 0.9987 0 -2.0 1e-06 
0.0 0.9988 0 -2.0 1e-06 
0.0 0.9989 0 -2.0 1e-06 
0.0 0.999 0 -2.0 1e-06 
0.0 0.9991 0 -2.0 1e-06 
0.0 0.9992 0 -2.0 1e-06 
0.0 0.9993 0 -2.0 1e-06 
0.0 0.9994 0 -2.0 1e-06 
0.0 0.9995 0 -2.0 1e-06 
0.0 0.9996 0 -2.0 1e-06 
0.0 0.9997 0 -2.0 1e-06 
0.0 0.9998 0 -2.0 1e-06 
0.0 0.9999 0 -2.0 1e-06 
0.0 1.0 0 -2.0 1e-06 
0.0 1.0001 0 -2.0 1e-06 
0.0 1.0002 0 -2.0 1e-06 
0.0 1.0003 0 -2.0 1e-06 
0.0 1.0004 0 -2.0 1e-06 
0.0 1.0005 0 -2.0 1e-06 
0.0 1.0006 0 -2.0 1e-06 
0.0 1.0007 0 -2.0 1e-06 
0.0 1.0008 0 -2.0 1e-06 
0.0 1.0009 0 -2.0 1e-06 
0.0 1.001 0 -2.0 1e-06 
0.0 1.0011 0 -2.0 1e-06 
0.0 1.0012 0 -2.0 1e-06 
0.0 1.0013 0 -2.0 1e-06 
0.0 1.0014 0 -2.0 1e-06 
0.0 1.0015 0 -2.0 1e-06 
0.0 1.0016 0 -2.0 1e-06 
0.0 1.0017 0 -2.0 1e-06 
0.0 1.0018 0 -2.0 1e-06 
0.0 1.0019 0 -2.0 1e-06 
0.0 1.002 0 -2.0 1e-06 
0.0 1.0021 0 -2.0 1e-06 
0.0 1.0022 0 -2.0 1e-06 
0.0 1.0023 0 -2.0 1e-06 
0.0 1.0024 0 -2.0 1e-06 
0.0 1.0025 0 -2.0 1e-06 
0.0 1.0026 0 -2.0 1e-06 
0.0 1.0027 0 -2.0 1e-06 
0.0 1.0028 0 -2.0 1e-06 
0.0 1.0029 0 -2.0 1e-06 
0.0 1.003 0 -2.0 1e-06 
0.0 1.0031 0 -2.0 1e-06 
0.0 1.0032 0 -2.0 1e-06 
0.0 1.0033 0 -2.0 1e-06 
0.0 1.0034 0 -2.0 1e-06 
0.0 1.0035 0 -2.0 1e-06 
0.0 1.0036 0 -2.0 1e-06 
0.0 1.0037 0 -2.0 1e-06 
0.0 1.0038 0 -2.0 1e-06 
0.0 1.0039 0 -2.0 1e-06 
0.0 1.004 0 -2.0 1e-06 
0.0 1.0041 0 -2.0 1e-06 
0.0 1.0042 0 -2.0 1e-06 
0.0 1.0043 0 -2.0 1e-06 
0.0 1.0044 0 -2.0 1e-06 
0.0 1.0045 0 -2.0 1e-06 
0.0 1.0046 0 -2.0 1e-06 
0.0 1.0047 0 -2.0 1e-06 
0.0 1.0048 0 -2.0 1e-06 
0.0 1.0049 0 -2.0 1e-06 
0.0 1.005 0 -2.0 1e-06 
0.0 1.0051 0 -2.0 1e-06 
0.0 1.0052 0 -2.0 1e-06 
0.0 1.0053 0 -2.0 1e-06 
0.0 1.0054 0 -2.0 1e-06 
0.0 1.0055 0 -2.0 1e-06 
0.0 1.0056 0 -2.0 1e-06 
0.0 1.0057 0 -2.0 1e-06 
0.0 1.0058 0 -2.0 1e-06 
0.0 1.0059 0 -2.0 1e-06 
0.0 1.006 0 -2.0 1e-06 
0.0 1.0061 0 -2.0 1e-06 
0.0 1.0062 0 -2.0 1e-06 
0.0 1.0063 0 -2.0 1e-06 
0.0 1.0064 0 -2.0 1e-06 
0.0 1.0065 0 -2.0 1e-06 
0.0 1.0066 0 -2.0 1e-06 
0.0 1.0067 0 -2.0 1e-06 
0.0 1.0068 0 -2.0 1e-06 
0.0 1.0069 0 -2.0 1e-06 
0.0 1.007 0 -2.0 1e-06 
0.0 1.0071 0 -2.0 1e-06 
0.0 1.0072 0 -2.0 1e-06 
0.0 1.0073 0 -2.0 1e-06 
0.0 1.0074 0 -2.0 1e-06 
0.0 1.0075 0 -2.0 1e-06 
0.0 1.0076 0 -2.0 1e-06 
0.0 1.0077 0 -2.0 1e-06 
0.0 1.0078 0 -2.0 1e-06 
0.0 1.0079 0 -2.0 1e-06 
0.0 1.008 0 -2.0 1e-06 
0.0 1.0081 0 -2.0 1e-06 
0.0 1.0082 0 -2.0 1e-06 
0.0 1.0083 0 -2.0 1e-06 
0.0 1.0084 0 -2.0 1e-06 
0.0 1.0085 0 -2.0 1e-06 
0.0 1.0086 0 -2.0 1e-06 
0.0 1.0087 0 -2.0 1e-06 
0.0 1.0088 0 -2.0 1e-06 
0.0 1.0089 0 -2.0 1e-06 
0.0 1.009 0 -2.0 1e-06 
0.0 1.0091 0 -2.0 1e-06 
0.0 1.0092 0 -2.0 1e-06 
0.0 1.0093 0 -2.0 1e-06 
0.0 1.0094 0 -2.0 1e-06 
0.0 1.0095 0 -2.0 1e-06 
0.0 1.0096 0 -2.0 1e-06 
0.0 1.0097 0 -2.0 1e-06 
0.0 1.0098 0 -2.0 1e-06 
0.0 1.0099 0 -2.0 1e-06 
0.0 1.01 0 -2.0 1e-06 
0.0 1.0101 0 -2.0 1e-06 
0.0 1.0102 0 -2.0 1e-06 
0.0 1.0103 0 -2.0 1e-06 
0.0 1.0104 0 -2.0 1e-06 
0.0 1.0105 0 -2.0 1e-06 
0.0 1.0106 0 -2.0 1e-06 
0.0 1.0107 0 -2.0 1e-06 
0.0 1.0108 0 -2.0 1e-06 
0.0 1.0109 0 -2.0 1e-06 
0.0 1.011 0 -2.0 1e-06 
0.0 1.0111 0 -2.0 1e-06 
0.0 1.0112 0 -2.0 1e-06 
0.0 1.0113 0 -2.0 1e-06 
0.0 1.0114 0 -2.0 1e-06 
0.0 1.0115 0 -2.0 1e-06 
0.0 1.0116 0 -2.0 1e-06 
0.0 1.0117 0 -2.0 1e-06 
0.0 1.0118 0 -2.0 1e-06 
0.0 1.0119 0 -2.0 1e-06 
0.0 1.012 0 -2.0 1e-06 
0.0 1.0121 0 -2.0 1e-06 
0.0 1.0122 0 -2.0 1e-06 
0.0 1.0123 0 -2.0 1e-06 
0.0 1.0124 0 -2.0 1e-06 
0.0 1.0125 0 -2.0 1e-06 
0.0 1.0126 0 -2.0 1e-06 
0.0 1.0127 0 -2.0 1e-06 
0.0 1.0128 0 -2.0 1e-06 
0.0 1.0129 0 -2.0 1e-06 
0.0 1.013 0 -2.0 1e-06 
0.0 1.0131 0 -2.0 1e-06 
0.0 1.0132 0 -2.0 1e-06 
0.0 1.0133 0 -2.0 1e-06 
0.0 1.0134 0 -2.0 1e-06 
0.0 1.0135 0 -2.0 1e-06 
0.0 1.0136 0 -2.0 1e-06 
0.0 1.0137 0 -2.0 1e-06 
0.0 1.0138 0 -2.0 1e-06 
0.0 1.0139 0 -2.0 1e-06 
0.0 1.014 0 -2.0 1e-06 
0.0 1.0141 0 -2.0 1e-06 
0.0 1.0142 0 -2.0 1e-06 
0.0 1.0143 0 -2.0 1e-06 
0.0 1.0144 0 -2.0 1e-06 
0.0 1.0145 0 -2.0 1e-06 
0.0 1.0146 0 -2.0 1e-06 
0.0 1.0147 0 -2.0 1e-06 
0.0 1.0148 0 -2.0 1e-06 
0.0 1.0149 0 -2.0 1e-06 
0.0 1.015 0 -2.0 1e-06 
0.0 1.0151 0 -2.0 1e-06 
0.0 1.0152 0 -2.0 1e-06 
0.0 1.0153 0 -2.0 1e-06 
0.0 1.0154 0 -2.0 1e-06 
0.0 1.0155 0 -2.0 1e-06 
0.0 1.0156 0 -2.0 1e-06 
0.0 1.0157 0 -2.0 1e-06 
0.0 1.0158 0 -2.0 1e-06 
0.0 1.0159 0 -2.0 1e-06 
0.0 1.016 0 -2.0 1e-06 
0.0 1.0161 0 -2.0 1e-06 
0.0 1.0162 0 -2.0 1e-06 
0.0 1.0163 0 -2.0 1e-06 
0.0 1.0164 0 -2.0 1e-06 
0.0 1.0165 0 -2.0 1e-06 
0.0 1.0166 0 -2.0 1e-06 
0.0 1.0167 0 -2.0 1e-06 
0.0 1.0168 0 -2.0 1e-06 
0.0 1.0169 0 -2.0 1e-06 
0.0 1.017 0 -2.0 1e-06 
0.0 1.0171 0 -2.0 1e-06 
0.0 1.0172 0 -2.0 1e-06 
0.0 1.0173 0 -2.0 1e-06 
0.0 1.0174 0 -2.0 1e-06 
0.0 1.0175 0 -2.0 1e-06 
0.0 1.0176 0 -2.0 1e-06 
0.0 1.0177 0 -2.0 1e-06 
0.0 1.0178 0 -2.0 1e-06 
0.0 1.0179 0 -2.0 1e-06 
0.0 1.018 0 -2.0 1e-06 
0.0 1.0181 0 -2.0 1e-06 
0.0 1.0182 0 -2.0 1e-06 
0.0 1.0183 0 -2.0 1e-06 
0.0 1.0184 0 -2.0 1e-06 
0.0 1.0185 0 -2.0 1e-06 
0.0 1.0186 0 -2.0 1e-06 
0.0 1.0187 0 -2.0 1e-06 
0.0 1.0188 0 -2.0 1e-06 
0.0 1.0189 0 -2.0 1e-06 
0.0 1.019 0 -2.0 1e-06 
0.0 1.0191 0 -2.0 1e-06 
0.0 1.0192 0 -2.0 1e-06 
0.0 1.0193 0 -2.0 1e-06 
0.0 1.0194 0 -2.0 1e-06 
0.0 1.0195 0 -2.0 1e-06 
0.0 1.0196 0 -2.0 1e-06 
0.0 1.0197 0 -2.0 1e-06 
0.0 1.0198 0 -2.0 1e-06 
0.0 1.0199 0 -2.0 1e-06 
0.0 1.02 0 -2.0 1e-06 
0.0 1.0201 0 -2.0 1e-06 
0.0 1.0202 0 -2.0 1e-06 
0.0 1.0203 0 -2.0 1e-06 
0.0 1.0204 0 -2.0 1e-06 
0.0 1.0205 0 -2.0 1e-06 
0.0 1.0206 0 -2.0 1e-06 
0.0 1.0207 0 -2.0 1e-06 
0.0 1.0208 0 -2.0 1e-06 
0.0 1.0209 0 -2.0 1e-06 
0.0 1.021 0 -2.0 1e-06 
0.0 1.0211 0 -2.0 1e-06 
0.0 1.0212 0 -2.0 1e-06 
0.0 1.0213 0 -2.0 1e-06 
0.0 1.0214 0 -2.0 1e-06 
0.0 1.0215 0 -2.0 1e-06 
0.0 1.0216 0 -2.0 1e-06 
0.0 1.0217 0 -2.0 1e-06 
0.0 1.0218 0 -2.0 1e-06 
0.0 1.0219 0 -2.0 1e-06 
0.0 1.022 0 -2.0 1e-06 
0.0 1.0221 0 -2.0 1e-06 
0.0 1.0222 0 -2.0 1e-06 
0.0 1.0223 0 -2.0 1e-06 
0.0 1.0224 0 -2.0 1e-06 
0.0 1.0225 0 -2.0 1e-06 
0.0 1.0226 0 -2.0 1e-06 
0.0 1.0227 0 -2.0 1e-06 
0.0 1.0228 0 -2.0 1e-06 
0.0 1.0229 0 -2.0 1e-06 
0.0 1.023 0 -2.0 1e-06 
0.0 1.0231 0 -2.0 1e-06 
0.0 1.0232 0 -2.0 1e-06 
0.0 1.0233 0 -2.0 1e-06 
0.0 1.0234 0 -2.0 1e-06 
0.0 1.0235 0 -2.0 1e-06 
0.0 1.0236 0 -2.0 1e-06 
0.0 1.0237 0 -2.0 1e-06 
0.0 1.0238 0 -2.0 1e-06 
0.0 1.0239 0 -2.0 1e-06 
0.0 1.024 0 -2.0 1e-06 
0.0 1.0241 0 -2.0 1e-06 
0.0 1.0242 0 -2.0 1e-06 
0.0 1.0243 0 -2.0 1e-06 
0.0 1.0244 0 -2.0 1e-06 
0.0 1.0245 0 -2.0 1e-06 
0.0 1.0246 0 -2.0 1e-06 
0.0 1.0247 0 -2.0 1e-06 
0.0 1.0248 0 -2.0 1e-06 
0.0 1.0249 0 -2.0 1e-06 
0.0 1.025 0 -2.0 1e-06 
0.0 1.0251 0 -2.0 1e-06 
0.0 1.0252 0 -2.0 1e-06 
0.0 1.0253 0 -2.0 1e-06 
0.0 1.0254 0 -2.0 1e-06 
0.0 1.0255 0 -2.0 1e-06 
0.0 1.0256 0 -2.0 1e-06 
0.0 1.0257 0 -2.0 1e-06 
0.0 1.0258 0 -2.0 1e-06 
0.0 1.0259 0 -2.0 1e-06 
0.0 1.026 0 -2.0 1e-06 
0.0 1.0261 0 -2.0 1e-06 
0.0 1.0262 0 -2.0 1e-06 
0.0 1.0263 0 -2.0 1e-06 
0.0 1.0264 0 -2.0 1e-06 
0.0 1.0265 0 -2.0 1e-06 
0.0 1.0266 0 -2.0 1e-06 
0.0 1.0267 0 -2.0 1e-06 
0.0 1.0268 0 -2.0 1e-06 
0.0 1.0269 0 -2.0 1e-06 
0.0 1.027 0 -2.0 1e-06 
0.0 1.0271 0 -2.0 1e-06 
0.0 1.0272 0 -2.0 1e-06 
0.0 1.0273 0 -2.0 1e-06 
0.0 1.0274 0 -2.0 1e-06 
0.0 1.0275 0 -2.0 1e-06 
0.0 1.0276 0 -2.0 1e-06 
0.0 1.0277 0 -2.0 1e-06 
0.0 1.0278 0 -2.0 1e-06 
0.0 1.0279 0 -2.0 1e-06 
0.0 1.028 0 -2.0 1e-06 
0.0 1.0281 0 -2.0 1e-06 
0.0 1.0282 0 -2.0 1e-06 
0.0 1.0283 0 -2.0 1e-06 
0.0 1.0284 0 -2.0 1e-06 
0.0 1.0285 0 -2.0 1e-06 
0.0 1.0286 0 -2.0 1e-06 
0.0 1.0287 0 -2.0 1e-06 
0.0 1.0288 0 -2.0 1e-06 
0.0 1.0289 0 -2.0 1e-06 
0.0 1.029 0 -2.0 1e-06 
0.0 1.0291 0 -2.0 1e-06 
0.0 1.0292 0 -2.0 1e-06 
0.0 1.0293 0 -2.0 1e-06 
0.0 1.0294 0 -2.0 1e-06 
0.0 1.0295 0 -2.0 1e-06 
0.0 1.0296 0 -2.0 1e-06 
0.0 1.0297 0 -2.0 1e-06 
0.0 1.0298 0 -2.0 1e-06 
0.0 1.0299 0 -2.0 1e-06 
0.0 1.03 0 -2.0 1e-06 
0.0 1.0301 0 -2.0 1e-06 
0.0 1.0302 0 -2.0 1e-06 
0.0 1.0303 0 -2.0 1e-06 
0.0 1.0304 0 -2.0 1e-06 
0.0 1.0305 0 -2.0 1e-06 
0.0 1.0306 0 -2.0 1e-06 
0.0 1.0307 0 -2.0 1e-06 
0.0 1.0308 0 -2.0 1e-06 
0.0 1.0309 0 -2.0 1e-06 
0.0 1.031 0 -2.0 1e-06 
0.0 1.0311 0 -2.0 1e-06 
0.0 1.0312 0 -2.0 1e-06 
0.0 1.0313 0 -2.0 1e-06 
0.0 1.0314 0 -2.0 1e-06 
0.0 1.0315 0 -2.0 1e-06 
0.0 1.0316 0 -2.0 1e-06 
0.0 1.0317 0 -2.0 1e-06 
0.0 1.0318 0 -2.0 1e-06 
0.0 1.0319 0 -2.0 1e-06 
0.0 1.032 0 -2.0 1e-06 
0.0 1.0321 0 -2.0 1e-06 
0.0 1.0322 0 -2.0 1e-06 
0.0 1.0323 0 -2.0 1e-06 
0.0 1.0324 0 -2.0 1e-06 
0.0 1.0325 0 -2.0 1e-06 
0.0 1.0326 0 -2.0 1e-06 
0.0 1.0327 0 -2.0 1e-06 
0.0 1.0328 0 -2.0 1e-06 
0.0 1.0329 0 -2.0 1e-06 
0.0 1.033 0 -2.0 1e-06 
0.0 1.0331 0 -2.0 1e-06 
0.0 1.0332 0 -2.0 1e-06 
0.0 1.0333 0 -2.0 1e-06 
0.0 1.0334 0 -2.0 1e-06 
0.0 1.0335 0 -2.0 1e-06 
0.0 1.0336 0 -2.0 1e-06 
0.0 1.0337 0 -2.0 1e-06 
0.0 1.0338 0 -2.0 1e-06 
0.0 1.0339 0 -2.0 1e-06 
0.0 1.034 0 -2.0 1e-06 
0.0 1.0341 0 -2.0 1e-06 
0.0 1.0342 0 -2.0 1e-06 
0.0 1.0343 0 -2.0 1e-06 
0.0 1.0344 0 -2.0 1e-06 
0.0 1.0345 0 -2.0 1e-06 
0.0 1.0346 0 -2.0 1e-06 
0.0 1.0347 0 -2.0 1e-06 
0.0 1.0348 0 -2.0 1e-06 
0.0 1.0349 0 -2.0 1e-06 
0.0 1.035 0 -2.0 1e-06 
0.0 1.0351 0 -2.0 1e-06 
0.0 1.0352 0 -2.0 1e-06 
0.0 1.0353 0 -2.0 1e-06 
0.0 1.0354 0 -2.0 1e-06 
0.0 1.0355 0 -2.0 1e-06 
0.0 1.0356 0 -2.0 1e-06 
0.0 1.0357 0 -2.0 1e-06 
0.0 1.0358 0 -2.0 1e-06 
0.0 1.0359 0 -2.0 1e-06 
0.0 1.036 0 -2.0 1e-06 
0.0 1.0361 0 -2.0 1e-06 
0.0 1.0362 0 -2.0 1e-06 
0.0 1.0363 0 -2.0 1e-06 
0.0 1.0364 0 -2.0 1e-06 
0.0 1.0365 0 -2.0 1e-06 
0.0 1.0366 0 -2.0 1e-06 
0.0 1.0367 0 -2.0 1e-06 
0.0 1.0368 0 -2.0 1e-06 
0.0 1.0369 0 -2.0 1e-06 
0.0 1.037 0 -2.0 1e-06 
0.0 1.0371 0 -2.0 1e-06 
0.0 1.0372 0 -2.0 1e-06 
0.0 1.0373 0 -2.0 1e-06 
0.0 1.0374 0 -2.0 1e-06 
0.0 1.0375 0 -2.0 1e-06 
0.0 1.0376 0 -2.0 1e-06 
0.0 1.0377 0 -2.0 1e-06 
0.0 1.0378 0 -2.0 1e-06 
0.0 1.0379 0 -2.0 1e-06 
0.0 1.038 0 -2.0 1e-06 
0.0 1.0381 0 -2.0 1e-06 
0.0 1.0382 0 -2.0 1e-06 
0.0 1.0383 0 -2.0 1e-06 
0.0 1.0384 0 -2.0 1e-06 
0.0 1.0385 0 -2.0 1e-06 
0.0 1.0386 0 -2.0 1e-06 
0.0 1.0387 0 -2.0 1e-06 
0.0 1.0388 0 -2.0 1e-06 
0.0 1.0389 0 -2.0 1e-06 
0.0 1.039 0 -2.0 1e-06 
0.0 1.0391 0 -2.0 1e-06 
0.0 1.0392 0 -2.0 1e-06 
0.0 1.0393 0 -2.0 1e-06 
0.0 1.0394 0 -2.0 1e-06 
0.0 1.0395 0 -2.0 1e-06 
0.0 1.0396 0 -2.0 1e-06 
0.0 1.0397 0 -2.0 1e-06 
0.0 1.0398 0 -2.0 1e-06 
0.0 1.0399 0 -2.0 1e-06 
0.0 1.04 0 -2.0 1e-06 
0.0 1.0401 0 -2.0 1e-06 
0.0 1.0402 0 -2.0 1e-06 
0.0 1.0403 0 -2.0 1e-06 
0.0 1.0404 0 -2.0 1e-06 
0.0 1.0405 0 -2.0 1e-06 
0.0 1.0406 0 -2.0 1e-06 
0.0 1.0407 0 -2.0 1e-06 
0.0 1.0408 0 -2.0 1e-06 
0.0 1.0409 0 -2.0 1e-06 
0.0 1.041 0 -2.0 1e-06 
0.0 1.0411 0 -2.0 1e-06 
0.0 1.0412 0 -2.0 1e-06 
0.0 1.0413 0 -2.0 1e-06 
0.0 1.0414 0 -2.0 1e-06 
0.0 1.0415 0 -2.0 1e-06 
0.0 1.0416 0 -2.0 1e-06 
0.0 1.0417 0 -2.0 1e-06 
0.0 1.0418 0 -2.0 1e-06 
0.0 1.0419 0 -2.0 1e-06 
0.0 1.042 0 -2.0 1e-06 
0.0 1.0421 0 -2.0 1e-06 
0.0 1.0422 0 -2.0 1e-06 
0.0 1.0423 0 -2.0 1e-06 
0.0 1.0424 0 -2.0 1e-06 
0.0 1.0425 0 -2.0 1e-06 
0.0 1.0426 0 -2.0 1e-06 
0.0 1.0427 0 -2.0 1e-06 
0.0 1.0428 0 -2.0 1e-06 
0.0 1.0429 0 -2.0 1e-06 
0.0 1.043 0 -2.0 1e-06 
0.0 1.0431 0 -2.0 1e-06 
0.0 1.0432 0 -2.0 1e-06 
0.0 1.0433 0 -2.0 1e-06 
0.0 1.0434 0 -2.0 1e-06 
0.0 1.0435 0 -2.0 1e-06 
0.0 1.0436 0 -2.0 1e-06 
0.0 1.0437 0 -2.0 1e-06 
0.0 1.0438 0 -2.0 1e-06 
0.0 1.0439 0 -2.0 1e-06 
0.0 1.044 0 -2.0 1e-06 
0.0 1.0441 0 -2.0 1e-06 
0.0 1.0442 0 -2.0 1e-06 
0.0 1.0443 0 -2.0 1e-06 
0.0 1.0444 0 -2.0 1e-06 
0.0 1.0445 0 -2.0 1e-06 
0.0 1.0446 0 -2.0 1e-06 
0.0 1.0447 0 -2.0 1e-06 
0.0 1.0448 0 -2.0 1e-06 
0.0 1.0449 0 -2.0 1e-06 
0.0 1.045 0 -2.0 1e-06 
0.0 1.0451 0 -2.0 1e-06 
0.0 1.0452 0 -2.0 1e-06 
0.0 1.0453 0 -2.0 1e-06 
0.0 1.0454 0 -2.0 1e-06 
0.0 1.0455 0 -2.0 1e-06 
0.0 1.0456 0 -2.0 1e-06 
0.0 1.0457 0 -2.0 1e-06 
0.0 1.0458 0 -2.0 1e-06 
0.0 1.0459 0 -2.0 1e-06 
0.0 1.046 0 -2.0 1e-06 
0.0 1.0461 0 -2.0 1e-06 
0.0 1.0462 0 -2.0 1e-06 
0.0 1.0463 0 -2.0 1e-06 
0.0 1.0464 0 -2.0 1e-06 
0.0 1.0465 0 -2.0 1e-06 
0.0 1.0466 0 -2.0 1e-06 
0.0 1.0467 0 -2.0 1e-06 
0.0 1.0468 0 -2.0 1e-06 
0.0 1.0469 0 -2.0 1e-06 
0.0 1.047 0 -2.0 1e-06 
0.0 1.0471 0 -2.0 1e-06 
0.0 1.0472 0 -2.0 1e-06 
0.0 1.0473 0 -2.0 1e-06 
0.0 1.0474 0 -2.0 1e-06 
0.0 1.0475 0 -2.0 1e-06 
0.0 1.0476 0 -2.0 1e-06 
0.0 1.0477 0 -2.0 1e-06 
0.0 1.0478 0 -2.0 1e-06 
0.0 1.0479 0 -2.0 1e-06 
0.0 1.048 0 -2.0 1e-06 
0.0 1.0481 0 -2.0 1e-06 
0.0 1.0482 0 -2.0 1e-06 
0.0 1.0483 0 -2.0 1e-06 
0.0 1.0484 0 -2.0 1e-06 
0.0 1.0485 0 -2.0 1e-06 
0.0 1.0486 0 -2.0 1e-06 
0.0 1.0487 0 -2.0 1e-06 
0.0 1.0488 0 -2.0 1e-06 
0.0 1.0489 0 -2.0 1e-06 
0.0 1.049 0 -2.0 1e-06 
0.0 1.0491 0 -2.0 1e-06 
0.0 1.0492 0 -2.0 1e-06 
0.0 1.0493 0 -2.0 1e-06 
0.0 1.0494 0 -2.0 1e-06 
0.0 1.0495 0 -2.0 1e-06 
0.0 1.0496 0 -2.0 1e-06 
0.0 1.0497 0 -2.0 1e-06 
0.0 1.0498 0 -2.0 1e-06 
0.0 1.0499 0 -2.0 1e-06 
0.0 1.05 0 -2.0 1e-06 
0.0 1.0501 0 -2.0 1e-06 
0.0 1.0502 0 -2.0 1e-06 
0.0 1.0503 0 -2.0 1e-06 
0.0 1.0504 0 -2.0 1e-06 
0.0 1.0505 0 -2.0 1e-06 
0.0 1.0506 0 -2.0 1e-06 
0.0 1.0507 0 -2.0 1e-06 
0.0 1.0508 0 -2.0 1e-06 
0.0 1.0509 0 -2.0 1e-06 
0.0 1.051 0 -2.0 1e-06 
0.0 1.0511 0 -2.0 1e-06 
0.0 1.0512 0 -2.0 1e-06 
0.0 1.0513 0 -2.0 1e-06 
0.0 1.0514 0 -2.0 1e-06 
0.0 1.0515 0 -2.0 1e-06 
0.0 1.0516 0 -2.0 1e-06 
0.0 1.0517 0 -2.0 1e-06 
0.0 1.0518 0 -2.0 1e-06 
0.0 1.0519 0 -2.0 1e-06 
0.0 1.052 0 -2.0 1e-06 
0.0 1.0521 0 -2.0 1e-06 
0.0 1.0522 0 -2.0 1e-06 
0.0 1.0523 0 -2.0 1e-06 
0.0 1.0524 0 -2.0 1e-06 
0.0 1.0525 0 -2.0 1e-06 
0.0 1.0526 0 -2.0 1e-06 
0.0 1.0527 0 -2.0 1e-06 
0.0 1.0528 0 -2.0 1e-06 
0.0 1.0529 0 -2.0 1e-06 
0.0 1.053 0 -2.0 1e-06 
0.0 1.0531 0 -2.0 1e-06 
0.0 1.0532 0 -2.0 1e-06 
0.0 1.0533 0 -2.0 1e-06 
0.0 1.0534 0 -2.0 1e-06 
0.0 1.0535 0 -2.0 1e-06 
0.0 1.0536 0 -2.0 1e-06 
0.0 1.0537 0 -2.0 1e-06 
0.0 1.0538 0 -2.0 1e-06 
0.0 1.0539 0 -2.0 1e-06 
0.0 1.054 0 -2.0 1e-06 
0.0 1.0541 0 -2.0 1e-06 
0.0 1.0542 0 -2.0 1e-06 
0.0 1.0543 0 -2.0 1e-06 
0.0 1.0544 0 -2.0 1e-06 
0.0 1.0545 0 -2.0 1e-06 
0.0 1.0546 0 -2.0 1e-06 
0.0 1.0547 0 -2.0 1e-06 
0.0 1.0548 0 -2.0 1e-06 
0.0 1.0549 0 -2.0 1e-06 
0.0 1.055 0 -2.0 1e-06 
0.0 1.0551 0 -2.0 1e-06 
0.0 1.0552 0 -2.0 1e-06 
0.0 1.0553 0 -2.0 1e-06 
0.0 1.0554 0 -2.0 1e-06 
0.0 1.0555 0 -2.0 1e-06 
0.0 1.0556 0 -2.0 1e-06 
0.0 1.0557 0 -2.0 1e-06 
0.0 1.0558 0 -2.0 1e-06 
0.0 1.0559 0 -2.0 1e-06 
0.0 1.056 0 -2.0 1e-06 
0.0 1.0561 0 -2.0 1e-06 
0.0 1.0562 0 -2.0 1e-06 
0.0 1.0563 0 -2.0 1e-06 
0.0 1.0564 0 -2.0 1e-06 
0.0 1.0565 0 -2.0 1e-06 
0.0 1.0566 0 -2.0 1e-06 
0.0 1.0567 0 -2.0 1e-06 
0.0 1.0568 0 -2.0 1e-06 
0.0 1.0569 0 -2.0 1e-06 
0.0 1.057 0 -2.0 1e-06 
0.0 1.0571 0 -2.0 1e-06 
0.0 1.0572 0 -2.0 1e-06 
0.0 1.0573 0 -2.0 1e-06 
0.0 1.0574 0 -2.0 1e-06 
0.0 1.0575 0 -2.0 1e-06 
0.0 1.0576 0 -2.0 1e-06 
0.0 1.0577 0 -2.0 1e-06 
0.0 1.0578 0 -2.0 1e-06 
0.0 1.0579 0 -2.0 1e-06 
0.0 1.058 0 -2.0 1e-06 
0.0 1.0581 0 -2.0 1e-06 
0.0 1.0582 0 -2.0 1e-06 
0.0 1.0583 0 -2.0 1e-06 
0.0 1.0584 0 -2.0 1e-06 
0.0 1.0585 0 -2.0 1e-06 
0.0 1.0586 0 -2.0 1e-06 
0.0 1.0587 0 -2.0 1e-06 
0.0 1.0588 0 -2.0 1e-06 
0.0 1.0589 0 -2.0 1e-06 
0.0 1.059 0 -2.0 1e-06 
0.0 1.0591 0 -2.0 1e-06 
0.0 1.0592 0 -2.0 1e-06 
0.0 1.0593 0 -2.0 1e-06 
0.0 1.0594 0 -2.0 1e-06 
0.0 1.0595 0 -2.0 1e-06 
0.0 1.0596 0 -2.0 1e-06 
0.0 1.0597 0 -2.0 1e-06 
0.0 1.0598 0 -2.0 1e-06 
0.0 1.0599 0 -2.0 1e-06 
0.0 1.06 0 -2.0 1e-06 
0.0 1.0601 0 -2.0 1e-06 
0.0 1.0602 0 -2.0 1e-06 
0.0 1.0603 0 -2.0 1e-06 
0.0 1.0604 0 -2.0 1e-06 
0.0 1.0605 0 -2.0 1e-06 
0.0 1.0606 0 -2.0 1e-06 
0.0 1.0607 0 -2.0 1e-06 
0.0 1.0608 0 -2.0 1e-06 
0.0 1.0609 0 -2.0 1e-06 
0.0 1.061 0 -2.0 1e-06 
0.0 1.0611 0 -2.0 1e-06 
0.0 1.0612 0 -2.0 1e-06 
0.0 1.0613 0 -2.0 1e-06 
0.0 1.0614 0 -2.0 1e-06 
0.0 1.0615 0 -2.0 1e-06 
0.0 1.0616 0 -2.0 1e-06 
0.0 1.0617 0 -2.0 1e-06 
0.0 1.0618 0 -2.0 1e-06 
0.0 1.0619 0 -2.0 1e-06 
0.0 1.062 0 -2.0 1e-06 
0.0 1.0621 0 -2.0 1e-06 
0.0 1.0622 0 -2.0 1e-06 
0.0 1.0623 0 -2.0 1e-06 
0.0 1.0624 0 -2.0 1e-06 
0.0 1.0625 0 -2.0 1e-06 
0.0 1.0626 0 -2.0 1e-06 
0.0 1.0627 0 -2.0 1e-06 
0.0 1.0628 0 -2.0 1e-06 
0.0 1.0629 0 -2.0 1e-06 
0.0 1.063 0 -2.0 1e-06 
0.0 1.0631 0 -2.0 1e-06 
0.0 1.0632 0 -2.0 1e-06 
0.0 1.0633 0 -2.0 1e-06 
0.0 1.0634 0 -2.0 1e-06 
0.0 1.0635 0 -2.0 1e-06 
0.0 1.0636 0 -2.0 1e-06 
0.0 1.0637 0 -2.0 1e-06 
0.0 1.0638 0 -2.0 1e-06 
0.0 1.0639 0 -2.0 1e-06 
0.0 1.064 0 -2.0 1e-06 
0.0 1.0641 0 -2.0 1e-06 
0.0 1.0642 0 -2.0 1e-06 
0.0 1.0643 0 -2.0 1e-06 
0.0 1.0644 0 -2.0 1e-06 
0.0 1.0645 0 -2.0 1e-06 
0.0 1.0646 0 -2.0 1e-06 
0.0 1.0647 0 -2.0 1e-06 
0.0 1.0648 0 -2.0 1e-06 
0.0 1.0649 0 -2.0 1e-06 
0.0 1.065 0 -2.0 1e-06 
0.0 1.0651 0 -2.0 1e-06 
0.0 1.0652 0 -2.0 1e-06 
0.0 1.0653 0 -2.0 1e-06 
0.0 1.0654 0 -2.0 1e-06 
0.0 1.0655 0 -2.0 1e-06 
0.0 1.0656 0 -2.0 1e-06 
0.0 1.0657 0 -2.0 1e-06 
0.0 1.0658 0 -2.0 1e-06 
0.0 1.0659 0 -2.0 1e-06 
0.0 1.066 0 -2.0 1e-06 
0.0 1.0661 0 -2.0 1e-06 
0.0 1.0662 0 -2.0 1e-06 
0.0 1.0663 0 -2.0 1e-06 
0.0 1.0664 0 -2.0 1e-06 
0.0 1.0665 0 -2.0 1e-06 
0.0 1.0666 0 -2.0 1e-06 
0.0 1.0667 0 -2.0 1e-06 
0.0 1.0668 0 -2.0 1e-06 
0.0 1.0669 0 -2.0 1e-06 
0.0 1.067 0 -2.0 1e-06 
0.0 1.0671 0 -2.0 1e-06 
0.0 1.0672 0 -2.0 1e-06 
0.0 1.0673 0 -2.0 1e-06 
0.0 1.0674 0 -2.0 1e-06 
0.0 1.0675 0 -2.0 1e-06 
0.0 1.0676 0 -2.0 1e-06 
0.0 1.0677 0 -2.0 1e-06 
0.0 1.0678 0 -2.0 1e-06 
0.0 1.0679 0 -2.0 1e-06 
0.0 1.068 0 -2.0 1e-06 
0.0 1.0681 0 -2.0 1e-06 
0.0 1.0682 0 -2.0 1e-06 
0.0 1.0683 0 -2.0 1e-06 
0.0 1.0684 0 -2.0 1e-06 
0.0 1.0685 0 -2.0 1e-06 
0.0 1.0686 0 -2.0 1e-06 
0.0 1.0687 0 -2.0 1e-06 
0.0 1.0688 0 -2.0 1e-06 
0.0 1.0689 0 -2.0 1e-06 
0.0 1.069 0 -2.0 1e-06 
0.0 1.0691 0 -2.0 1e-06 
0.0 1.0692 0 -2.0 1e-06 
0.0 1.0693 0 -2.0 1e-06 
0.0 1.0694 0 -2.0 1e-06 
0.0 1.0695 0 -2.0 1e-06 
0.0 1.0696 0 -2.0 1e-06 
0.0 1.0697 0 -2.0 1e-06 
0.0 1.0698 0 -2.0 1e-06 
0.0 1.0699 0 -2.0 1e-06 
0.0 1.07 0 -2.0 1e-06 
0.0 1.0701 0 -2.0 1e-06 
0.0 1.0702 0 -2.0 1e-06 
0.0 1.0703 0 -2.0 1e-06 
0.0 1.0704 0 -2.0 1e-06 
0.0 1.0705 0 -2.0 1e-06 
0.0 1.0706 0 -2.0 1e-06 
0.0 1.0707 0 -2.0 1e-06 
0.0 1.0708 0 -2.0 1e-06 
0.0 1.0709 0 -2.0 1e-06 
0.0 1.071 0 -2.0 1e-06 
0.0 1.0711 0 -2.0 1e-06 
0.0 1.0712 0 -2.0 1e-06 
0.0 1.0713 0 -2.0 1e-06 
0.0 1.0714 0 -2.0 1e-06 
0.0 1.0715 0 -2.0 1e-06 
0.0 1.0716 0 -2.0 1e-06 
0.0 1.0717 0 -2.0 1e-06 
0.0 1.0718 0 -2.0 1e-06 
0.0 1.0719 0 -2.0 1e-06 
0.0 1.072 0 -2.0 1e-06 
0.0 1.0721 0 -2.0 1e-06 
0.0 1.0722 0 -2.0 1e-06 
0.0 1.0723 0 -2.0 1e-06 
0.0 1.0724 0 -2.0 1e-06 
0.0 1.0725 0 -2.0 1e-06 
0.0 1.0726 0 -2.0 1e-06 
0.0 1.0727 0 -2.0 1e-06 
0.0 1.0728 0 -2.0 1e-06 
0.0 1.0729 0 -2.0 1e-06 
0.0 1.073 0 -2.0 1e-06 
0.0 1.0731 0 -2.0 1e-06 
0.0 1.0732 0 -2.0 1e-06 
0.0 1.0733 0 -2.0 1e-06 
0.0 1.0734 0 -2.0 1e-06 
0.0 1.0735 0 -2.0 1e-06 
0.0 1.0736 0 -2.0 1e-06 
0.0 1.0737 0 -2.0 1e-06 
0.0 1.0738 0 -2.0 1e-06 
0.0 1.0739 0 -2.0 1e-06 
0.0 1.074 0 -2.0 1e-06 
0.0 1.0741 0 -2.0 1e-06 
0.0 1.0742 0 -2.0 1e-06 
0.0 1.0743 0 -2.0 1e-06 
0.0 1.0744 0 -2.0 1e-06 
0.0 1.0745 0 -2.0 1e-06 
0.0 1.0746 0 -2.0 1e-06 
0.0 1.0747 0 -2.0 1e-06 
0.0 1.0748 0 -2.0 1e-06 
0.0 1.0749 0 -2.0 1e-06 
0.0 1.075 0 -2.0 1e-06 
0.0 1.0751 0 -2.0 1e-06 
0.0 1.0752 0 -2.0 1e-06 
0.0 1.0753 0 -2.0 1e-06 
0.0 1.0754 0 -2.0 1e-06 
0.0 1.0755 0 -2.0 1e-06 
0.0 1.0756 0 -2.0 1e-06 
0.0 1.0757 0 -2.0 1e-06 
0.0 1.0758 0 -2.0 1e-06 
0.0 1.0759 0 -2.0 1e-06 
0.0 1.076 0 -2.0 1e-06 
0.0 1.0761 0 -2.0 1e-06 
0.0 1.0762 0 -2.0 1e-06 
0.0 1.0763 0 -2.0 1e-06 
0.0 1.0764 0 -2.0 1e-06 
0.0 1.0765 0 -2.0 1e-06 
0.0 1.0766 0 -2.0 1e-06 
0.0 1.0767 0 -2.0 1e-06 
0.0 1.0768 0 -2.0 1e-06 
0.0 1.0769 0 -2.0 1e-06 
0.0 1.077 0 -2.0 1e-06 
0.0 1.0771 0 -2.0 1e-06 
0.0 1.0772 0 -2.0 1e-06 
0.0 1.0773 0 -2.0 1e-06 
0.0 1.0774 0 -2.0 1e-06 
0.0 1.0775 0 -2.0 1e-06 
0.0 1.0776 0 -2.0 1e-06 
0.0 1.0777 0 -2.0 1e-06 
0.0 1.0778 0 -2.0 1e-06 
0.0 1.0779 0 -2.0 1e-06 
0.0 1.078 0 -2.0 1e-06 
0.0 1.0781 0 -2.0 1e-06 
0.0 1.0782 0 -2.0 1e-06 
0.0 1.0783 0 -2.0 1e-06 
0.0 1.0784 0 -2.0 1e-06 
0.0 1.0785 0 -2.0 1e-06 
0.0 1.0786 0 -2.0 1e-06 
0.0 1.0787 0 -2.0 1e-06 
0.0 1.0788 0 -2.0 1e-06 
0.0 1.0789 0 -2.0 1e-06 
0.0 1.079 0 -2.0 1e-06 
0.0 1.0791 0 -2.0 1e-06 
0.0 1.0792 0 -2.0 1e-06 
0.0 1.0793 0 -2.0 1e-06 
0.0 1.0794 0 -2.0 1e-06 
0.0 1.0795 0 -2.0 1e-06 
0.0 1.0796 0 -2.0 1e-06 
0.0 1.0797 0 -2.0 1e-06 
0.0 1.0798 0 -2.0 1e-06 
0.0 1.0799 0 -2.0 1e-06 
0.0 1.08 0 -2.0 1e-06 
0.0 1.0801 0 -2.0 1e-06 
0.0 1.0802 0 -2.0 1e-06 
0.0 1.0803 0 -2.0 1e-06 
0.0 1.0804 0 -2.0 1e-06 
0.0 1.0805 0 -2.0 1e-06 
0.0 1.0806 0 -2.0 1e-06 
0.0 1.0807 0 -2.0 1e-06 
0.0 1.0808 0 -2.0 1e-06 
0.0 1.0809 0 -2.0 1e-06 
0.0 1.081 0 -2.0 1e-06 
0.0 1.0811 0 -2.0 1e-06 
0.0 1.0812 0 -2.0 1e-06 
0.0 1.0813 0 -2.0 1e-06 
0.0 1.0814 0 -2.0 1e-06 
0.0 1.0815 0 -2.0 1e-06 
0.0 1.0816 0 -2.0 1e-06 
0.0 1.0817 0 -2.0 1e-06 
0.0 1.0818 0 -2.0 1e-06 
0.0 1.0819 0 -2.0 1e-06 
0.0 1.082 0 -2.0 1e-06 
0.0 1.0821 0 -2.0 1e-06 
0.0 1.0822 0 -2.0 1e-06 
0.0 1.0823 0 -2.0 1e-06 
0.0 1.0824 0 -2.0 1e-06 
0.0 1.0825 0 -2.0 1e-06 
0.0 1.0826 0 -2.0 1e-06 
0.0 1.0827 0 -2.0 1e-06 
0.0 1.0828 0 -2.0 1e-06 
0.0 1.0829 0 -2.0 1e-06 
0.0 1.083 0 -2.0 1e-06 
0.0 1.0831 0 -2.0 1e-06 
0.0 1.0832 0 -2.0 1e-06 
0.0 1.0833 0 -2.0 1e-06 
0.0 1.0834 0 -2.0 1e-06 
0.0 1.0835 0 -2.0 1e-06 
0.0 1.0836 0 -2.0 1e-06 
0.0 1.0837 0 -2.0 1e-06 
0.0 1.0838 0 -2.0 1e-06 
0.0 1.0839 0 -2.0 1e-06 
0.0 1.084 0 -2.0 1e-06 
0.0 1.0841 0 -2.0 1e-06 
0.0 1.0842 0 -2.0 1e-06 
0.0 1.0843 0 -2.0 1e-06 
0.0 1.0844 0 -2.0 1e-06 
0.0 1.0845 0 -2.0 1e-06 
0.0 1.0846 0 -2.0 1e-06 
0.0 1.0847 0 -2.0 1e-06 
0.0 1.0848 0 -2.0 1e-06 
0.0 1.0849 0 -2.0 1e-06 
0.0 1.085 0 -2.0 1e-06 
0.0 1.0851 0 -2.0 1e-06 
0.0 1.0852 0 -2.0 1e-06 
0.0 1.0853 0 -2.0 1e-06 
0.0 1.0854 0 -2.0 1e-06 
0.0 1.0855 0 -2.0 1e-06 
0.0 1.0856 0 -2.0 1e-06 
0.0 1.0857 0 -2.0 1e-06 
0.0 1.0858 0 -2.0 1e-06 
0.0 1.0859 0 -2.0 1e-06 
0.0 1.086 0 -2.0 1e-06 
0.0 1.0861 0 -2.0 1e-06 
0.0 1.0862 0 -2.0 1e-06 
0.0 1.0863 0 -2.0 1e-06 
0.0 1.0864 0 -2.0 1e-06 
0.0 1.0865 0 -2.0 1e-06 
0.0 1.0866 0 -2.0 1e-06 
0.0 1.0867 0 -2.0 1e-06 
0.0 1.0868 0 -2.0 1e-06 
0.0 1.0869 0 -2.0 1e-06 
0.0 1.087 0 -2.0 1e-06 
0.0 1.0871 0 -2.0 1e-06 
0.0 1.0872 0 -2.0 1e-06 
0.0 1.0873 0 -2.0 1e-06 
0.0 1.0874 0 -2.0 1e-06 
0.0 1.0875 0 -2.0 1e-06 
0.0 1.0876 0 -2.0 1e-06 
0.0 1.0877 0 -2.0 1e-06 
0.0 1.0878 0 -2.0 1e-06 
0.0 1.0879 0 -2.0 1e-06 
0.0 1.088 0 -2.0 1e-06 
0.0 1.0881 0 -2.0 1e-06 
0.0 1.0882 0 -2.0 1e-06 
0.0 1.0883 0 -2.0 1e-06 
0.0 1.0884 0 -2.0 1e-06 
0.0 1.0885 0 -2.0 1e-06 
0.0 1.0886 0 -2.0 1e-06 
0.0 1.0887 0 -2.0 1e-06 
0.0 1.0888 0 -2.0 1e-06 
0.0 1.0889 0 -2.0 1e-06 
0.0 1.089 0 -2.0 1e-06 
0.0 1.0891 0 -2.0 1e-06 
0.0 1.0892 0 -2.0 1e-06 
0.0 1.0893 0 -2.0 1e-06 
0.0 1.0894 0 -2.0 1e-06 
0.0 1.0895 0 -2.0 1e-06 
0.0 1.0896 0 -2.0 1e-06 
0.0 1.0897 0 -2.0 1e-06 
0.0 1.0898 0 -2.0 1e-06 
0.0 1.0899 0 -2.0 1e-06 
0.0 1.09 0 -2.0 1e-06 
0.0 1.0901 0 -2.0 1e-06 
0.0 1.0902 0 -2.0 1e-06 
0.0 1.0903 0 -2.0 1e-06 
0.0 1.0904 0 -2.0 1e-06 
0.0 1.0905 0 -2.0 1e-06 
0.0 1.0906 0 -2.0 1e-06 
0.0 1.0907 0 -2.0 1e-06 
0.0 1.0908 0 -2.0 1e-06 
0.0 1.0909 0 -2.0 1e-06 
0.0 1.091 0 -2.0 1e-06 
0.0 1.0911 0 -2.0 1e-06 
0.0 1.0912 0 -2.0 1e-06 
0.0 1.0913 0 -2.0 1e-06 
0.0 1.0914 0 -2.0 1e-06 
0.0 1.0915 0 -2.0 1e-06 
0.0 1.0916 0 -2.0 1e-06 
0.0 1.0917 0 -2.0 1e-06 
0.0 1.0918 0 -2.0 1e-06 
0.0 1.0919 0 -2.0 1e-06 
0.0 1.092 0 -2.0 1e-06 
0.0 1.0921 0 -2.0 1e-06 
0.0 1.0922 0 -2.0 1e-06 
0.0 1.0923 0 -2.0 1e-06 
0.0 1.0924 0 -2.0 1e-06 
0.0 1.0925 0 -2.0 1e-06 
0.0 1.0926 0 -2.0 1e-06 
0.0 1.0927 0 -2.0 1e-06 
0.0 1.0928 0 -2.0 1e-06 
0.0 1.0929 0 -2.0 1e-06 
0.0 1.093 0 -2.0 1e-06 
0.0 1.0931 0 -2.0 1e-06 
0.0 1.0932 0 -2.0 1e-06 
0.0 1.0933 0 -2.0 1e-06 
0.0 1.0934 0 -2.0 1e-06 
0.0 1.0935 0 -2.0 1e-06 
0.0 1.0936 0 -2.0 1e-06 
0.0 1.0937 0 -2.0 1e-06 
0.0 1.0938 0 -2.0 1e-06 
0.0 1.0939 0 -2.0 1e-06 
0.0 1.094 0 -2.0 1e-06 
0.0 1.0941 0 -2.0 1e-06 
0.0 1.0942 0 -2.0 1e-06 
0.0 1.0943 0 -2.0 1e-06 
0.0 1.0944 0 -2.0 1e-06 
0.0 1.0945 0 -2.0 1e-06 
0.0 1.0946 0 -2.0 1e-06 
0.0 1.0947 0 -2.0 1e-06 
0.0 1.0948 0 -2.0 1e-06 
0.0 1.0949 0 -2.0 1e-06 
0.0 1.095 0 -2.0 1e-06 
0.0 1.0951 0 -2.0 1e-06 
0.0 1.0952 0 -2.0 1e-06 
0.0 1.0953 0 -2.0 1e-06 
0.0 1.0954 0 -2.0 1e-06 
0.0 1.0955 0 -2.0 1e-06 
0.0 1.0956 0 -2.0 1e-06 
0.0 1.0957 0 -2.0 1e-06 
0.0 1.0958 0 -2.0 1e-06 
0.0 1.0959 0 -2.0 1e-06 
0.0 1.096 0 -2.0 1e-06 
0.0 1.0961 0 -2.0 1e-06 
0.0 1.0962 0 -2.0 1e-06 
0.0 1.0963 0 -2.0 1e-06 
0.0 1.0964 0 -2.0 1e-06 
0.0 1.0965 0 -2.0 1e-06 
0.0 1.0966 0 -2.0 1e-06 
0.0 1.0967 0 -2.0 1e-06 
0.0 1.0968 0 -2.0 1e-06 
0.0 1.0969 0 -2.0 1e-06 
0.0 1.097 0 -2.0 1e-06 
0.0 1.0971 0 -2.0 1e-06 
0.0 1.0972 0 -2.0 1e-06 
0.0 1.0973 0 -2.0 1e-06 
0.0 1.0974 0 -2.0 1e-06 
0.0 1.0975 0 -2.0 1e-06 
0.0 1.0976 0 -2.0 1e-06 
0.0 1.0977 0 -2.0 1e-06 
0.0 1.0978 0 -2.0 1e-06 
0.0 1.0979 0 -2.0 1e-06 
0.0 1.098 0 -2.0 1e-06 
0.0 1.0981 0 -2.0 1e-06 
0.0 1.0982 0 -2.0 1e-06 
0.0 1.0983 0 -2.0 1e-06 
0.0 1.0984 0 -2.0 1e-06 
0.0 1.0985 0 -2.0 1e-06 
0.0 1.0986 0 -2.0 1e-06 
0.0 1.0987 0 -2.0 1e-06 
0.0 1.0988 0 -2.0 1e-06 
0.0 1.0989 0 -2.0 1e-06 
0.0 1.099 0 -2.0 1e-06 
0.0 1.0991 0 -2.0 1e-06 
0.0 1.0992 0 -2.0 1e-06 
0.0 1.0993 0 -2.0 1e-06 
0.0 1.0994 0 -2.0 1e-06 
0.0 1.0995 0 -2.0 1e-06 
0.0 1.0996 0 -2.0 1e-06 
0.0 1.0997 0 -2.0 1e-06 
0.0 1.0998 0 -2.0 1e-06 
0.0 1.0999 0 -2.0 1e-06 
0.0 1.1 0 -2.0 1e-06 
0.0 1.1001 0 -2.0 1e-06 
0.0 1.1002 0 -2.0 1e-06 
0.0 1.1003 0 -2.0 1e-06 
0.0 1.1004 0 -2.0 1e-06 
0.0 1.1005 0 -2.0 1e-06 
0.0 1.1006 0 -2.0 1e-06 
0.0 1.1007 0 -2.0 1e-06 
0.0 1.1008 0 -2.0 1e-06 
0.0 1.1009 0 -2.0 1e-06 
0.0 1.101 0 -2.0 1e-06 
0.0 1.1011 0 -2.0 1e-06 
0.0 1.1012 0 -2.0 1e-06 
0.0 1.1013 0 -2.0 1e-06 
0.0 1.1014 0 -2.0 1e-06 
0.0 1.1015 0 -2.0 1e-06 
0.0 1.1016 0 -2.0 1e-06 
0.0 1.1017 0 -2.0 1e-06 
0.0 1.1018 0 -2.0 1e-06 
0.0 1.1019 0 -2.0 1e-06 
0.0 1.102 0 -2.0 1e-06 
0.0 1.1021 0 -2.0 1e-06 
0.0 1.1022 0 -2.0 1e-06 
0.0 1.1023 0 -2.0 1e-06 
0.0 1.1024 0 -2.0 1e-06 
0.0 1.1025 0 -2.0 1e-06 
0.0 1.1026 0 -2.0 1e-06 
0.0 1.1027 0 -2.0 1e-06 
0.0 1.1028 0 -2.0 1e-06 
0.0 1.1029 0 -2.0 1e-06 
0.0 1.103 0 -2.0 1e-06 
0.0 1.1031 0 -2.0 1e-06 
0.0 1.1032 0 -2.0 1e-06 
0.0 1.1033 0 -2.0 1e-06 
0.0 1.1034 0 -2.0 1e-06 
0.0 1.1035 0 -2.0 1e-06 
0.0 1.1036 0 -2.0 1e-06 
0.0 1.1037 0 -2.0 1e-06 
0.0 1.1038 0 -2.0 1e-06 
0.0 1.1039 0 -2.0 1e-06 
0.0 1.104 0 -2.0 1e-06 
0.0 1.1041 0 -2.0 1e-06 
0.0 1.1042 0 -2.0 1e-06 
0.0 1.1043 0 -2.0 1e-06 
0.0 1.1044 0 -2.0 1e-06 
0.0 1.1045 0 -2.0 1e-06 
0.0 1.1046 0 -2.0 1e-06 
0.0 1.1047 0 -2.0 1e-06 
0.0 1.1048 0 -2.0 1e-06 
0.0 1.1049 0 -2.0 1e-06 
0.0 1.105 0 -2.0 1e-06 
0.0 1.1051 0 -2.0 1e-06 
0.0 1.1052 0 -2.0 1e-06 
0.0 1.1053 0 -2.0 1e-06 
0.0 1.1054 0 -2.0 1e-06 
0.0 1.1055 0 -2.0 1e-06 
0.0 1.1056 0 -2.0 1e-06 
0.0 1.1057 0 -2.0 1e-06 
0.0 1.1058 0 -2.0 1e-06 
0.0 1.1059 0 -2.0 1e-06 
0.0 1.106 0 -2.0 1e-06 
0.0 1.1061 0 -2.0 1e-06 
0.0 1.1062 0 -2.0 1e-06 
0.0 1.1063 0 -2.0 1e-06 
0.0 1.1064 0 -2.0 1e-06 
0.0 1.1065 0 -2.0 1e-06 
0.0 1.1066 0 -2.0 1e-06 
0.0 1.1067 0 -2.0 1e-06 
0.0 1.1068 0 -2.0 1e-06 
0.0 1.1069 0 -2.0 1e-06 
0.0 1.107 0 -2.0 1e-06 
0.0 1.1071 0 -2.0 1e-06 
0.0 1.1072 0 -2.0 1e-06 
0.0 1.1073 0 -2.0 1e-06 
0.0 1.1074 0 -2.0 1e-06 
0.0 1.1075 0 -2.0 1e-06 
0.0 1.1076 0 -2.0 1e-06 
0.0 1.1077 0 -2.0 1e-06 
0.0 1.1078 0 -2.0 1e-06 
0.0 1.1079 0 -2.0 1e-06 
0.0 1.108 0 -2.0 1e-06 
0.0 1.1081 0 -2.0 1e-06 
0.0 1.1082 0 -2.0 1e-06 
0.0 1.1083 0 -2.0 1e-06 
0.0 1.1084 0 -2.0 1e-06 
0.0 1.1085 0 -2.0 1e-06 
0.0 1.1086 0 -2.0 1e-06 
0.0 1.1087 0 -2.0 1e-06 
0.0 1.1088 0 -2.0 1e-06 
0.0 1.1089 0 -2.0 1e-06 
0.0 1.109 0 -2.0 1e-06 
0.0 1.1091 0 -2.0 1e-06 
0.0 1.1092 0 -2.0 1e-06 
0.0 1.1093 0 -2.0 1e-06 
0.0 1.1094 0 -2.0 1e-06 
0.0 1.1095 0 -2.0 1e-06 
0.0 1.1096 0 -2.0 1e-06 
0.0 1.1097 0 -2.0 1e-06 
0.0 1.1098 0 -2.0 1e-06 
0.0 1.1099 0 -2.0 1e-06 
0.0 1.11 0 -2.0 1e-06 
0.0 1.1101 0 -2.0 1e-06 
0.0 1.1102 0 -2.0 1e-06 
0.0 1.1103 0 -2.0 1e-06 
0.0 1.1104 0 -2.0 1e-06 
0.0 1.1105 0 -2.0 1e-06 
0.0 1.1106 0 -2.0 1e-06 
0.0 1.1107 0 -2.0 1e-06 
0.0 1.1108 0 -2.0 1e-06 
0.0 1.1109 0 -2.0 1e-06 
0.0 1.111 0 -2.0 1e-06 
0.0 1.1111 0 -2.0 1e-06 
0.0 1.1112 0 -2.0 1e-06 
0.0 1.1113 0 -2.0 1e-06 
0.0 1.1114 0 -2.0 1e-06 
0.0 1.1115 0 -2.0 1e-06 
0.0 1.1116 0 -2.0 1e-06 
0.0 1.1117 0 -2.0 1e-06 
0.0 1.1118 0 -2.0 1e-06 
0.0 1.1119 0 -2.0 1e-06 
0.0 1.112 0 -2.0 1e-06 
0.0 1.1121 0 -2.0 1e-06 
0.0 1.1122 0 -2.0 1e-06 
0.0 1.1123 0 -2.0 1e-06 
0.0 1.1124 0 -2.0 1e-06 
0.0 1.1125 0 -2.0 1e-06 
0.0 1.1126 0 -2.0 1e-06 
0.0 1.1127 0 -2.0 1e-06 
0.0 1.1128 0 -2.0 1e-06 
0.0 1.1129 0 -2.0 1e-06 
0.0 1.113 0 -2.0 1e-06 
0.0 1.1131 0 -2.0 1e-06 
0.0 1.1132 0 -2.0 1e-06 
0.0 1.1133 0 -2.0 1e-06 
0.0 1.1134 0 -2.0 1e-06 
0.0 1.1135 0 -2.0 1e-06 
0.0 1.1136 0 -2.0 1e-06 
0.0 1.1137 0 -2.0 1e-06 
0.0 1.1138 0 -2.0 1e-06 
0.0 1.1139 0 -2.0 1e-06 
0.0 1.114 0 -2.0 1e-06 
0.0 1.1141 0 -2.0 1e-06 
0.0 1.1142 0 -2.0 1e-06 
0.0 1.1143 0 -2.0 1e-06 
0.0 1.1144 0 -2.0 1e-06 
0.0 1.1145 0 -2.0 1e-06 
0.0 1.1146 0 -2.0 1e-06 
0.0 1.1147 0 -2.0 1e-06 
0.0 1.1148 0 -2.0 1e-06 
0.0 1.1149 0 -2.0 1e-06 
0.0 1.115 0 -2.0 1e-06 
0.0 1.1151 0 -2.0 1e-06 
0.0 1.1152 0 -2.0 1e-06 
0.0 1.1153 0 -2.0 1e-06 
0.0 1.1154 0 -2.0 1e-06 
0.0 1.1155 0 -2.0 1e-06 
0.0 1.1156 0 -2.0 1e-06 
0.0 1.1157 0 -2.0 1e-06 
0.0 1.1158 0 -2.0 1e-06 
0.0 1.1159 0 -2.0 1e-06 
0.0 1.116 0 -2.0 1e-06 
0.0 1.1161 0 -2.0 1e-06 
0.0 1.1162 0 -2.0 1e-06 
0.0 1.1163 0 -2.0 1e-06 
0.0 1.1164 0 -2.0 1e-06 
0.0 1.1165 0 -2.0 1e-06 
0.0 1.1166 0 -2.0 1e-06 
0.0 1.1167 0 -2.0 1e-06 
0.0 1.1168 0 -2.0 1e-06 
0.0 1.1169 0 -2.0 1e-06 
0.0 1.117 0 -2.0 1e-06 
0.0 1.1171 0 -2.0 1e-06 
0.0 1.1172 0 -2.0 1e-06 
0.0 1.1173 0 -2.0 1e-06 
0.0 1.1174 0 -2.0 1e-06 
0.0 1.1175 0 -2.0 1e-06 
0.0 1.1176 0 -2.0 1e-06 
0.0 1.1177 0 -2.0 1e-06 
0.0 1.1178 0 -2.0 1e-06 
0.0 1.1179 0 -2.0 1e-06 
0.0 1.118 0 -2.0 1e-06 
0.0 1.1181 0 -2.0 1e-06 
0.0 1.1182 0 -2.0 1e-06 
0.0 1.1183 0 -2.0 1e-06 
0.0 1.1184 0 -2.0 1e-06 
0.0 1.1185 0 -2.0 1e-06 
0.0 1.1186 0 -2.0 1e-06 
0.0 1.1187 0 -2.0 1e-06 
0.0 1.1188 0 -2.0 1e-06 
0.0 1.1189 0 -2.0 1e-06 
0.0 1.119 0 -2.0 1e-06 
0.0 1.1191 0 -2.0 1e-06 
0.0 1.1192 0 -2.0 1e-06 
0.0 1.1193 0 -2.0 1e-06 
0.0 1.1194 0 -2.0 1e-06 
0.0 1.1195 0 -2.0 1e-06 
0.0 1.1196 0 -2.0 1e-06 
0.0 1.1197 0 -2.0 1e-06 
0.0 1.1198 0 -2.0 1e-06 
0.0 1.1199 0 -2.0 1e-06 
0.0 1.12 0 -2.0 1e-06 
0.0 1.1201 0 -2.0 1e-06 
0.0 1.1202 0 -2.0 1e-06 
0.0 1.1203 0 -2.0 1e-06 
0.0 1.1204 0 -2.0 1e-06 
0.0 1.1205 0 -2.0 1e-06 
0.0 1.1206 0 -2.0 1e-06 
0.0 1.1207 0 -2.0 1e-06 
0.0 1.1208 0 -2.0 1e-06 
0.0 1.1209 0 -2.0 1e-06 
0.0 1.121 0 -2.0 1e-06 
0.0 1.1211 0 -2.0 1e-06 
0.0 1.1212 0 -2.0 1e-06 
0.0 1.1213 0 -2.0 1e-06 
0.0 1.1214 0 -2.0 1e-06 
0.0 1.1215 0 -2.0 1e-06 
0.0 1.1216 0 -2.0 1e-06 
0.0 1.1217 0 -2.0 1e-06 
0.0 1.1218 0 -2.0 1e-06 
0.0 1.1219 0 -2.0 1e-06 
0.0 1.122 0 -2.0 1e-06 
0.0 1.1221 0 -2.0 1e-06 
0.0 1.1222 0 -2.0 1e-06 
0.0 1.1223 0 -2.0 1e-06 
0.0 1.1224 0 -2.0 1e-06 
0.0 1.1225 0 -2.0 1e-06 
0.0 1.1226 0 -2.0 1e-06 
0.0 1.1227 0 -2.0 1e-06 
0.0 1.1228 0 -2.0 1e-06 
0.0 1.1229 0 -2.0 1e-06 
0.0 1.123 0 -2.0 1e-06 
0.0 1.1231 0 -2.0 1e-06 
0.0 1.1232 0 -2.0 1e-06 
0.0 1.1233 0 -2.0 1e-06 
0.0 1.1234 0 -2.0 1e-06 
0.0 1.1235 0 -2.0 1e-06 
0.0 1.1236 0 -2.0 1e-06 
0.0 1.1237 0 -2.0 1e-06 
0.0 1.1238 0 -2.0 1e-06 
0.0 1.1239 0 -2.0 1e-06 
0.0 1.124 0 -2.0 1e-06 
0.0 1.1241 0 -2.0 1e-06 
0.0 1.1242 0 -2.0 1e-06 
0.0 1.1243 0 -2.0 1e-06 
0.0 1.1244 0 -2.0 1e-06 
0.0 1.1245 0 -2.0 1e-06 
0.0 1.1246 0 -2.0 1e-06 
0.0 1.1247 0 -2.0 1e-06 
0.0 1.1248 0 -2.0 1e-06 
0.0 1.1249 0 -2.0 1e-06 
0.0 1.125 0 -2.0 1e-06 
0.0 1.1251 0 -2.0 1e-06 
0.0 1.1252 0 -2.0 1e-06 
0.0 1.1253 0 -2.0 1e-06 
0.0 1.1254 0 -2.0 1e-06 
0.0 1.1255 0 -2.0 1e-06 
0.0 1.1256 0 -2.0 1e-06 
0.0 1.1257 0 -2.0 1e-06 
0.0 1.1258 0 -2.0 1e-06 
0.0 1.1259 0 -2.0 1e-06 
0.0 1.126 0 -2.0 1e-06 
0.0 1.1261 0 -2.0 1e-06 
0.0 1.1262 0 -2.0 1e-06 
0.0 1.1263 0 -2.0 1e-06 
0.0 1.1264 0 -2.0 1e-06 
0.0 1.1265 0 -2.0 1e-06 
0.0 1.1266 0 -2.0 1e-06 
0.0 1.1267 0 -2.0 1e-06 
0.0 1.1268 0 -2.0 1e-06 
0.0 1.1269 0 -2.0 1e-06 
0.0 1.127 0 -2.0 1e-06 
0.0 1.1271 0 -2.0 1e-06 
0.0 1.1272 0 -2.0 1e-06 
0.0 1.1273 0 -2.0 1e-06 
0.0 1.1274 0 -2.0 1e-06 
0.0 1.1275 0 -2.0 1e-06 
0.0 1.1276 0 -2.0 1e-06 
0.0 1.1277 0 -2.0 1e-06 
0.0 1.1278 0 -2.0 1e-06 
0.0 1.1279 0 -2.0 1e-06 
0.0 1.128 0 -2.0 1e-06 
0.0 1.1281 0 -2.0 1e-06 
0.0 1.1282 0 -2.0 1e-06 
0.0 1.1283 0 -2.0 1e-06 
0.0 1.1284 0 -2.0 1e-06 
0.0 1.1285 0 -2.0 1e-06 
0.0 1.1286 0 -2.0 1e-06 
0.0 1.1287 0 -2.0 1e-06 
0.0 1.1288 0 -2.0 1e-06 
0.0 1.1289 0 -2.0 1e-06 
0.0 1.129 0 -2.0 1e-06 
0.0 1.1291 0 -2.0 1e-06 
0.0 1.1292 0 -2.0 1e-06 
0.0 1.1293 0 -2.0 1e-06 
0.0 1.1294 0 -2.0 1e-06 
0.0 1.1295 0 -2.0 1e-06 
0.0 1.1296 0 -2.0 1e-06 
0.0 1.1297 0 -2.0 1e-06 
0.0 1.1298 0 -2.0 1e-06 
0.0 1.1299 0 -2.0 1e-06 
0.0 1.13 0 -2.0 1e-06 
0.0 1.1301 0 -2.0 1e-06 
0.0 1.1302 0 -2.0 1e-06 
0.0 1.1303 0 -2.0 1e-06 
0.0 1.1304 0 -2.0 1e-06 
0.0 1.1305 0 -2.0 1e-06 
0.0 1.1306 0 -2.0 1e-06 
0.0 1.1307 0 -2.0 1e-06 
0.0 1.1308 0 -2.0 1e-06 
0.0 1.1309 0 -2.0 1e-06 
0.0 1.131 0 -2.0 1e-06 
0.0 1.1311 0 -2.0 1e-06 
0.0 1.1312 0 -2.0 1e-06 
0.0 1.1313 0 -2.0 1e-06 
0.0 1.1314 0 -2.0 1e-06 
0.0 1.1315 0 -2.0 1e-06 
0.0 1.1316 0 -2.0 1e-06 
0.0 1.1317 0 -2.0 1e-06 
0.0 1.1318 0 -2.0 1e-06 
0.0 1.1319 0 -2.0 1e-06 
0.0 1.132 0 -2.0 1e-06 
0.0 1.1321 0 -2.0 1e-06 
0.0 1.1322 0 -2.0 1e-06 
0.0 1.1323 0 -2.0 1e-06 
0.0 1.1324 0 -2.0 1e-06 
0.0 1.1325 0 -2.0 1e-06 
0.0 1.1326 0 -2.0 1e-06 
0.0 1.1327 0 -2.0 1e-06 
0.0 1.1328 0 -2.0 1e-06 
0.0 1.1329 0 -2.0 1e-06 
0.0 1.133 0 -2.0 1e-06 
0.0 1.1331 0 -2.0 1e-06 
0.0 1.1332 0 -2.0 1e-06 
0.0 1.1333 0 -2.0 1e-06 
0.0 1.1334 0 -2.0 1e-06 
0.0 1.1335 0 -2.0 1e-06 
0.0 1.1336 0 -2.0 1e-06 
0.0 1.1337 0 -2.0 1e-06 
0.0 1.1338 0 -2.0 1e-06 
0.0 1.1339 0 -2.0 1e-06 
0.0 1.134 0 -2.0 1e-06 
0.0 1.1341 0 -2.0 1e-06 
0.0 1.1342 0 -2.0 1e-06 
0.0 1.1343 0 -2.0 1e-06 
0.0 1.1344 0 -2.0 1e-06 
0.0 1.1345 0 -2.0 1e-06 
0.0 1.1346 0 -2.0 1e-06 
0.0 1.1347 0 -2.0 1e-06 
0.0 1.1348 0 -2.0 1e-06 
0.0 1.1349 0 -2.0 1e-06 
0.0 1.135 0 -2.0 1e-06 
0.0 1.1351 0 -2.0 1e-06 
0.0 1.1352 0 -2.0 1e-06 
0.0 1.1353 0 -2.0 1e-06 
0.0 1.1354 0 -2.0 1e-06 
0.0 1.1355 0 -2.0 1e-06 
0.0 1.1356 0 -2.0 1e-06 
0.0 1.1357 0 -2.0 1e-06 
0.0 1.1358 0 -2.0 1e-06 
0.0 1.1359 0 -2.0 1e-06 
0.0 1.136 0 -2.0 1e-06 
0.0 1.1361 0 -2.0 1e-06 
0.0 1.1362 0 -2.0 1e-06 
0.0 1.1363 0 -2.0 1e-06 
0.0 1.1364 0 -2.0 1e-06 
0.0 1.1365 0 -2.0 1e-06 
0.0 1.1366 0 -2.0 1e-06 
0.0 1.1367 0 -2.0 1e-06 
0.0 1.1368 0 -2.0 1e-06 
0.0 1.1369 0 -2.0 1e-06 
0.0 1.137 0 -2.0 1e-06 
0.0 1.1371 0 -2.0 1e-06 
0.0 1.1372 0 -2.0 1e-06 
0.0 1.1373 0 -2.0 1e-06 
0.0 1.1374 0 -2.0 1e-06 
0.0 1.1375 0 -2.0 1e-06 
0.0 1.1376 0 -2.0 1e-06 
0.0 1.1377 0 -2.0 1e-06 
0.0 1.1378 0 -2.0 1e-06 
0.0 1.1379 0 -2.0 1e-06 
0.0 1.138 0 -2.0 1e-06 
0.0 1.1381 0 -2.0 1e-06 
0.0 1.1382 0 -2.0 1e-06 
0.0 1.1383 0 -2.0 1e-06 
0.0 1.1384 0 -2.0 1e-06 
0.0 1.1385 0 -2.0 1e-06 
0.0 1.1386 0 -2.0 1e-06 
0.0 1.1387 0 -2.0 1e-06 
0.0 1.1388 0 -2.0 1e-06 
0.0 1.1389 0 -2.0 1e-06 
0.0 1.139 0 -2.0 1e-06 
0.0 1.1391 0 -2.0 1e-06 
0.0 1.1392 0 -2.0 1e-06 
0.0 1.1393 0 -2.0 1e-06 
0.0 1.1394 0 -2.0 1e-06 
0.0 1.1395 0 -2.0 1e-06 
0.0 1.1396 0 -2.0 1e-06 
0.0 1.1397 0 -2.0 1e-06 
0.0 1.1398 0 -2.0 1e-06 
0.0 1.1399 0 -2.0 1e-06 
0.0 1.14 0 -2.0 1e-06 
0.0 1.1401 0 -2.0 1e-06 
0.0 1.1402 0 -2.0 1e-06 
0.0 1.1403 0 -2.0 1e-06 
0.0 1.1404 0 -2.0 1e-06 
0.0 1.1405 0 -2.0 1e-06 
0.0 1.1406 0 -2.0 1e-06 
0.0 1.1407 0 -2.0 1e-06 
0.0 1.1408 0 -2.0 1e-06 
0.0 1.1409 0 -2.0 1e-06 
0.0 1.141 0 -2.0 1e-06 
0.0 1.1411 0 -2.0 1e-06 
0.0 1.1412 0 -2.0 1e-06 
0.0 1.1413 0 -2.0 1e-06 
0.0 1.1414 0 -2.0 1e-06 
0.0 1.1415 0 -2.0 1e-06 
0.0 1.1416 0 -2.0 1e-06 
0.0 1.1417 0 -2.0 1e-06 
0.0 1.1418 0 -2.0 1e-06 
0.0 1.1419 0 -2.0 1e-06 
0.0 1.142 0 -2.0 1e-06 
0.0 1.1421 0 -2.0 1e-06 
0.0 1.1422 0 -2.0 1e-06 
0.0 1.1423 0 -2.0 1e-06 
0.0 1.1424 0 -2.0 1e-06 
0.0 1.1425 0 -2.0 1e-06 
0.0 1.1426 0 -2.0 1e-06 
0.0 1.1427 0 -2.0 1e-06 
0.0 1.1428 0 -2.0 1e-06 
0.0 1.1429 0 -2.0 1e-06 
0.0 1.143 0 -2.0 1e-06 
0.0 1.1431 0 -2.0 1e-06 
0.0 1.1432 0 -2.0 1e-06 
0.0 1.1433 0 -2.0 1e-06 
0.0 1.1434 0 -2.0 1e-06 
0.0 1.1435 0 -2.0 1e-06 
0.0 1.1436 0 -2.0 1e-06 
0.0 1.1437 0 -2.0 1e-06 
0.0 1.1438 0 -2.0 1e-06 
0.0 1.1439 0 -2.0 1e-06 
0.0 1.144 0 -2.0 1e-06 
0.0 1.1441 0 -2.0 1e-06 
0.0 1.1442 0 -2.0 1e-06 
0.0 1.1443 0 -2.0 1e-06 
0.0 1.1444 0 -2.0 1e-06 
0.0 1.1445 0 -2.0 1e-06 
0.0 1.1446 0 -2.0 1e-06 
0.0 1.1447 0 -2.0 1e-06 
0.0 1.1448 0 -2.0 1e-06 
0.0 1.1449 0 -2.0 1e-06 
0.0 1.145 0 -2.0 1e-06 
0.0 1.1451 0 -2.0 1e-06 
0.0 1.1452 0 -2.0 1e-06 
0.0 1.1453 0 -2.0 1e-06 
0.0 1.1454 0 -2.0 1e-06 
0.0 1.1455 0 -2.0 1e-06 
0.0 1.1456 0 -2.0 1e-06 
0.0 1.1457 0 -2.0 1e-06 
0.0 1.1458 0 -2.0 1e-06 
0.0 1.1459 0 -2.0 1e-06 
0.0 1.146 0 -2.0 1e-06 
0.0 1.1461 0 -2.0 1e-06 
0.0 1.1462 0 -2.0 1e-06 
0.0 1.1463 0 -2.0 1e-06 
0.0 1.1464 0 -2.0 1e-06 
0.0 1.1465 0 -2.0 1e-06 
0.0 1.1466 0 -2.0 1e-06 
0.0 1.1467 0 -2.0 1e-06 
0.0 1.1468 0 -2.0 1e-06 
0.0 1.1469 0 -2.0 1e-06 
0.0 1.147 0 -2.0 1e-06 
0.0 1.1471 0 -2.0 1e-06 
0.0 1.1472 0 -2.0 1e-06 
0.0 1.1473 0 -2.0 1e-06 
0.0 1.1474 0 -2.0 1e-06 
0.0 1.1475 0 -2.0 1e-06 
0.0 1.1476 0 -2.0 1e-06 
0.0 1.1477 0 -2.0 1e-06 
0.0 1.1478 0 -2.0 1e-06 
0.0 1.1479 0 -2.0 1e-06 
0.0 1.148 0 -2.0 1e-06 
0.0 1.1481 0 -2.0 1e-06 
0.0 1.1482 0 -2.0 1e-06 
0.0 1.1483 0 -2.0 1e-06 
0.0 1.1484 0 -2.0 1e-06 
0.0 1.1485 0 -2.0 1e-06 
0.0 1.1486 0 -2.0 1e-06 
0.0 1.1487 0 -2.0 1e-06 
0.0 1.1488 0 -2.0 1e-06 
0.0 1.1489 0 -2.0 1e-06 
0.0 1.149 0 -2.0 1e-06 
0.0 1.1491 0 -2.0 1e-06 
0.0 1.1492 0 -2.0 1e-06 
0.0 1.1493 0 -2.0 1e-06 
0.0 1.1494 0 -2.0 1e-06 
0.0 1.1495 0 -2.0 1e-06 
0.0 1.1496 0 -2.0 1e-06 
0.0 1.1497 0 -2.0 1e-06 
0.0 1.1498 0 -2.0 1e-06 
0.0 1.1499 0 -2.0 1e-06 
0.0 1.15 0 -2.0 1e-06 
0.0 1.1501 0 -2.0 1e-06 
0.0 1.1502 0 -2.0 1e-06 
0.0 1.1503 0 -2.0 1e-06 
0.0 1.1504 0 -2.0 1e-06 
0.0 1.1505 0 -2.0 1e-06 
0.0 1.1506 0 -2.0 1e-06 
0.0 1.1507 0 -2.0 1e-06 
0.0 1.1508 0 -2.0 1e-06 
0.0 1.1509 0 -2.0 1e-06 
0.0 1.151 0 -2.0 1e-06 
0.0 1.1511 0 -2.0 1e-06 
0.0 1.1512 0 -2.0 1e-06 
0.0 1.1513 0 -2.0 1e-06 
0.0 1.1514 0 -2.0 1e-06 
0.0 1.1515 0 -2.0 1e-06 
0.0 1.1516 0 -2.0 1e-06 
0.0 1.1517 0 -2.0 1e-06 
0.0 1.1518 0 -2.0 1e-06 
0.0 1.1519 0 -2.0 1e-06 
0.0 1.152 0 -2.0 1e-06 
0.0 1.1521 0 -2.0 1e-06 
0.0 1.1522 0 -2.0 1e-06 
0.0 1.1523 0 -2.0 1e-06 
0.0 1.1524 0 -2.0 1e-06 
0.0 1.1525 0 -2.0 1e-06 
0.0 1.1526 0 -2.0 1e-06 
0.0 1.1527 0 -2.0 1e-06 
0.0 1.1528 0 -2.0 1e-06 
0.0 1.1529 0 -2.0 1e-06 
0.0 1.153 0 -2.0 1e-06 
0.0 1.1531 0 -2.0 1e-06 
0.0 1.1532 0 -2.0 1e-06 
0.0 1.1533 0 -2.0 1e-06 
0.0 1.1534 0 -2.0 1e-06 
0.0 1.1535 0 -2.0 1e-06 
0.0 1.1536 0 -2.0 1e-06 
0.0 1.1537 0 -2.0 1e-06 
0.0 1.1538 0 -2.0 1e-06 
0.0 1.1539 0 -2.0 1e-06 
0.0 1.154 0 -2.0 1e-06 
0.0 1.1541 0 -2.0 1e-06 
0.0 1.1542 0 -2.0 1e-06 
0.0 1.1543 0 -2.0 1e-06 
0.0 1.1544 0 -2.0 1e-06 
0.0 1.1545 0 -2.0 1e-06 
0.0 1.1546 0 -2.0 1e-06 
0.0 1.1547 0 -2.0 1e-06 
0.0 1.1548 0 -2.0 1e-06 
0.0 1.1549 0 -2.0 1e-06 
0.0 1.155 0 -2.0 1e-06 
0.0 1.1551 0 -2.0 1e-06 
0.0 1.1552 0 -2.0 1e-06 
0.0 1.1553 0 -2.0 1e-06 
0.0 1.1554 0 -2.0 1e-06 
0.0 1.1555 0 -2.0 1e-06 
0.0 1.1556 0 -2.0 1e-06 
0.0 1.1557 0 -2.0 1e-06 
0.0 1.1558 0 -2.0 1e-06 
0.0 1.1559 0 -2.0 1e-06 
0.0 1.156 0 -2.0 1e-06 
0.0 1.1561 0 -2.0 1e-06 
0.0 1.1562 0 -2.0 1e-06 
0.0 1.1563 0 -2.0 1e-06 
0.0 1.1564 0 -2.0 1e-06 
0.0 1.1565 0 -2.0 1e-06 
0.0 1.1566 0 -2.0 1e-06 
0.0 1.1567 0 -2.0 1e-06 
0.0 1.1568 0 -2.0 1e-06 
0.0 1.1569 0 -2.0 1e-06 
0.0 1.157 0 -2.0 1e-06 
0.0 1.1571 0 -2.0 1e-06 
0.0 1.1572 0 -2.0 1e-06 
0.0 1.1573 0 -2.0 1e-06 
0.0 1.1574 0 -2.0 1e-06 
0.0 1.1575 0 -2.0 1e-06 
0.0 1.1576 0 -2.0 1e-06 
0.0 1.1577 0 -2.0 1e-06 
0.0 1.1578 0 -2.0 1e-06 
0.0 1.1579 0 -2.0 1e-06 
0.0 1.158 0 -2.0 1e-06 
0.0 1.1581 0 -2.0 1e-06 
0.0 1.1582 0 -2.0 1e-06 
0.0 1.1583 0 -2.0 1e-06 
0.0 1.1584 0 -2.0 1e-06 
0.0 1.1585 0 -2.0 1e-06 
0.0 1.1586 0 -2.0 1e-06 
0.0 1.1587 0 -2.0 1e-06 
0.0 1.1588 0 -2.0 1e-06 
0.0 1.1589 0 -2.0 1e-06 
0.0 1.159 0 -2.0 1e-06 
0.0 1.1591 0 -2.0 1e-06 
0.0 1.1592 0 -2.0 1e-06 
0.0 1.1593 0 -2.0 1e-06 
0.0 1.1594 0 -2.0 1e-06 
0.0 1.1595 0 -2.0 1e-06 
0.0 1.1596 0 -2.0 1e-06 
0.0 1.1597 0 -2.0 1e-06 
0.0 1.1598 0 -2.0 1e-06 
0.0 1.1599 0 -2.0 1e-06 
0.0 1.16 0 -2.0 1e-06 
0.0 1.1601 0 -2.0 1e-06 
0.0 1.1602 0 -2.0 1e-06 
0.0 1.1603 0 -2.0 1e-06 
0.0 1.1604 0 -2.0 1e-06 
0.0 1.1605 0 -2.0 1e-06 
0.0 1.1606 0 -2.0 1e-06 
0.0 1.1607 0 -2.0 1e-06 
0.0 1.1608 0 -2.0 1e-06 
0.0 1.1609 0 -2.0 1e-06 
0.0 1.161 0 -2.0 1e-06 
0.0 1.1611 0 -2.0 1e-06 
0.0 1.1612 0 -2.0 1e-06 
0.0 1.1613 0 -2.0 1e-06 
0.0 1.1614 0 -2.0 1e-06 
0.0 1.1615 0 -2.0 1e-06 
0.0 1.1616 0 -2.0 1e-06 
0.0 1.1617 0 -2.0 1e-06 
0.0 1.1618 0 -2.0 1e-06 
0.0 1.1619 0 -2.0 1e-06 
0.0 1.162 0 -2.0 1e-06 
0.0 1.1621 0 -2.0 1e-06 
0.0 1.1622 0 -2.0 1e-06 
0.0 1.1623 0 -2.0 1e-06 
0.0 1.1624 0 -2.0 1e-06 
0.0 1.1625 0 -2.0 1e-06 
0.0 1.1626 0 -2.0 1e-06 
0.0 1.1627 0 -2.0 1e-06 
0.0 1.1628 0 -2.0 1e-06 
0.0 1.1629 0 -2.0 1e-06 
0.0 1.163 0 -2.0 1e-06 
0.0 1.1631 0 -2.0 1e-06 
0.0 1.1632 0 -2.0 1e-06 
0.0 1.1633 0 -2.0 1e-06 
0.0 1.1634 0 -2.0 1e-06 
0.0 1.1635 0 -2.0 1e-06 
0.0 1.1636 0 -2.0 1e-06 
0.0 1.1637 0 -2.0 1e-06 
0.0 1.1638 0 -2.0 1e-06 
0.0 1.1639 0 -2.0 1e-06 
0.0 1.164 0 -2.0 1e-06 
0.0 1.1641 0 -2.0 1e-06 
0.0 1.1642 0 -2.0 1e-06 
0.0 1.1643 0 -2.0 1e-06 
0.0 1.1644 0 -2.0 1e-06 
0.0 1.1645 0 -2.0 1e-06 
0.0 1.1646 0 -2.0 1e-06 
0.0 1.1647 0 -2.0 1e-06 
0.0 1.1648 0 -2.0 1e-06 
0.0 1.1649 0 -2.0 1e-06 
0.0 1.165 0 -2.0 1e-06 
0.0 1.1651 0 -2.0 1e-06 
0.0 1.1652 0 -2.0 1e-06 
0.0 1.1653 0 -2.0 1e-06 
0.0 1.1654 0 -2.0 1e-06 
0.0 1.1655 0 -2.0 1e-06 
0.0 1.1656 0 -2.0 1e-06 
0.0 1.1657 0 -2.0 1e-06 
0.0 1.1658 0 -2.0 1e-06 
0.0 1.1659 0 -2.0 1e-06 
0.0 1.166 0 -2.0 1e-06 
0.0 1.1661 0 -2.0 1e-06 
0.0 1.1662 0 -2.0 1e-06 
0.0 1.1663 0 -2.0 1e-06 
0.0 1.1664 0 -2.0 1e-06 
0.0 1.1665 0 -2.0 1e-06 
0.0 1.1666 0 -2.0 1e-06 
0.0 1.1667 0 -2.0 1e-06 
0.0 1.1668 0 -2.0 1e-06 
0.0 1.1669 0 -2.0 1e-06 
0.0 1.167 0 -2.0 1e-06 
0.0 1.1671 0 -2.0 1e-06 
0.0 1.1672 0 -2.0 1e-06 
0.0 1.1673 0 -2.0 1e-06 
0.0 1.1674 0 -2.0 1e-06 
0.0 1.1675 0 -2.0 1e-06 
0.0 1.1676 0 -2.0 1e-06 
0.0 1.1677 0 -2.0 1e-06 
0.0 1.1678 0 -2.0 1e-06 
0.0 1.1679 0 -2.0 1e-06 
0.0 1.168 0 -2.0 1e-06 
0.0 1.1681 0 -2.0 1e-06 
0.0 1.1682 0 -2.0 1e-06 
0.0 1.1683 0 -2.0 1e-06 
0.0 1.1684 0 -2.0 1e-06 
0.0 1.1685 0 -2.0 1e-06 
0.0 1.1686 0 -2.0 1e-06 
0.0 1.1687 0 -2.0 1e-06 
0.0 1.1688 0 -2.0 1e-06 
0.0 1.1689 0 -2.0 1e-06 
0.0 1.169 0 -2.0 1e-06 
0.0 1.1691 0 -2.0 1e-06 
0.0 1.1692 0 -2.0 1e-06 
0.0 1.1693 0 -2.0 1e-06 
0.0 1.1694 0 -2.0 1e-06 
0.0 1.1695 0 -2.0 1e-06 
0.0 1.1696 0 -2.0 1e-06 
0.0 1.1697 0 -2.0 1e-06 
0.0 1.1698 0 -2.0 1e-06 
0.0 1.1699 0 -2.0 1e-06 
0.0 1.17 0 -2.0 1e-06 
0.0 1.1701 0 -2.0 1e-06 
0.0 1.1702 0 -2.0 1e-06 
0.0 1.1703 0 -2.0 1e-06 
0.0 1.1704 0 -2.0 1e-06 
0.0 1.1705 0 -2.0 1e-06 
0.0 1.1706 0 -2.0 1e-06 
0.0 1.1707 0 -2.0 1e-06 
0.0 1.1708 0 -2.0 1e-06 
0.0 1.1709 0 -2.0 1e-06 
0.0 1.171 0 -2.0 1e-06 
0.0 1.1711 0 -2.0 1e-06 
0.0 1.1712 0 -2.0 1e-06 
0.0 1.1713 0 -2.0 1e-06 
0.0 1.1714 0 -2.0 1e-06 
0.0 1.1715 0 -2.0 1e-06 
0.0 1.1716 0 -2.0 1e-06 
0.0 1.1717 0 -2.0 1e-06 
0.0 1.1718 0 -2.0 1e-06 
0.0 1.1719 0 -2.0 1e-06 
0.0 1.172 0 -2.0 1e-06 
0.0 1.1721 0 -2.0 1e-06 
0.0 1.1722 0 -2.0 1e-06 
0.0 1.1723 0 -2.0 1e-06 
0.0 1.1724 0 -2.0 1e-06 
0.0 1.1725 0 -2.0 1e-06 
0.0 1.1726 0 -2.0 1e-06 
0.0 1.1727 0 -2.0 1e-06 
0.0 1.1728 0 -2.0 1e-06 
0.0 1.1729 0 -2.0 1e-06 
0.0 1.173 0 -2.0 1e-06 
0.0 1.1731 0 -2.0 1e-06 
0.0 1.1732 0 -2.0 1e-06 
0.0 1.1733 0 -2.0 1e-06 
0.0 1.1734 0 -2.0 1e-06 
0.0 1.1735 0 -2.0 1e-06 
0.0 1.1736 0 -2.0 1e-06 
0.0 1.1737 0 -2.0 1e-06 
0.0 1.1738 0 -2.0 1e-06 
0.0 1.1739 0 -2.0 1e-06 
0.0 1.174 0 -2.0 1e-06 
0.0 1.1741 0 -2.0 1e-06 
0.0 1.1742 0 -2.0 1e-06 
0.0 1.1743 0 -2.0 1e-06 
0.0 1.1744 0 -2.0 1e-06 
0.0 1.1745 0 -2.0 1e-06 
0.0 1.1746 0 -2.0 1e-06 
0.0 1.1747 0 -2.0 1e-06 
0.0 1.1748 0 -2.0 1e-06 
0.0 1.1749 0 -2.0 1e-06 
0.0 1.175 0 -2.0 1e-06 
0.0 1.1751 0 -2.0 1e-06 
0.0 1.1752 0 -2.0 1e-06 
0.0 1.1753 0 -2.0 1e-06 
0.0 1.1754 0 -2.0 1e-06 
0.0 1.1755 0 -2.0 1e-06 
0.0 1.1756 0 -2.0 1e-06 
0.0 1.1757 0 -2.0 1e-06 
0.0 1.1758 0 -2.0 1e-06 
0.0 1.1759 0 -2.0 1e-06 
0.0 1.176 0 -2.0 1e-06 
0.0 1.1761 0 -2.0 1e-06 
0.0 1.1762 0 -2.0 1e-06 
0.0 1.1763 0 -2.0 1e-06 
0.0 1.1764 0 -2.0 1e-06 
0.0 1.1765 0 -2.0 1e-06 
0.0 1.1766 0 -2.0 1e-06 
0.0 1.1767 0 -2.0 1e-06 
0.0 1.1768 0 -2.0 1e-06 
0.0 1.1769 0 -2.0 1e-06 
0.0 1.177 0 -2.0 1e-06 
0.0 1.1771 0 -2.0 1e-06 
0.0 1.1772 0 -2.0 1e-06 
0.0 1.1773 0 -2.0 1e-06 
0.0 1.1774 0 -2.0 1e-06 
0.0 1.1775 0 -2.0 1e-06 
0.0 1.1776 0 -2.0 1e-06 
0.0 1.1777 0 -2.0 1e-06 
0.0 1.1778 0 -2.0 1e-06 
0.0 1.1779 0 -2.0 1e-06 
0.0 1.178 0 -2.0 1e-06 
0.0 1.1781 0 -2.0 1e-06 
0.0 1.1782 0 -2.0 1e-06 
0.0 1.1783 0 -2.0 1e-06 
0.0 1.1784 0 -2.0 1e-06 
0.0 1.1785 0 -2.0 1e-06 
0.0 1.1786 0 -2.0 1e-06 
0.0 1.1787 0 -2.0 1e-06 
0.0 1.1788 0 -2.0 1e-06 
0.0 1.1789 0 -2.0 1e-06 
0.0 1.179 0 -2.0 1e-06 
0.0 1.1791 0 -2.0 1e-06 
0.0 1.1792 0 -2.0 1e-06 
0.0 1.1793 0 -2.0 1e-06 
0.0 1.1794 0 -2.0 1e-06 
0.0 1.1795 0 -2.0 1e-06 
0.0 1.1796 0 -2.0 1e-06 
0.0 1.1797 0 -2.0 1e-06 
0.0 1.1798 0 -2.0 1e-06 
0.0 1.1799 0 -2.0 1e-06 
0.0 1.18 0 -2.0 1e-06 
0.0 1.1801 0 -2.0 1e-06 
0.0 1.1802 0 -2.0 1e-06 
0.0 1.1803 0 -2.0 1e-06 
0.0 1.1804 0 -2.0 1e-06 
0.0 1.1805 0 -2.0 1e-06 
0.0 1.1806 0 -2.0 1e-06 
0.0 1.1807 0 -2.0 1e-06 
0.0 1.1808 0 -2.0 1e-06 
0.0 1.1809 0 -2.0 1e-06 
0.0 1.181 0 -2.0 1e-06 
0.0 1.1811 0 -2.0 1e-06 
0.0 1.1812 0 -2.0 1e-06 
0.0 1.1813 0 -2.0 1e-06 
0.0 1.1814 0 -2.0 1e-06 
0.0 1.1815 0 -2.0 1e-06 
0.0 1.1816 0 -2.0 1e-06 
0.0 1.1817 0 -2.0 1e-06 
0.0 1.1818 0 -2.0 1e-06 
0.0 1.1819 0 -2.0 1e-06 
0.0 1.182 0 -2.0 1e-06 
0.0 1.1821 0 -2.0 1e-06 
0.0 1.1822 0 -2.0 1e-06 
0.0 1.1823 0 -2.0 1e-06 
0.0 1.1824 0 -2.0 1e-06 
0.0 1.1825 0 -2.0 1e-06 
0.0 1.1826 0 -2.0 1e-06 
0.0 1.1827 0 -2.0 1e-06 
0.0 1.1828 0 -2.0 1e-06 
0.0 1.1829 0 -2.0 1e-06 
0.0 1.183 0 -2.0 1e-06 
0.0 1.1831 0 -2.0 1e-06 
0.0 1.1832 0 -2.0 1e-06 
0.0 1.1833 0 -2.0 1e-06 
0.0 1.1834 0 -2.0 1e-06 
0.0 1.1835 0 -2.0 1e-06 
0.0 1.1836 0 -2.0 1e-06 
0.0 1.1837 0 -2.0 1e-06 
0.0 1.1838 0 -2.0 1e-06 
0.0 1.1839 0 -2.0 1e-06 
0.0 1.184 0 -2.0 1e-06 
0.0 1.1841 0 -2.0 1e-06 
0.0 1.1842 0 -2.0 1e-06 
0.0 1.1843 0 -2.0 1e-06 
0.0 1.1844 0 -2.0 1e-06 
0.0 1.1845 0 -2.0 1e-06 
0.0 1.1846 0 -2.0 1e-06 
0.0 1.1847 0 -2.0 1e-06 
0.0 1.1848 0 -2.0 1e-06 
0.0 1.1849 0 -2.0 1e-06 
0.0 1.185 0 -2.0 1e-06 
0.0 1.1851 0 -2.0 1e-06 
0.0 1.1852 0 -2.0 1e-06 
0.0 1.1853 0 -2.0 1e-06 
0.0 1.1854 0 -2.0 1e-06 
0.0 1.1855 0 -2.0 1e-06 
0.0 1.1856 0 -2.0 1e-06 
0.0 1.1857 0 -2.0 1e-06 
0.0 1.1858 0 -2.0 1e-06 
0.0 1.1859 0 -2.0 1e-06 
0.0 1.186 0 -2.0 1e-06 
0.0 1.1861 0 -2.0 1e-06 
0.0 1.1862 0 -2.0 1e-06 
0.0 1.1863 0 -2.0 1e-06 
0.0 1.1864 0 -2.0 1e-06 
0.0 1.1865 0 -2.0 1e-06 
0.0 1.1866 0 -2.0 1e-06 
0.0 1.1867 0 -2.0 1e-06 
0.0 1.1868 0 -2.0 1e-06 
0.0 1.1869 0 -2.0 1e-06 
0.0 1.187 0 -2.0 1e-06 
0.0 1.1871 0 -2.0 1e-06 
0.0 1.1872 0 -2.0 1e-06 
0.0 1.1873 0 -2.0 1e-06 
0.0 1.1874 0 -2.0 1e-06 
0.0 1.1875 0 -2.0 1e-06 
0.0 1.1876 0 -2.0 1e-06 
0.0 1.1877 0 -2.0 1e-06 
0.0 1.1878 0 -2.0 1e-06 
0.0 1.1879 0 -2.0 1e-06 
0.0 1.188 0 -2.0 1e-06 
0.0 1.1881 0 -2.0 1e-06 
0.0 1.1882 0 -2.0 1e-06 
0.0 1.1883 0 -2.0 1e-06 
0.0 1.1884 0 -2.0 1e-06 
0.0 1.1885 0 -2.0 1e-06 
0.0 1.1886 0 -2.0 1e-06 
0.0 1.1887 0 -2.0 1e-06 
0.0 1.1888 0 -2.0 1e-06 
0.0 1.1889 0 -2.0 1e-06 
0.0 1.189 0 -2.0 1e-06 
0.0 1.1891 0 -2.0 1e-06 
0.0 1.1892 0 -2.0 1e-06 
0.0 1.1893 0 -2.0 1e-06 
0.0 1.1894 0 -2.0 1e-06 
0.0 1.1895 0 -2.0 1e-06 
0.0 1.1896 0 -2.0 1e-06 
0.0 1.1897 0 -2.0 1e-06 
0.0 1.1898 0 -2.0 1e-06 
0.0 1.1899 0 -2.0 1e-06 
0.0 1.19 0 -2.0 1e-06 
0.0 1.1901 0 -2.0 1e-06 
0.0 1.1902 0 -2.0 1e-06 
0.0 1.1903 0 -2.0 1e-06 
0.0 1.1904 0 -2.0 1e-06 
0.0 1.1905 0 -2.0 1e-06 
0.0 1.1906 0 -2.0 1e-06 
0.0 1.1907 0 -2.0 1e-06 
0.0 1.1908 0 -2.0 1e-06 
0.0 1.1909 0 -2.0 1e-06 
0.0 1.191 0 -2.0 1e-06 
0.0 1.1911 0 -2.0 1e-06 
0.0 1.1912 0 -2.0 1e-06 
0.0 1.1913 0 -2.0 1e-06 
0.0 1.1914 0 -2.0 1e-06 
0.0 1.1915 0 -2.0 1e-06 
0.0 1.1916 0 -2.0 1e-06 
0.0 1.1917 0 -2.0 1e-06 
0.0 1.1918 0 -2.0 1e-06 
0.0 1.1919 0 -2.0 1e-06 
0.0 1.192 0 -2.0 1e-06 
0.0 1.1921 0 -2.0 1e-06 
0.0 1.1922 0 -2.0 1e-06 
0.0 1.1923 0 -2.0 1e-06 
0.0 1.1924 0 -2.0 1e-06 
0.0 1.1925 0 -2.0 1e-06 
0.0 1.1926 0 -2.0 1e-06 
0.0 1.1927 0 -2.0 1e-06 
0.0 1.1928 0 -2.0 1e-06 
0.0 1.1929 0 -2.0 1e-06 
0.0 1.193 0 -2.0 1e-06 
0.0 1.1931 0 -2.0 1e-06 
0.0 1.1932 0 -2.0 1e-06 
0.0 1.1933 0 -2.0 1e-06 
0.0 1.1934 0 -2.0 1e-06 
0.0 1.1935 0 -2.0 1e-06 
0.0 1.1936 0 -2.0 1e-06 
0.0 1.1937 0 -2.0 1e-06 
0.0 1.1938 0 -2.0 1e-06 
0.0 1.1939 0 -2.0 1e-06 
0.0 1.194 0 -2.0 1e-06 
0.0 1.1941 0 -2.0 1e-06 
0.0 1.1942 0 -2.0 1e-06 
0.0 1.1943 0 -2.0 1e-06 
0.0 1.1944 0 -2.0 1e-06 
0.0 1.1945 0 -2.0 1e-06 
0.0 1.1946 0 -2.0 1e-06 
0.0 1.1947 0 -2.0 1e-06 
0.0 1.1948 0 -2.0 1e-06 
0.0 1.1949 0 -2.0 1e-06 
0.0 1.195 0 -2.0 1e-06 
0.0 1.1951 0 -2.0 1e-06 
0.0 1.1952 0 -2.0 1e-06 
0.0 1.1953 0 -2.0 1e-06 
0.0 1.1954 0 -2.0 1e-06 
0.0 1.1955 0 -2.0 1e-06 
0.0 1.1956 0 -2.0 1e-06 
0.0 1.1957 0 -2.0 1e-06 
0.0 1.1958 0 -2.0 1e-06 
0.0 1.1959 0 -2.0 1e-06 
0.0 1.196 0 -2.0 1e-06 
0.0 1.1961 0 -2.0 1e-06 
0.0 1.1962 0 -2.0 1e-06 
0.0 1.1963 0 -2.0 1e-06 
0.0 1.1964 0 -2.0 1e-06 
0.0 1.1965 0 -2.0 1e-06 
0.0 1.1966 0 -2.0 1e-06 
0.0 1.1967 0 -2.0 1e-06 
0.0 1.1968 0 -2.0 1e-06 
0.0 1.1969 0 -2.0 1e-06 
0.0 1.197 0 -2.0 1e-06 
0.0 1.1971 0 -2.0 1e-06 
0.0 1.1972 0 -2.0 1e-06 
0.0 1.1973 0 -2.0 1e-06 
0.0 1.1974 0 -2.0 1e-06 
0.0 1.1975 0 -2.0 1e-06 
0.0 1.1976 0 -2.0 1e-06 
0.0 1.1977 0 -2.0 1e-06 
0.0 1.1978 0 -2.0 1e-06 
0.0 1.1979 0 -2.0 1e-06 
0.0 1.198 0 -2.0 1e-06 
0.0 1.1981 0 -2.0 1e-06 
0.0 1.1982 0 -2.0 1e-06 
0.0 1.1983 0 -2.0 1e-06 
0.0 1.1984 0 -2.0 1e-06 
0.0 1.1985 0 -2.0 1e-06 
0.0 1.1986 0 -2.0 1e-06 
0.0 1.1987 0 -2.0 1e-06 
0.0 1.1988 0 -2.0 1e-06 
0.0 1.1989 0 -2.0 1e-06 
0.0 1.199 0 -2.0 1e-06 
0.0 1.1991 0 -2.0 1e-06 
0.0 1.1992 0 -2.0 1e-06 
0.0 1.1993 0 -2.0 1e-06 
0.0 1.1994 0 -2.0 1e-06 
0.0 1.1995 0 -2.0 1e-06 
0.0 1.1996 0 -2.0 1e-06 
0.0 1.1997 0 -2.0 1e-06 
0.0 1.1998 0 -2.0 1e-06 
0.0 1.1999 0 -2.0 1e-06 
0.0 1.2 0 -2.0 1e-06 
0.0 1.2001 0 -2.0 1e-06 
0.0 1.2002 0 -2.0 1e-06 
0.0 1.2003 0 -2.0 1e-06 
0.0 1.2004 0 -2.0 1e-06 
0.0 1.2005 0 -2.0 1e-06 
0.0 1.2006 0 -2.0 1e-06 
0.0 1.2007 0 -2.0 1e-06 
0.0 1.2008 0 -2.0 1e-06 
0.0 1.2009 0 -2.0 1e-06 
0.0 1.201 0 -2.0 1e-06 
0.0 1.2011 0 -2.0 1e-06 
0.0 1.2012 0 -2.0 1e-06 
0.0 1.2013 0 -2.0 1e-06 
0.0 1.2014 0 -2.0 1e-06 
0.0 1.2015 0 -2.0 1e-06 
0.0 1.2016 0 -2.0 1e-06 
0.0 1.2017 0 -2.0 1e-06 
0.0 1.2018 0 -2.0 1e-06 
0.0 1.2019 0 -2.0 1e-06 
0.0 1.202 0 -2.0 1e-06 
0.0 1.2021 0 -2.0 1e-06 
0.0 1.2022 0 -2.0 1e-06 
0.0 1.2023 0 -2.0 1e-06 
0.0 1.2024 0 -2.0 1e-06 
0.0 1.2025 0 -2.0 1e-06 
0.0 1.2026 0 -2.0 1e-06 
0.0 1.2027 0 -2.0 1e-06 
0.0 1.2028 0 -2.0 1e-06 
0.0 1.2029 0 -2.0 1e-06 
0.0 1.203 0 -2.0 1e-06 
0.0 1.2031 0 -2.0 1e-06 
0.0 1.2032 0 -2.0 1e-06 
0.0 1.2033 0 -2.0 1e-06 
0.0 1.2034 0 -2.0 1e-06 
0.0 1.2035 0 -2.0 1e-06 
0.0 1.2036 0 -2.0 1e-06 
0.0 1.2037 0 -2.0 1e-06 
0.0 1.2038 0 -2.0 1e-06 
0.0 1.2039 0 -2.0 1e-06 
0.0 1.204 0 -2.0 1e-06 
0.0 1.2041 0 -2.0 1e-06 
0.0 1.2042 0 -2.0 1e-06 
0.0 1.2043 0 -2.0 1e-06 
0.0 1.2044 0 -2.0 1e-06 
0.0 1.2045 0 -2.0 1e-06 
0.0 1.2046 0 -2.0 1e-06 
0.0 1.2047 0 -2.0 1e-06 
0.0 1.2048 0 -2.0 1e-06 
0.0 1.2049 0 -2.0 1e-06 
0.0 1.205 0 -2.0 1e-06 
0.0 1.2051 0 -2.0 1e-06 
0.0 1.2052 0 -2.0 1e-06 
0.0 1.2053 0 -2.0 1e-06 
0.0 1.2054 0 -2.0 1e-06 
0.0 1.2055 0 -2.0 1e-06 
0.0 1.2056 0 -2.0 1e-06 
0.0 1.2057 0 -2.0 1e-06 
0.0 1.2058 0 -2.0 1e-06 
0.0 1.2059 0 -2.0 1e-06 
0.0 1.206 0 -2.0 1e-06 
0.0 1.2061 0 -2.0 1e-06 
0.0 1.2062 0 -2.0 1e-06 
0.0 1.2063 0 -2.0 1e-06 
0.0 1.2064 0 -2.0 1e-06 
0.0 1.2065 0 -2.0 1e-06 
0.0 1.2066 0 -2.0 1e-06 
0.0 1.2067 0 -2.0 1e-06 
0.0 1.2068 0 -2.0 1e-06 
0.0 1.2069 0 -2.0 1e-06 
0.0 1.207 0 -2.0 1e-06 
0.0 1.2071 0 -2.0 1e-06 
0.0 1.2072 0 -2.0 1e-06 
0.0 1.2073 0 -2.0 1e-06 
0.0 1.2074 0 -2.0 1e-06 
0.0 1.2075 0 -2.0 1e-06 
0.0 1.2076 0 -2.0 1e-06 
0.0 1.2077 0 -2.0 1e-06 
0.0 1.2078 0 -2.0 1e-06 
0.0 1.2079 0 -2.0 1e-06 
0.0 1.208 0 -2.0 1e-06 
0.0 1.2081 0 -2.0 1e-06 
0.0 1.2082 0 -2.0 1e-06 
0.0 1.2083 0 -2.0 1e-06 
0.0 1.2084 0 -2.0 1e-06 
0.0 1.2085 0 -2.0 1e-06 
0.0 1.2086 0 -2.0 1e-06 
0.0 1.2087 0 -2.0 1e-06 
0.0 1.2088 0 -2.0 1e-06 
0.0 1.2089 0 -2.0 1e-06 
0.0 1.209 0 -2.0 1e-06 
0.0 1.2091 0 -2.0 1e-06 
0.0 1.2092 0 -2.0 1e-06 
0.0 1.2093 0 -2.0 1e-06 
0.0 1.2094 0 -2.0 1e-06 
0.0 1.2095 0 -2.0 1e-06 
0.0 1.2096 0 -2.0 1e-06 
0.0 1.2097 0 -2.0 1e-06 
0.0 1.2098 0 -2.0 1e-06 
0.0 1.2099 0 -2.0 1e-06 
0.0 1.21 0 -2.0 1e-06 
0.0 1.2101 0 -2.0 1e-06 
0.0 1.2102 0 -2.0 1e-06 
0.0 1.2103 0 -2.0 1e-06 
0.0 1.2104 0 -2.0 1e-06 
0.0 1.2105 0 -2.0 1e-06 
0.0 1.2106 0 -2.0 1e-06 
0.0 1.2107 0 -2.0 1e-06 
0.0 1.2108 0 -2.0 1e-06 
0.0 1.2109 0 -2.0 1e-06 
0.0 1.211 0 -2.0 1e-06 
0.0 1.2111 0 -2.0 1e-06 
0.0 1.2112 0 -2.0 1e-06 
0.0 1.2113 0 -2.0 1e-06 
0.0 1.2114 0 -2.0 1e-06 
0.0 1.2115 0 -2.0 1e-06 
0.0 1.2116 0 -2.0 1e-06 
0.0 1.2117 0 -2.0 1e-06 
0.0 1.2118 0 -2.0 1e-06 
0.0 1.2119 0 -2.0 1e-06 
0.0 1.212 0 -2.0 1e-06 
0.0 1.2121 0 -2.0 1e-06 
0.0 1.2122 0 -2.0 1e-06 
0.0 1.2123 0 -2.0 1e-06 
0.0 1.2124 0 -2.0 1e-06 
0.0 1.2125 0 -2.0 1e-06 
0.0 1.2126 0 -2.0 1e-06 
0.0 1.2127 0 -2.0 1e-06 
0.0 1.2128 0 -2.0 1e-06 
0.0 1.2129 0 -2.0 1e-06 
0.0 1.213 0 -2.0 1e-06 
0.0 1.2131 0 -2.0 1e-06 
0.0 1.2132 0 -2.0 1e-06 
0.0 1.2133 0 -2.0 1e-06 
0.0 1.2134 0 -2.0 1e-06 
0.0 1.2135 0 -2.0 1e-06 
0.0 1.2136 0 -2.0 1e-06 
0.0 1.2137 0 -2.0 1e-06 
0.0 1.2138 0 -2.0 1e-06 
0.0 1.2139 0 -2.0 1e-06 
0.0 1.214 0 -2.0 1e-06 
0.0 1.2141 0 -2.0 1e-06 
0.0 1.2142 0 -2.0 1e-06 
0.0 1.2143 0 -2.0 1e-06 
0.0 1.2144 0 -2.0 1e-06 
0.0 1.2145 0 -2.0 1e-06 
0.0 1.2146 0 -2.0 1e-06 
0.0 1.2147 0 -2.0 1e-06 
0.0 1.2148 0 -2.0 1e-06 
0.0 1.2149 0 -2.0 1e-06 
0.0 1.215 0 -2.0 1e-06 
0.0 1.2151 0 -2.0 1e-06 
0.0 1.2152 0 -2.0 1e-06 
0.0 1.2153 0 -2.0 1e-06 
0.0 1.2154 0 -2.0 1e-06 
0.0 1.2155 0 -2.0 1e-06 
0.0 1.2156 0 -2.0 1e-06 
0.0 1.2157 0 -2.0 1e-06 
0.0 1.2158 0 -2.0 1e-06 
0.0 1.2159 0 -2.0 1e-06 
0.0 1.216 0 -2.0 1e-06 
0.0 1.2161 0 -2.0 1e-06 
0.0 1.2162 0 -2.0 1e-06 
0.0 1.2163 0 -2.0 1e-06 
0.0 1.2164 0 -2.0 1e-06 
0.0 1.2165 0 -2.0 1e-06 
0.0 1.2166 0 -2.0 1e-06 
0.0 1.2167 0 -2.0 1e-06 
0.0 1.2168 0 -2.0 1e-06 
0.0 1.2169 0 -2.0 1e-06 
0.0 1.217 0 -2.0 1e-06 
0.0 1.2171 0 -2.0 1e-06 
0.0 1.2172 0 -2.0 1e-06 
0.0 1.2173 0 -2.0 1e-06 
0.0 1.2174 0 -2.0 1e-06 
0.0 1.2175 0 -2.0 1e-06 
0.0 1.2176 0 -2.0 1e-06 
0.0 1.2177 0 -2.0 1e-06 
0.0 1.2178 0 -2.0 1e-06 
0.0 1.2179 0 -2.0 1e-06 
0.0 1.218 0 -2.0 1e-06 
0.0 1.2181 0 -2.0 1e-06 
0.0 1.2182 0 -2.0 1e-06 
0.0 1.2183 0 -2.0 1e-06 
0.0 1.2184 0 -2.0 1e-06 
0.0 1.2185 0 -2.0 1e-06 
0.0 1.2186 0 -2.0 1e-06 
0.0 1.2187 0 -2.0 1e-06 
0.0 1.2188 0 -2.0 1e-06 
0.0 1.2189 0 -2.0 1e-06 
0.0 1.219 0 -2.0 1e-06 
0.0 1.2191 0 -2.0 1e-06 
0.0 1.2192 0 -2.0 1e-06 
0.0 1.2193 0 -2.0 1e-06 
0.0 1.2194 0 -2.0 1e-06 
0.0 1.2195 0 -2.0 1e-06 
0.0 1.2196 0 -2.0 1e-06 
0.0 1.2197 0 -2.0 1e-06 
0.0 1.2198 0 -2.0 1e-06 
0.0 1.2199 0 -2.0 1e-06 
0.0 1.22 0 -2.0 1e-06 
0.0 1.2201 0 -2.0 1e-06 
0.0 1.2202 0 -2.0 1e-06 
0.0 1.2203 0 -2.0 1e-06 
0.0 1.2204 0 -2.0 1e-06 
0.0 1.2205 0 -2.0 1e-06 
0.0 1.2206 0 -2.0 1e-06 
0.0 1.2207 0 -2.0 1e-06 
0.0 1.2208 0 -2.0 1e-06 
0.0 1.2209 0 -2.0 1e-06 
0.0 1.221 0 -2.0 1e-06 
0.0 1.2211 0 -2.0 1e-06 
0.0 1.2212 0 -2.0 1e-06 
0.0 1.2213 0 -2.0 1e-06 
0.0 1.2214 0 -2.0 1e-06 
0.0 1.2215 0 -2.0 1e-06 
0.0 1.2216 0 -2.0 1e-06 
0.0 1.2217 0 -2.0 1e-06 
0.0 1.2218 0 -2.0 1e-06 
0.0 1.2219 0 -2.0 1e-06 
0.0 1.222 0 -2.0 1e-06 
0.0 1.2221 0 -2.0 1e-06 
0.0 1.2222 0 -2.0 1e-06 
0.0 1.2223 0 -2.0 1e-06 
0.0 1.2224 0 -2.0 1e-06 
0.0 1.2225 0 -2.0 1e-06 
0.0 1.2226 0 -2.0 1e-06 
0.0 1.2227 0 -2.0 1e-06 
0.0 1.2228 0 -2.0 1e-06 
0.0 1.2229 0 -2.0 1e-06 
0.0 1.223 0 -2.0 1e-06 
0.0 1.2231 0 -2.0 1e-06 
0.0 1.2232 0 -2.0 1e-06 
0.0 1.2233 0 -2.0 1e-06 
0.0 1.2234 0 -2.0 1e-06 
0.0 1.2235 0 -2.0 1e-06 
0.0 1.2236 0 -2.0 1e-06 
0.0 1.2237 0 -2.0 1e-06 
0.0 1.2238 0 -2.0 1e-06 
0.0 1.2239 0 -2.0 1e-06 
0.0 1.224 0 -2.0 1e-06 
0.0 1.2241 0 -2.0 1e-06 
0.0 1.2242 0 -2.0 1e-06 
0.0 1.2243 0 -2.0 1e-06 
0.0 1.2244 0 -2.0 1e-06 
0.0 1.2245 0 -2.0 1e-06 
0.0 1.2246 0 -2.0 1e-06 
0.0 1.2247 0 -2.0 1e-06 
0.0 1.2248 0 -2.0 1e-06 
0.0 1.2249 0 -2.0 1e-06 
0.0 1.225 0 -2.0 1e-06 
0.0 1.2251 0 -2.0 1e-06 
0.0 1.2252 0 -2.0 1e-06 
0.0 1.2253 0 -2.0 1e-06 
0.0 1.2254 0 -2.0 1e-06 
0.0 1.2255 0 -2.0 1e-06 
0.0 1.2256 0 -2.0 1e-06 
0.0 1.2257 0 -2.0 1e-06 
0.0 1.2258 0 -2.0 1e-06 
0.0 1.2259 0 -2.0 1e-06 
0.0 1.226 0 -2.0 1e-06 
0.0 1.2261 0 -2.0 1e-06 
0.0 1.2262 0 -2.0 1e-06 
0.0 1.2263 0 -2.0 1e-06 
0.0 1.2264 0 -2.0 1e-06 
0.0 1.2265 0 -2.0 1e-06 
0.0 1.2266 0 -2.0 1e-06 
0.0 1.2267 0 -2.0 1e-06 
0.0 1.2268 0 -2.0 1e-06 
0.0 1.2269 0 -2.0 1e-06 
0.0 1.227 0 -2.0 1e-06 
0.0 1.2271 0 -2.0 1e-06 
0.0 1.2272 0 -2.0 1e-06 
0.0 1.2273 0 -2.0 1e-06 
0.0 1.2274 0 -2.0 1e-06 
0.0 1.2275 0 -2.0 1e-06 
0.0 1.2276 0 -2.0 1e-06 
0.0 1.2277 0 -2.0 1e-06 
0.0 1.2278 0 -2.0 1e-06 
0.0 1.2279 0 -2.0 1e-06 
0.0 1.228 0 -2.0 1e-06 
0.0 1.2281 0 -2.0 1e-06 
0.0 1.2282 0 -2.0 1e-06 
0.0 1.2283 0 -2.0 1e-06 
0.0 1.2284 0 -2.0 1e-06 
0.0 1.2285 0 -2.0 1e-06 
0.0 1.2286 0 -2.0 1e-06 
0.0 1.2287 0 -2.0 1e-06 
0.0 1.2288 0 -2.0 1e-06 
0.0 1.2289 0 -2.0 1e-06 
0.0 1.229 0 -2.0 1e-06 
0.0 1.2291 0 -2.0 1e-06 
0.0 1.2292 0 -2.0 1e-06 
0.0 1.2293 0 -2.0 1e-06 
0.0 1.2294 0 -2.0 1e-06 
0.0 1.2295 0 -2.0 1e-06 
0.0 1.2296 0 -2.0 1e-06 
0.0 1.2297 0 -2.0 1e-06 
0.0 1.2298 0 -2.0 1e-06 
0.0 1.2299 0 -2.0 1e-06 
0.0 1.23 0 -2.0 1e-06 
0.0 1.2301 0 -2.0 1e-06 
0.0 1.2302 0 -2.0 1e-06 
0.0 1.2303 0 -2.0 1e-06 
0.0 1.2304 0 -2.0 1e-06 
0.0 1.2305 0 -2.0 1e-06 
0.0 1.2306 0 -2.0 1e-06 
0.0 1.2307 0 -2.0 1e-06 
0.0 1.2308 0 -2.0 1e-06 
0.0 1.2309 0 -2.0 1e-06 
0.0 1.231 0 -2.0 1e-06 
0.0 1.2311 0 -2.0 1e-06 
0.0 1.2312 0 -2.0 1e-06 
0.0 1.2313 0 -2.0 1e-06 
0.0 1.2314 0 -2.0 1e-06 
0.0 1.2315 0 -2.0 1e-06 
0.0 1.2316 0 -2.0 1e-06 
0.0 1.2317 0 -2.0 1e-06 
0.0 1.2318 0 -2.0 1e-06 
0.0 1.2319 0 -2.0 1e-06 
0.0 1.232 0 -2.0 1e-06 
0.0 1.2321 0 -2.0 1e-06 
0.0 1.2322 0 -2.0 1e-06 
0.0 1.2323 0 -2.0 1e-06 
0.0 1.2324 0 -2.0 1e-06 
0.0 1.2325 0 -2.0 1e-06 
0.0 1.2326 0 -2.0 1e-06 
0.0 1.2327 0 -2.0 1e-06 
0.0 1.2328 0 -2.0 1e-06 
0.0 1.2329 0 -2.0 1e-06 
0.0 1.233 0 -2.0 1e-06 
0.0 1.2331 0 -2.0 1e-06 
0.0 1.2332 0 -2.0 1e-06 
0.0 1.2333 0 -2.0 1e-06 
0.0 1.2334 0 -2.0 1e-06 
0.0 1.2335 0 -2.0 1e-06 
0.0 1.2336 0 -2.0 1e-06 
0.0 1.2337 0 -2.0 1e-06 
0.0 1.2338 0 -2.0 1e-06 
0.0 1.2339 0 -2.0 1e-06 
0.0 1.234 0 -2.0 1e-06 
0.0 1.2341 0 -2.0 1e-06 
0.0 1.2342 0 -2.0 1e-06 
0.0 1.2343 0 -2.0 1e-06 
0.0 1.2344 0 -2.0 1e-06 
0.0 1.2345 0 -2.0 1e-06 
0.0 1.2346 0 -2.0 1e-06 
0.0 1.2347 0 -2.0 1e-06 
0.0 1.2348 0 -2.0 1e-06 
0.0 1.2349 0 -2.0 1e-06 
0.0 1.235 0 -2.0 1e-06 
0.0 1.2351 0 -2.0 1e-06 
0.0 1.2352 0 -2.0 1e-06 
0.0 1.2353 0 -2.0 1e-06 
0.0 1.2354 0 -2.0 1e-06 
0.0 1.2355 0 -2.0 1e-06 
0.0 1.2356 0 -2.0 1e-06 
0.0 1.2357 0 -2.0 1e-06 
0.0 1.2358 0 -2.0 1e-06 
0.0 1.2359 0 -2.0 1e-06 
0.0 1.236 0 -2.0 1e-06 
0.0 1.2361 0 -2.0 1e-06 
0.0 1.2362 0 -2.0 1e-06 
0.0 1.2363 0 -2.0 1e-06 
0.0 1.2364 0 -2.0 1e-06 
0.0 1.2365 0 -2.0 1e-06 
0.0 1.2366 0 -2.0 1e-06 
0.0 1.2367 0 -2.0 1e-06 
0.0 1.2368 0 -2.0 1e-06 
0.0 1.2369 0 -2.0 1e-06 
0.0 1.237 0 -2.0 1e-06 
0.0 1.2371 0 -2.0 1e-06 
0.0 1.2372 0 -2.0 1e-06 
0.0 1.2373 0 -2.0 1e-06 
0.0 1.2374 0 -2.0 1e-06 
0.0 1.2375 0 -2.0 1e-06 
0.0 1.2376 0 -2.0 1e-06 
0.0 1.2377 0 -2.0 1e-06 
0.0 1.2378 0 -2.0 1e-06 
0.0 1.2379 0 -2.0 1e-06 
0.0 1.238 0 -2.0 1e-06 
0.0 1.2381 0 -2.0 1e-06 
0.0 1.2382 0 -2.0 1e-06 
0.0 1.2383 0 -2.0 1e-06 
0.0 1.2384 0 -2.0 1e-06 
0.0 1.2385 0 -2.0 1e-06 
0.0 1.2386 0 -2.0 1e-06 
0.0 1.2387 0 -2.0 1e-06 
0.0 1.2388 0 -2.0 1e-06 
0.0 1.2389 0 -2.0 1e-06 
0.0 1.239 0 -2.0 1e-06 
0.0 1.2391 0 -2.0 1e-06 
0.0 1.2392 0 -2.0 1e-06 
0.0 1.2393 0 -2.0 1e-06 
0.0 1.2394 0 -2.0 1e-06 
0.0 1.2395 0 -2.0 1e-06 
0.0 1.2396 0 -2.0 1e-06 
0.0 1.2397 0 -2.0 1e-06 
0.0 1.2398 0 -2.0 1e-06 
0.0 1.2399 0 -2.0 1e-06 
0.0 1.24 0 -2.0 1e-06 
0.0 1.2401 0 -2.0 1e-06 
0.0 1.2402 0 -2.0 1e-06 
0.0 1.2403 0 -2.0 1e-06 
0.0 1.2404 0 -2.0 1e-06 
0.0 1.2405 0 -2.0 1e-06 
0.0 1.2406 0 -2.0 1e-06 
0.0 1.2407 0 -2.0 1e-06 
0.0 1.2408 0 -2.0 1e-06 
0.0 1.2409 0 -2.0 1e-06 
0.0 1.241 0 -2.0 1e-06 
0.0 1.2411 0 -2.0 1e-06 
0.0 1.2412 0 -2.0 1e-06 
0.0 1.2413 0 -2.0 1e-06 
0.0 1.2414 0 -2.0 1e-06 
0.0 1.2415 0 -2.0 1e-06 
0.0 1.2416 0 -2.0 1e-06 
0.0 1.2417 0 -2.0 1e-06 
0.0 1.2418 0 -2.0 1e-06 
0.0 1.2419 0 -2.0 1e-06 
0.0 1.242 0 -2.0 1e-06 
0.0 1.2421 0 -2.0 1e-06 
0.0 1.2422 0 -2.0 1e-06 
0.0 1.2423 0 -2.0 1e-06 
0.0 1.2424 0 -2.0 1e-06 
0.0 1.2425 0 -2.0 1e-06 
0.0 1.2426 0 -2.0 1e-06 
0.0 1.2427 0 -2.0 1e-06 
0.0 1.2428 0 -2.0 1e-06 
0.0 1.2429 0 -2.0 1e-06 
0.0 1.243 0 -2.0 1e-06 
0.0 1.2431 0 -2.0 1e-06 
0.0 1.2432 0 -2.0 1e-06 
0.0 1.2433 0 -2.0 1e-06 
0.0 1.2434 0 -2.0 1e-06 
0.0 1.2435 0 -2.0 1e-06 
0.0 1.2436 0 -2.0 1e-06 
0.0 1.2437 0 -2.0 1e-06 
0.0 1.2438 0 -2.0 1e-06 
0.0 1.2439 0 -2.0 1e-06 
0.0 1.244 0 -2.0 1e-06 
0.0 1.2441 0 -2.0 1e-06 
0.0 1.2442 0 -2.0 1e-06 
0.0 1.2443 0 -2.0 1e-06 
0.0 1.2444 0 -2.0 1e-06 
0.0 1.2445 0 -2.0 1e-06 
0.0 1.2446 0 -2.0 1e-06 
0.0 1.2447 0 -2.0 1e-06 
0.0 1.2448 0 -2.0 1e-06 
0.0 1.2449 0 -2.0 1e-06 
0.0 1.245 0 -2.0 1e-06 
0.0 1.2451 0 -2.0 1e-06 
0.0 1.2452 0 -2.0 1e-06 
0.0 1.2453 0 -2.0 1e-06 
0.0 1.2454 0 -2.0 1e-06 
0.0 1.2455 0 -2.0 1e-06 
0.0 1.2456 0 -2.0 1e-06 
0.0 1.2457 0 -2.0 1e-06 
0.0 1.2458 0 -2.0 1e-06 
0.0 1.2459 0 -2.0 1e-06 
0.0 1.246 0 -2.0 1e-06 
0.0 1.2461 0 -2.0 1e-06 
0.0 1.2462 0 -2.0 1e-06 
0.0 1.2463 0 -2.0 1e-06 
0.0 1.2464 0 -2.0 1e-06 
0.0 1.2465 0 -2.0 1e-06 
0.0 1.2466 0 -2.0 1e-06 
0.0 1.2467 0 -2.0 1e-06 
0.0 1.2468 0 -2.0 1e-06 
0.0 1.2469 0 -2.0 1e-06 
0.0 1.247 0 -2.0 1e-06 
0.0 1.2471 0 -2.0 1e-06 
0.0 1.2472 0 -2.0 1e-06 
0.0 1.2473 0 -2.0 1e-06 
0.0 1.2474 0 -2.0 1e-06 
0.0 1.2475 0 -2.0 1e-06 
0.0 1.2476 0 -2.0 1e-06 
0.0 1.2477 0 -2.0 1e-06 
0.0 1.2478 0 -2.0 1e-06 
0.0 1.2479 0 -2.0 1e-06 
0.0 1.248 0 -2.0 1e-06 
0.0 1.2481 0 -2.0 1e-06 
0.0 1.2482 0 -2.0 1e-06 
0.0 1.2483 0 -2.0 1e-06 
0.0 1.2484 0 -2.0 1e-06 
0.0 1.2485 0 -2.0 1e-06 
0.0 1.2486 0 -2.0 1e-06 
0.0 1.2487 0 -2.0 1e-06 
0.0 1.2488 0 -2.0 1e-06 
0.0 1.2489 0 -2.0 1e-06 
0.0 1.249 0 -2.0 1e-06 
0.0 1.2491 0 -2.0 1e-06 
0.0 1.2492 0 -2.0 1e-06 
0.0 1.2493 0 -2.0 1e-06 
0.0 1.2494 0 -2.0 1e-06 
0.0 1.2495 0 -2.0 1e-06 
0.0 1.2496 0 -2.0 1e-06 
0.0 1.2497 0 -2.0 1e-06 
0.0 1.2498 0 -2.0 1e-06 
0.0 1.2499 0 -2.0 1e-06 
0.0 1.25 0 -2.0 1e-06 
0.0 1.2501 0 -2.0 1e-06 
0.0 1.2502 0 -2.0 1e-06 
0.0 1.2503 0 -2.0 1e-06 
0.0 1.2504 0 -2.0 1e-06 
0.0 1.2505 0 -2.0 1e-06 
0.0 1.2506 0 -2.0 1e-06 
0.0 1.2507 0 -2.0 1e-06 
0.0 1.2508 0 -2.0 1e-06 
0.0 1.2509 0 -2.0 1e-06 
0.0 1.251 0 -2.0 1e-06 
0.0 1.2511 0 -2.0 1e-06 
0.0 1.2512 0 -2.0 1e-06 
0.0 1.2513 0 -2.0 1e-06 
0.0 1.2514 0 -2.0 1e-06 
0.0 1.2515 0 -2.0 1e-06 
0.0 1.2516 0 -2.0 1e-06 
0.0 1.2517 0 -2.0 1e-06 
0.0 1.2518 0 -2.0 1e-06 
0.0 1.2519 0 -2.0 1e-06 
0.0 1.252 0 -2.0 1e-06 
0.0 1.2521 0 -2.0 1e-06 
0.0 1.2522 0 -2.0 1e-06 
0.0 1.2523 0 -2.0 1e-06 
0.0 1.2524 0 -2.0 1e-06 
0.0 1.2525 0 -2.0 1e-06 
0.0 1.2526 0 -2.0 1e-06 
0.0 1.2527 0 -2.0 1e-06 
0.0 1.2528 0 -2.0 1e-06 
0.0 1.2529 0 -2.0 1e-06 
0.0 1.253 0 -2.0 1e-06 
0.0 1.2531 0 -2.0 1e-06 
0.0 1.2532 0 -2.0 1e-06 
0.0 1.2533 0 -2.0 1e-06 
0.0 1.2534 0 -2.0 1e-06 
0.0 1.2535 0 -2.0 1e-06 
0.0 1.2536 0 -2.0 1e-06 
0.0 1.2537 0 -2.0 1e-06 
0.0 1.2538 0 -2.0 1e-06 
0.0 1.2539 0 -2.0 1e-06 
0.0 1.254 0 -2.0 1e-06 
0.0 1.2541 0 -2.0 1e-06 
0.0 1.2542 0 -2.0 1e-06 
0.0 1.2543 0 -2.0 1e-06 
0.0 1.2544 0 -2.0 1e-06 
0.0 1.2545 0 -2.0 1e-06 
0.0 1.2546 0 -2.0 1e-06 
0.0 1.2547 0 -2.0 1e-06 
0.0 1.2548 0 -2.0 1e-06 
0.0 1.2549 0 -2.0 1e-06 
0.0 1.255 0 -2.0 1e-06 
0.0 1.2551 0 -2.0 1e-06 
0.0 1.2552 0 -2.0 1e-06 
0.0 1.2553 0 -2.0 1e-06 
0.0 1.2554 0 -2.0 1e-06 
0.0 1.2555 0 -2.0 1e-06 
0.0 1.2556 0 -2.0 1e-06 
0.0 1.2557 0 -2.0 1e-06 
0.0 1.2558 0 -2.0 1e-06 
0.0 1.2559 0 -2.0 1e-06 
0.0 1.256 0 -2.0 1e-06 
0.0 1.2561 0 -2.0 1e-06 
0.0 1.2562 0 -2.0 1e-06 
0.0 1.2563 0 -2.0 1e-06 
0.0 1.2564 0 -2.0 1e-06 
0.0 1.2565 0 -2.0 1e-06 
0.0 1.2566 0 -2.0 1e-06 
0.0 1.2567 0 -2.0 1e-06 
0.0 1.2568 0 -2.0 1e-06 
0.0 1.2569 0 -2.0 1e-06 
0.0 1.257 0 -2.0 1e-06 
0.0 1.2571 0 -2.0 1e-06 
0.0 1.2572 0 -2.0 1e-06 
0.0 1.2573 0 -2.0 1e-06 
0.0 1.2574 0 -2.0 1e-06 
0.0 1.2575 0 -2.0 1e-06 
0.0 1.2576 0 -2.0 1e-06 
0.0 1.2577 0 -2.0 1e-06 
0.0 1.2578 0 -2.0 1e-06 
0.0 1.2579 0 -2.0 1e-06 
0.0 1.258 0 -2.0 1e-06 
0.0 1.2581 0 -2.0 1e-06 
0.0 1.2582 0 -2.0 1e-06 
0.0 1.2583 0 -2.0 1e-06 
0.0 1.2584 0 -2.0 1e-06 
0.0 1.2585 0 -2.0 1e-06 
0.0 1.2586 0 -2.0 1e-06 
0.0 1.2587 0 -2.0 1e-06 
0.0 1.2588 0 -2.0 1e-06 
0.0 1.2589 0 -2.0 1e-06 
0.0 1.259 0 -2.0 1e-06 
0.0 1.2591 0 -2.0 1e-06 
0.0 1.2592 0 -2.0 1e-06 
0.0 1.2593 0 -2.0 1e-06 
0.0 1.2594 0 -2.0 1e-06 
0.0 1.2595 0 -2.0 1e-06 
0.0 1.2596 0 -2.0 1e-06 
0.0 1.2597 0 -2.0 1e-06 
0.0 1.2598 0 -2.0 1e-06 
0.0 1.2599 0 -2.0 1e-06 
0.0 1.26 0 -2.0 1e-06 
0.0 1.2601 0 -2.0 1e-06 
0.0 1.2602 0 -2.0 1e-06 
0.0 1.2603 0 -2.0 1e-06 
0.0 1.2604 0 -2.0 1e-06 
0.0 1.2605 0 -2.0 1e-06 
0.0 1.2606 0 -2.0 1e-06 
0.0 1.2607 0 -2.0 1e-06 
0.0 1.2608 0 -2.0 1e-06 
0.0 1.2609 0 -2.0 1e-06 
0.0 1.261 0 -2.0 1e-06 
0.0 1.2611 0 -2.0 1e-06 
0.0 1.2612 0 -2.0 1e-06 
0.0 1.2613 0 -2.0 1e-06 
0.0 1.2614 0 -2.0 1e-06 
0.0 1.2615 0 -2.0 1e-06 
0.0 1.2616 0 -2.0 1e-06 
0.0 1.2617 0 -2.0 1e-06 
0.0 1.2618 0 -2.0 1e-06 
0.0 1.2619 0 -2.0 1e-06 
0.0 1.262 0 -2.0 1e-06 
0.0 1.2621 0 -2.0 1e-06 
0.0 1.2622 0 -2.0 1e-06 
0.0 1.2623 0 -2.0 1e-06 
0.0 1.2624 0 -2.0 1e-06 
0.0 1.2625 0 -2.0 1e-06 
0.0 1.2626 0 -2.0 1e-06 
0.0 1.2627 0 -2.0 1e-06 
0.0 1.2628 0 -2.0 1e-06 
0.0 1.2629 0 -2.0 1e-06 
0.0 1.263 0 -2.0 1e-06 
0.0 1.2631 0 -2.0 1e-06 
0.0 1.2632 0 -2.0 1e-06 
0.0 1.2633 0 -2.0 1e-06 
0.0 1.2634 0 -2.0 1e-06 
0.0 1.2635 0 -2.0 1e-06 
0.0 1.2636 0 -2.0 1e-06 
0.0 1.2637 0 -2.0 1e-06 
0.0 1.2638 0 -2.0 1e-06 
0.0 1.2639 0 -2.0 1e-06 
0.0 1.264 0 -2.0 1e-06 
0.0 1.2641 0 -2.0 1e-06 
0.0 1.2642 0 -2.0 1e-06 
0.0 1.2643 0 -2.0 1e-06 
0.0 1.2644 0 -2.0 1e-06 
0.0 1.2645 0 -2.0 1e-06 
0.0 1.2646 0 -2.0 1e-06 
0.0 1.2647 0 -2.0 1e-06 
0.0 1.2648 0 -2.0 1e-06 
0.0 1.2649 0 -2.0 1e-06 
0.0 1.265 0 -2.0 1e-06 
0.0 1.2651 0 -2.0 1e-06 
0.0 1.2652 0 -2.0 1e-06 
0.0 1.2653 0 -2.0 1e-06 
0.0 1.2654 0 -2.0 1e-06 
0.0 1.2655 0 -2.0 1e-06 
0.0 1.2656 0 -2.0 1e-06 
0.0 1.2657 0 -2.0 1e-06 
0.0 1.2658 0 -2.0 1e-06 
0.0 1.2659 0 -2.0 1e-06 
0.0 1.266 0 -2.0 1e-06 
0.0 1.2661 0 -2.0 1e-06 
0.0 1.2662 0 -2.0 1e-06 
0.0 1.2663 0 -2.0 1e-06 
0.0 1.2664 0 -2.0 1e-06 
0.0 1.2665 0 -2.0 1e-06 
0.0 1.2666 0 -2.0 1e-06 
0.0 1.2667 0 -2.0 1e-06 
0.0 1.2668 0 -2.0 1e-06 
0.0 1.2669 0 -2.0 1e-06 
0.0 1.267 0 -2.0 1e-06 
0.0 1.2671 0 -2.0 1e-06 
0.0 1.2672 0 -2.0 1e-06 
0.0 1.2673 0 -2.0 1e-06 
0.0 1.2674 0 -2.0 1e-06 
0.0 1.2675 0 -2.0 1e-06 
0.0 1.2676 0 -2.0 1e-06 
0.0 1.2677 0 -2.0 1e-06 
0.0 1.2678 0 -2.0 1e-06 
0.0 1.2679 0 -2.0 1e-06 
0.0 1.268 0 -2.0 1e-06 
0.0 1.2681 0 -2.0 1e-06 
0.0 1.2682 0 -2.0 1e-06 
0.0 1.2683 0 -2.0 1e-06 
0.0 1.2684 0 -2.0 1e-06 
0.0 1.2685 0 -2.0 1e-06 
0.0 1.2686 0 -2.0 1e-06 
0.0 1.2687 0 -2.0 1e-06 
0.0 1.2688 0 -2.0 1e-06 
0.0 1.2689 0 -2.0 1e-06 
0.0 1.269 0 -2.0 1e-06 
0.0 1.2691 0 -2.0 1e-06 
0.0 1.2692 0 -2.0 1e-06 
0.0 1.2693 0 -2.0 1e-06 
0.0 1.2694 0 -2.0 1e-06 
0.0 1.2695 0 -2.0 1e-06 
0.0 1.2696 0 -2.0 1e-06 
0.0 1.2697 0 -2.0 1e-06 
0.0 1.2698 0 -2.0 1e-06 
0.0 1.2699 0 -2.0 1e-06 
0.0 1.27 0 -2.0 1e-06 
0.0 1.2701 0 -2.0 1e-06 
0.0 1.2702 0 -2.0 1e-06 
0.0 1.2703 0 -2.0 1e-06 
0.0 1.2704 0 -2.0 1e-06 
0.0 1.2705 0 -2.0 1e-06 
0.0 1.2706 0 -2.0 1e-06 
0.0 1.2707 0 -2.0 1e-06 
0.0 1.2708 0 -2.0 1e-06 
0.0 1.2709 0 -2.0 1e-06 
0.0 1.271 0 -2.0 1e-06 
0.0 1.2711 0 -2.0 1e-06 
0.0 1.2712 0 -2.0 1e-06 
0.0 1.2713 0 -2.0 1e-06 
0.0 1.2714 0 -2.0 1e-06 
0.0 1.2715 0 -2.0 1e-06 
0.0 1.2716 0 -2.0 1e-06 
0.0 1.2717 0 -2.0 1e-06 
0.0 1.2718 0 -2.0 1e-06 
0.0 1.2719 0 -2.0 1e-06 
0.0 1.272 0 -2.0 1e-06 
0.0 1.2721 0 -2.0 1e-06 
0.0 1.2722 0 -2.0 1e-06 
0.0 1.2723 0 -2.0 1e-06 
0.0 1.2724 0 -2.0 1e-06 
0.0 1.2725 0 -2.0 1e-06 
0.0 1.2726 0 -2.0 1e-06 
0.0 1.2727 0 -2.0 1e-06 
0.0 1.2728 0 -2.0 1e-06 
0.0 1.2729 0 -2.0 1e-06 
0.0 1.273 0 -2.0 1e-06 
0.0 1.2731 0 -2.0 1e-06 
0.0 1.2732 0 -2.0 1e-06 
0.0 1.2733 0 -2.0 1e-06 
0.0 1.2734 0 -2.0 1e-06 
0.0 1.2735 0 -2.0 1e-06 
0.0 1.2736 0 -2.0 1e-06 
0.0 1.2737 0 -2.0 1e-06 
0.0 1.2738 0 -2.0 1e-06 
0.0 1.2739 0 -2.0 1e-06 
0.0 1.274 0 -2.0 1e-06 
0.0 1.2741 0 -2.0 1e-06 
0.0 1.2742 0 -2.0 1e-06 
0.0 1.2743 0 -2.0 1e-06 
0.0 1.2744 0 -2.0 1e-06 
0.0 1.2745 0 -2.0 1e-06 
0.0 1.2746 0 -2.0 1e-06 
0.0 1.2747 0 -2.0 1e-06 
0.0 1.2748 0 -2.0 1e-06 
0.0 1.2749 0 -2.0 1e-06 
0.0 1.275 0 -2.0 1e-06 
0.0 1.2751 0 -2.0 1e-06 
0.0 1.2752 0 -2.0 1e-06 
0.0 1.2753 0 -2.0 1e-06 
0.0 1.2754 0 -2.0 1e-06 
0.0 1.2755 0 -2.0 1e-06 
0.0 1.2756 0 -2.0 1e-06 
0.0 1.2757 0 -2.0 1e-06 
0.0 1.2758 0 -2.0 1e-06 
0.0 1.2759 0 -2.0 1e-06 
0.0 1.276 0 -2.0 1e-06 
0.0 1.2761 0 -2.0 1e-06 
0.0 1.2762 0 -2.0 1e-06 
0.0 1.2763 0 -2.0 1e-06 
0.0 1.2764 0 -2.0 1e-06 
0.0 1.2765 0 -2.0 1e-06 
0.0 1.2766 0 -2.0 1e-06 
0.0 1.2767 0 -2.0 1e-06 
0.0 1.2768 0 -2.0 1e-06 
0.0 1.2769 0 -2.0 1e-06 
0.0 1.277 0 -2.0 1e-06 
0.0 1.2771 0 -2.0 1e-06 
0.0 1.2772 0 -2.0 1e-06 
0.0 1.2773 0 -2.0 1e-06 
0.0 1.2774 0 -2.0 1e-06 
0.0 1.2775 0 -2.0 1e-06 
0.0 1.2776 0 -2.0 1e-06 
0.0 1.2777 0 -2.0 1e-06 
0.0 1.2778 0 -2.0 1e-06 
0.0 1.2779 0 -2.0 1e-06 
0.0 1.278 0 -2.0 1e-06 
0.0 1.2781 0 -2.0 1e-06 
0.0 1.2782 0 -2.0 1e-06 
0.0 1.2783 0 -2.0 1e-06 
0.0 1.2784 0 -2.0 1e-06 
0.0 1.2785 0 -2.0 1e-06 
0.0 1.2786 0 -2.0 1e-06 
0.0 1.2787 0 -2.0 1e-06 
0.0 1.2788 0 -2.0 1e-06 
0.0 1.2789 0 -2.0 1e-06 
0.0 1.279 0 -2.0 1e-06 
0.0 1.2791 0 -2.0 1e-06 
0.0 1.2792 0 -2.0 1e-06 
0.0 1.2793 0 -2.0 1e-06 
0.0 1.2794 0 -2.0 1e-06 
0.0 1.2795 0 -2.0 1e-06 
0.0 1.2796 0 -2.0 1e-06 
0.0 1.2797 0 -2.0 1e-06 
0.0 1.2798 0 -2.0 1e-06 
0.0 1.2799 0 -2.0 1e-06 
0.0 1.28 0 -2.0 1e-06 
0.0 1.2801 0 -2.0 1e-06 
0.0 1.2802 0 -2.0 1e-06 
0.0 1.2803 0 -2.0 1e-06 
0.0 1.2804 0 -2.0 1e-06 
0.0 1.2805 0 -2.0 1e-06 
0.0 1.2806 0 -2.0 1e-06 
0.0 1.2807 0 -2.0 1e-06 
0.0 1.2808 0 -2.0 1e-06 
0.0 1.2809 0 -2.0 1e-06 
0.0 1.281 0 -2.0 1e-06 
0.0 1.2811 0 -2.0 1e-06 
0.0 1.2812 0 -2.0 1e-06 
0.0 1.2813 0 -2.0 1e-06 
0.0 1.2814 0 -2.0 1e-06 
0.0 1.2815 0 -2.0 1e-06 
0.0 1.2816 0 -2.0 1e-06 
0.0 1.2817 0 -2.0 1e-06 
0.0 1.2818 0 -2.0 1e-06 
0.0 1.2819 0 -2.0 1e-06 
0.0 1.282 0 -2.0 1e-06 
0.0 1.2821 0 -2.0 1e-06 
0.0 1.2822 0 -2.0 1e-06 
0.0 1.2823 0 -2.0 1e-06 
0.0 1.2824 0 -2.0 1e-06 
0.0 1.2825 0 -2.0 1e-06 
0.0 1.2826 0 -2.0 1e-06 
0.0 1.2827 0 -2.0 1e-06 
0.0 1.2828 0 -2.0 1e-06 
0.0 1.2829 0 -2.0 1e-06 
0.0 1.283 0 -2.0 1e-06 
0.0 1.2831 0 -2.0 1e-06 
0.0 1.2832 0 -2.0 1e-06 
0.0 1.2833 0 -2.0 1e-06 
0.0 1.2834 0 -2.0 1e-06 
0.0 1.2835 0 -2.0 1e-06 
0.0 1.2836 0 -2.0 1e-06 
0.0 1.2837 0 -2.0 1e-06 
0.0 1.2838 0 -2.0 1e-06 
0.0 1.2839 0 -2.0 1e-06 
0.0 1.284 0 -2.0 1e-06 
0.0 1.2841 0 -2.0 1e-06 
0.0 1.2842 0 -2.0 1e-06 
0.0 1.2843 0 -2.0 1e-06 
0.0 1.2844 0 -2.0 1e-06 
0.0 1.2845 0 -2.0 1e-06 
0.0 1.2846 0 -2.0 1e-06 
0.0 1.2847 0 -2.0 1e-06 
0.0 1.2848 0 -2.0 1e-06 
0.0 1.2849 0 -2.0 1e-06 
0.0 1.285 0 -2.0 1e-06 
0.0 1.2851 0 -2.0 1e-06 
0.0 1.2852 0 -2.0 1e-06 
0.0 1.2853 0 -2.0 1e-06 
0.0 1.2854 0 -2.0 1e-06 
0.0 1.2855 0 -2.0 1e-06 
0.0 1.2856 0 -2.0 1e-06 
0.0 1.2857 0 -2.0 1e-06 
0.0 1.2858 0 -2.0 1e-06 
0.0 1.2859 0 -2.0 1e-06 
0.0 1.286 0 -2.0 1e-06 
0.0 1.2861 0 -2.0 1e-06 
0.0 1.2862 0 -2.0 1e-06 
0.0 1.2863 0 -2.0 1e-06 
0.0 1.2864 0 -2.0 1e-06 
0.0 1.2865 0 -2.0 1e-06 
0.0 1.2866 0 -2.0 1e-06 
0.0 1.2867 0 -2.0 1e-06 
0.0 1.2868 0 -2.0 1e-06 
0.0 1.2869 0 -2.0 1e-06 
0.0 1.287 0 -2.0 1e-06 
0.0 1.2871 0 -2.0 1e-06 
0.0 1.2872 0 -2.0 1e-06 
0.0 1.2873 0 -2.0 1e-06 
0.0 1.2874 0 -2.0 1e-06 
0.0 1.2875 0 -2.0 1e-06 
0.0 1.2876 0 -2.0 1e-06 
0.0 1.2877 0 -2.0 1e-06 
0.0 1.2878 0 -2.0 1e-06 
0.0 1.2879 0 -2.0 1e-06 
0.0 1.288 0 -2.0 1e-06 
0.0 1.2881 0 -2.0 1e-06 
0.0 1.2882 0 -2.0 1e-06 
0.0 1.2883 0 -2.0 1e-06 
0.0 1.2884 0 -2.0 1e-06 
0.0 1.2885 0 -2.0 1e-06 
0.0 1.2886 0 -2.0 1e-06 
0.0 1.2887 0 -2.0 1e-06 
0.0 1.2888 0 -2.0 1e-06 
0.0 1.2889 0 -2.0 1e-06 
0.0 1.289 0 -2.0 1e-06 
0.0 1.2891 0 -2.0 1e-06 
0.0 1.2892 0 -2.0 1e-06 
0.0 1.2893 0 -2.0 1e-06 
0.0 1.2894 0 -2.0 1e-06 
0.0 1.2895 0 -2.0 1e-06 
0.0 1.2896 0 -2.0 1e-06 
0.0 1.2897 0 -2.0 1e-06 
0.0 1.2898 0 -2.0 1e-06 
0.0 1.2899 0 -2.0 1e-06 
0.0 1.29 0 -2.0 1e-06 
0.0 1.2901 0 -2.0 1e-06 
0.0 1.2902 0 -2.0 1e-06 
0.0 1.2903 0 -2.0 1e-06 
0.0 1.2904 0 -2.0 1e-06 
0.0 1.2905 0 -2.0 1e-06 
0.0 1.2906 0 -2.0 1e-06 
0.0 1.2907 0 -2.0 1e-06 
0.0 1.2908 0 -2.0 1e-06 
0.0 1.2909 0 -2.0 1e-06 
0.0 1.291 0 -2.0 1e-06 
0.0 1.2911 0 -2.0 1e-06 
0.0 1.2912 0 -2.0 1e-06 
0.0 1.2913 0 -2.0 1e-06 
0.0 1.2914 0 -2.0 1e-06 
0.0 1.2915 0 -2.0 1e-06 
0.0 1.2916 0 -2.0 1e-06 
0.0 1.2917 0 -2.0 1e-06 
0.0 1.2918 0 -2.0 1e-06 
0.0 1.2919 0 -2.0 1e-06 
0.0 1.292 0 -2.0 1e-06 
0.0 1.2921 0 -2.0 1e-06 
0.0 1.2922 0 -2.0 1e-06 
0.0 1.2923 0 -2.0 1e-06 
0.0 1.2924 0 -2.0 1e-06 
0.0 1.2925 0 -2.0 1e-06 
0.0 1.2926 0 -2.0 1e-06 
0.0 1.2927 0 -2.0 1e-06 
0.0 1.2928 0 -2.0 1e-06 
0.0 1.2929 0 -2.0 1e-06 
0.0 1.293 0 -2.0 1e-06 
0.0 1.2931 0 -2.0 1e-06 
0.0 1.2932 0 -2.0 1e-06 
0.0 1.2933 0 -2.0 1e-06 
0.0 1.2934 0 -2.0 1e-06 
0.0 1.2935 0 -2.0 1e-06 
0.0 1.2936 0 -2.0 1e-06 
0.0 1.2937 0 -2.0 1e-06 
0.0 1.2938 0 -2.0 1e-06 
0.0 1.2939 0 -2.0 1e-06 
0.0 1.294 0 -2.0 1e-06 
0.0 1.2941 0 -2.0 1e-06 
0.0 1.2942 0 -2.0 1e-06 
0.0 1.2943 0 -2.0 1e-06 
0.0 1.2944 0 -2.0 1e-06 
0.0 1.2945 0 -2.0 1e-06 
0.0 1.2946 0 -2.0 1e-06 
0.0 1.2947 0 -2.0 1e-06 
0.0 1.2948 0 -2.0 1e-06 
0.0 1.2949 0 -2.0 1e-06 
0.0 1.295 0 -2.0 1e-06 
0.0 1.2951 0 -2.0 1e-06 
0.0 1.2952 0 -2.0 1e-06 
0.0 1.2953 0 -2.0 1e-06 
0.0 1.2954 0 -2.0 1e-06 
0.0 1.2955 0 -2.0 1e-06 
0.0 1.2956 0 -2.0 1e-06 
0.0 1.2957 0 -2.0 1e-06 
0.0 1.2958 0 -2.0 1e-06 
0.0 1.2959 0 -2.0 1e-06 
0.0 1.296 0 -2.0 1e-06 
0.0 1.2961 0 -2.0 1e-06 
0.0 1.2962 0 -2.0 1e-06 
0.0 1.2963 0 -2.0 1e-06 
0.0 1.2964 0 -2.0 1e-06 
0.0 1.2965 0 -2.0 1e-06 
0.0 1.2966 0 -2.0 1e-06 
0.0 1.2967 0 -2.0 1e-06 
0.0 1.2968 0 -2.0 1e-06 
0.0 1.2969 0 -2.0 1e-06 
0.0 1.297 0 -2.0 1e-06 
0.0 1.2971 0 -2.0 1e-06 
0.0 1.2972 0 -2.0 1e-06 
0.0 1.2973 0 -2.0 1e-06 
0.0 1.2974 0 -2.0 1e-06 
0.0 1.2975 0 -2.0 1e-06 
0.0 1.2976 0 -2.0 1e-06 
0.0 1.2977 0 -2.0 1e-06 
0.0 1.2978 0 -2.0 1e-06 
0.0 1.2979 0 -2.0 1e-06 
0.0 1.298 0 -2.0 1e-06 
0.0 1.2981 0 -2.0 1e-06 
0.0 1.2982 0 -2.0 1e-06 
0.0 1.2983 0 -2.0 1e-06 
0.0 1.2984 0 -2.0 1e-06 
0.0 1.2985 0 -2.0 1e-06 
0.0 1.2986 0 -2.0 1e-06 
0.0 1.2987 0 -2.0 1e-06 
0.0 1.2988 0 -2.0 1e-06 
0.0 1.2989 0 -2.0 1e-06 
0.0 1.299 0 -2.0 1e-06 
0.0 1.2991 0 -2.0 1e-06 
0.0 1.2992 0 -2.0 1e-06 
0.0 1.2993 0 -2.0 1e-06 
0.0 1.2994 0 -2.0 1e-06 
0.0 1.2995 0 -2.0 1e-06 
0.0 1.2996 0 -2.0 1e-06 
0.0 1.2997 0 -2.0 1e-06 
0.0 1.2998 0 -2.0 1e-06 
0.0 1.2999 0 -2.0 1e-06 
0.0 1.3 0 -2.0 1e-06 
0.0 1.3001 0 -2.0 1e-06 
0.0 1.3002 0 -2.0 1e-06 
0.0 1.3003 0 -2.0 1e-06 
0.0 1.3004 0 -2.0 1e-06 
0.0 1.3005 0 -2.0 1e-06 
0.0 1.3006 0 -2.0 1e-06 
0.0 1.3007 0 -2.0 1e-06 
0.0 1.3008 0 -2.0 1e-06 
0.0 1.3009 0 -2.0 1e-06 
0.0 1.301 0 -2.0 1e-06 
0.0 1.3011 0 -2.0 1e-06 
0.0 1.3012 0 -2.0 1e-06 
0.0 1.3013 0 -2.0 1e-06 
0.0 1.3014 0 -2.0 1e-06 
0.0 1.3015 0 -2.0 1e-06 
0.0 1.3016 0 -2.0 1e-06 
0.0 1.3017 0 -2.0 1e-06 
0.0 1.3018 0 -2.0 1e-06 
0.0 1.3019 0 -2.0 1e-06 
0.0 1.302 0 -2.0 1e-06 
0.0 1.3021 0 -2.0 1e-06 
0.0 1.3022 0 -2.0 1e-06 
0.0 1.3023 0 -2.0 1e-06 
0.0 1.3024 0 -2.0 1e-06 
0.0 1.3025 0 -2.0 1e-06 
0.0 1.3026 0 -2.0 1e-06 
0.0 1.3027 0 -2.0 1e-06 
0.0 1.3028 0 -2.0 1e-06 
0.0 1.3029 0 -2.0 1e-06 
0.0 1.303 0 -2.0 1e-06 
0.0 1.3031 0 -2.0 1e-06 
0.0 1.3032 0 -2.0 1e-06 
0.0 1.3033 0 -2.0 1e-06 
0.0 1.3034 0 -2.0 1e-06 
0.0 1.3035 0 -2.0 1e-06 
0.0 1.3036 0 -2.0 1e-06 
0.0 1.3037 0 -2.0 1e-06 
0.0 1.3038 0 -2.0 1e-06 
0.0 1.3039 0 -2.0 1e-06 
0.0 1.304 0 -2.0 1e-06 
0.0 1.3041 0 -2.0 1e-06 
0.0 1.3042 0 -2.0 1e-06 
0.0 1.3043 0 -2.0 1e-06 
0.0 1.3044 0 -2.0 1e-06 
0.0 1.3045 0 -2.0 1e-06 
0.0 1.3046 0 -2.0 1e-06 
0.0 1.3047 0 -2.0 1e-06 
0.0 1.3048 0 -2.0 1e-06 
0.0 1.3049 0 -2.0 1e-06 
0.0 1.305 0 -2.0 1e-06 
0.0 1.3051 0 -2.0 1e-06 
0.0 1.3052 0 -2.0 1e-06 
0.0 1.3053 0 -2.0 1e-06 
0.0 1.3054 0 -2.0 1e-06 
0.0 1.3055 0 -2.0 1e-06 
0.0 1.3056 0 -2.0 1e-06 
0.0 1.3057 0 -2.0 1e-06 
0.0 1.3058 0 -2.0 1e-06 
0.0 1.3059 0 -2.0 1e-06 
0.0 1.306 0 -2.0 1e-06 
0.0 1.3061 0 -2.0 1e-06 
0.0 1.3062 0 -2.0 1e-06 
0.0 1.3063 0 -2.0 1e-06 
0.0 1.3064 0 -2.0 1e-06 
0.0 1.3065 0 -2.0 1e-06 
0.0 1.3066 0 -2.0 1e-06 
0.0 1.3067 0 -2.0 1e-06 
0.0 1.3068 0 -2.0 1e-06 
0.0 1.3069 0 -2.0 1e-06 
0.0 1.307 0 -2.0 1e-06 
0.0 1.3071 0 -2.0 1e-06 
0.0 1.3072 0 -2.0 1e-06 
0.0 1.3073 0 -2.0 1e-06 
0.0 1.3074 0 -2.0 1e-06 
0.0 1.3075 0 -2.0 1e-06 
0.0 1.3076 0 -2.0 1e-06 
0.0 1.3077 0 -2.0 1e-06 
0.0 1.3078 0 -2.0 1e-06 
0.0 1.3079 0 -2.0 1e-06 
0.0 1.308 0 -2.0 1e-06 
0.0 1.3081 0 -2.0 1e-06 
0.0 1.3082 0 -2.0 1e-06 
0.0 1.3083 0 -2.0 1e-06 
0.0 1.3084 0 -2.0 1e-06 
0.0 1.3085 0 -2.0 1e-06 
0.0 1.3086 0 -2.0 1e-06 
0.0 1.3087 0 -2.0 1e-06 
0.0 1.3088 0 -2.0 1e-06 
0.0 1.3089 0 -2.0 1e-06 
0.0 1.309 0 -2.0 1e-06 
0.0 1.3091 0 -2.0 1e-06 
0.0 1.3092 0 -2.0 1e-06 
0.0 1.3093 0 -2.0 1e-06 
0.0 1.3094 0 -2.0 1e-06 
0.0 1.3095 0 -2.0 1e-06 
0.0 1.3096 0 -2.0 1e-06 
0.0 1.3097 0 -2.0 1e-06 
0.0 1.3098 0 -2.0 1e-06 
0.0 1.3099 0 -2.0 1e-06 
0.0 1.31 0 -2.0 1e-06 
0.0 1.3101 0 -2.0 1e-06 
0.0 1.3102 0 -2.0 1e-06 
0.0 1.3103 0 -2.0 1e-06 
0.0 1.3104 0 -2.0 1e-06 
0.0 1.3105 0 -2.0 1e-06 
0.0 1.3106 0 -2.0 1e-06 
0.0 1.3107 0 -2.0 1e-06 
0.0 1.3108 0 -2.0 1e-06 
0.0 1.3109 0 -2.0 1e-06 
0.0 1.311 0 -2.0 1e-06 
0.0 1.3111 0 -2.0 1e-06 
0.0 1.3112 0 -2.0 1e-06 
0.0 1.3113 0 -2.0 1e-06 
0.0 1.3114 0 -2.0 1e-06 
0.0 1.3115 0 -2.0 1e-06 
0.0 1.3116 0 -2.0 1e-06 
0.0 1.3117 0 -2.0 1e-06 
0.0 1.3118 0 -2.0 1e-06 
0.0 1.3119 0 -2.0 1e-06 
0.0 1.312 0 -2.0 1e-06 
0.0 1.3121 0 -2.0 1e-06 
0.0 1.3122 0 -2.0 1e-06 
0.0 1.3123 0 -2.0 1e-06 
0.0 1.3124 0 -2.0 1e-06 
0.0 1.3125 0 -2.0 1e-06 
0.0 1.3126 0 -2.0 1e-06 
0.0 1.3127 0 -2.0 1e-06 
0.0 1.3128 0 -2.0 1e-06 
0.0 1.3129 0 -2.0 1e-06 
0.0 1.313 0 -2.0 1e-06 
0.0 1.3131 0 -2.0 1e-06 
0.0 1.3132 0 -2.0 1e-06 
0.0 1.3133 0 -2.0 1e-06 
0.0 1.3134 0 -2.0 1e-06 
0.0 1.3135 0 -2.0 1e-06 
0.0 1.3136 0 -2.0 1e-06 
0.0 1.3137 0 -2.0 1e-06 
0.0 1.3138 0 -2.0 1e-06 
0.0 1.3139 0 -2.0 1e-06 
0.0 1.314 0 -2.0 1e-06 
0.0 1.3141 0 -2.0 1e-06 
0.0 1.3142 0 -2.0 1e-06 
0.0 1.3143 0 -2.0 1e-06 
0.0 1.3144 0 -2.0 1e-06 
0.0 1.3145 0 -2.0 1e-06 
0.0 1.3146 0 -2.0 1e-06 
0.0 1.3147 0 -2.0 1e-06 
0.0 1.3148 0 -2.0 1e-06 
0.0 1.3149 0 -2.0 1e-06 
0.0 1.315 0 -2.0 1e-06 
0.0 1.3151 0 -2.0 1e-06 
0.0 1.3152 0 -2.0 1e-06 
0.0 1.3153 0 -2.0 1e-06 
0.0 1.3154 0 -2.0 1e-06 
0.0 1.3155 0 -2.0 1e-06 
0.0 1.3156 0 -2.0 1e-06 
0.0 1.3157 0 -2.0 1e-06 
0.0 1.3158 0 -2.0 1e-06 
0.0 1.3159 0 -2.0 1e-06 
0.0 1.316 0 -2.0 1e-06 
0.0 1.3161 0 -2.0 1e-06 
0.0 1.3162 0 -2.0 1e-06 
0.0 1.3163 0 -2.0 1e-06 
0.0 1.3164 0 -2.0 1e-06 
0.0 1.3165 0 -2.0 1e-06 
0.0 1.3166 0 -2.0 1e-06 
0.0 1.3167 0 -2.0 1e-06 
0.0 1.3168 0 -2.0 1e-06 
0.0 1.3169 0 -2.0 1e-06 
0.0 1.317 0 -2.0 1e-06 
0.0 1.3171 0 -2.0 1e-06 
0.0 1.3172 0 -2.0 1e-06 
0.0 1.3173 0 -2.0 1e-06 
0.0 1.3174 0 -2.0 1e-06 
0.0 1.3175 0 -2.0 1e-06 
0.0 1.3176 0 -2.0 1e-06 
0.0 1.3177 0 -2.0 1e-06 
0.0 1.3178 0 -2.0 1e-06 
0.0 1.3179 0 -2.0 1e-06 
0.0 1.318 0 -2.0 1e-06 
0.0 1.3181 0 -2.0 1e-06 
0.0 1.3182 0 -2.0 1e-06 
0.0 1.3183 0 -2.0 1e-06 
0.0 1.3184 0 -2.0 1e-06 
0.0 1.3185 0 -2.0 1e-06 
0.0 1.3186 0 -2.0 1e-06 
0.0 1.3187 0 -2.0 1e-06 
0.0 1.3188 0 -2.0 1e-06 
0.0 1.3189 0 -2.0 1e-06 
0.0 1.319 0 -2.0 1e-06 
0.0 1.3191 0 -2.0 1e-06 
0.0 1.3192 0 -2.0 1e-06 
0.0 1.3193 0 -2.0 1e-06 
0.0 1.3194 0 -2.0 1e-06 
0.0 1.3195 0 -2.0 1e-06 
0.0 1.3196 0 -2.0 1e-06 
0.0 1.3197 0 -2.0 1e-06 
0.0 1.3198 0 -2.0 1e-06 
0.0 1.3199 0 -2.0 1e-06 
0.0 1.32 0 -2.0 1e-06 
0.0 1.3201 0 -2.0 1e-06 
0.0 1.3202 0 -2.0 1e-06 
0.0 1.3203 0 -2.0 1e-06 
0.0 1.3204 0 -2.0 1e-06 
0.0 1.3205 0 -2.0 1e-06 
0.0 1.3206 0 -2.0 1e-06 
0.0 1.3207 0 -2.0 1e-06 
0.0 1.3208 0 -2.0 1e-06 
0.0 1.3209 0 -2.0 1e-06 
0.0 1.321 0 -2.0 1e-06 
0.0 1.3211 0 -2.0 1e-06 
0.0 1.3212 0 -2.0 1e-06 
0.0 1.3213 0 -2.0 1e-06 
0.0 1.3214 0 -2.0 1e-06 
0.0 1.3215 0 -2.0 1e-06 
0.0 1.3216 0 -2.0 1e-06 
0.0 1.3217 0 -2.0 1e-06 
0.0 1.3218 0 -2.0 1e-06 
0.0 1.3219 0 -2.0 1e-06 
0.0 1.322 0 -2.0 1e-06 
0.0 1.3221 0 -2.0 1e-06 
0.0 1.3222 0 -2.0 1e-06 
0.0 1.3223 0 -2.0 1e-06 
0.0 1.3224 0 -2.0 1e-06 
0.0 1.3225 0 -2.0 1e-06 
0.0 1.3226 0 -2.0 1e-06 
0.0 1.3227 0 -2.0 1e-06 
0.0 1.3228 0 -2.0 1e-06 
0.0 1.3229 0 -2.0 1e-06 
0.0 1.323 0 -2.0 1e-06 
0.0 1.3231 0 -2.0 1e-06 
0.0 1.3232 0 -2.0 1e-06 
0.0 1.3233 0 -2.0 1e-06 
0.0 1.3234 0 -2.0 1e-06 
0.0 1.3235 0 -2.0 1e-06 
0.0 1.3236 0 -2.0 1e-06 
0.0 1.3237 0 -2.0 1e-06 
0.0 1.3238 0 -2.0 1e-06 
0.0 1.3239 0 -2.0 1e-06 
0.0 1.324 0 -2.0 1e-06 
0.0 1.3241 0 -2.0 1e-06 
0.0 1.3242 0 -2.0 1e-06 
0.0 1.3243 0 -2.0 1e-06 
0.0 1.3244 0 -2.0 1e-06 
0.0 1.3245 0 -2.0 1e-06 
0.0 1.3246 0 -2.0 1e-06 
0.0 1.3247 0 -2.0 1e-06 
0.0 1.3248 0 -2.0 1e-06 
0.0 1.3249 0 -2.0 1e-06 
0.0 1.325 0 -2.0 1e-06 
0.0 1.3251 0 -2.0 1e-06 
0.0 1.3252 0 -2.0 1e-06 
0.0 1.3253 0 -2.0 1e-06 
0.0 1.3254 0 -2.0 1e-06 
0.0 1.3255 0 -2.0 1e-06 
0.0 1.3256 0 -2.0 1e-06 
0.0 1.3257 0 -2.0 1e-06 
0.0 1.3258 0 -2.0 1e-06 
0.0 1.3259 0 -2.0 1e-06 
0.0 1.326 0 -2.0 1e-06 
0.0 1.3261 0 -2.0 1e-06 
0.0 1.3262 0 -2.0 1e-06 
0.0 1.3263 0 -2.0 1e-06 
0.0 1.3264 0 -2.0 1e-06 
0.0 1.3265 0 -2.0 1e-06 
0.0 1.3266 0 -2.0 1e-06 
0.0 1.3267 0 -2.0 1e-06 
0.0 1.3268 0 -2.0 1e-06 
0.0 1.3269 0 -2.0 1e-06 
0.0 1.327 0 -2.0 1e-06 
0.0 1.3271 0 -2.0 1e-06 
0.0 1.3272 0 -2.0 1e-06 
0.0 1.3273 0 -2.0 1e-06 
0.0 1.3274 0 -2.0 1e-06 
0.0 1.3275 0 -2.0 1e-06 
0.0 1.3276 0 -2.0 1e-06 
0.0 1.3277 0 -2.0 1e-06 
0.0 1.3278 0 -2.0 1e-06 
0.0 1.3279 0 -2.0 1e-06 
0.0 1.328 0 -2.0 1e-06 
0.0 1.3281 0 -2.0 1e-06 
0.0 1.3282 0 -2.0 1e-06 
0.0 1.3283 0 -2.0 1e-06 
0.0 1.3284 0 -2.0 1e-06 
0.0 1.3285 0 -2.0 1e-06 
0.0 1.3286 0 -2.0 1e-06 
0.0 1.3287 0 -2.0 1e-06 
0.0 1.3288 0 -2.0 1e-06 
0.0 1.3289 0 -2.0 1e-06 
0.0 1.329 0 -2.0 1e-06 
0.0 1.3291 0 -2.0 1e-06 
0.0 1.3292 0 -2.0 1e-06 
0.0 1.3293 0 -2.0 1e-06 
0.0 1.3294 0 -2.0 1e-06 
0.0 1.3295 0 -2.0 1e-06 
0.0 1.3296 0 -2.0 1e-06 
0.0 1.3297 0 -2.0 1e-06 
0.0 1.3298 0 -2.0 1e-06 
0.0 1.3299 0 -2.0 1e-06 
0.0 1.33 0 -2.0 1e-06 
0.0 1.3301 0 -2.0 1e-06 
0.0 1.3302 0 -2.0 1e-06 
0.0 1.3303 0 -2.0 1e-06 
0.0 1.3304 0 -2.0 1e-06 
0.0 1.3305 0 -2.0 1e-06 
0.0 1.3306 0 -2.0 1e-06 
0.0 1.3307 0 -2.0 1e-06 
0.0 1.3308 0 -2.0 1e-06 
0.0 1.3309 0 -2.0 1e-06 
0.0 1.331 0 -2.0 1e-06 
0.0 1.3311 0 -2.0 1e-06 
0.0 1.3312 0 -2.0 1e-06 
0.0 1.3313 0 -2.0 1e-06 
0.0 1.3314 0 -2.0 1e-06 
0.0 1.3315 0 -2.0 1e-06 
0.0 1.3316 0 -2.0 1e-06 
0.0 1.3317 0 -2.0 1e-06 
0.0 1.3318 0 -2.0 1e-06 
0.0 1.3319 0 -2.0 1e-06 
0.0 1.332 0 -2.0 1e-06 
0.0 1.3321 0 -2.0 1e-06 
0.0 1.3322 0 -2.0 1e-06 
0.0 1.3323 0 -2.0 1e-06 
0.0 1.3324 0 -2.0 1e-06 
0.0 1.3325 0 -2.0 1e-06 
0.0 1.3326 0 -2.0 1e-06 
0.0 1.3327 0 -2.0 1e-06 
0.0 1.3328 0 -2.0 1e-06 
0.0 1.3329 0 -2.0 1e-06 
0.0 1.333 0 -2.0 1e-06 
0.0 1.3331 0 -2.0 1e-06 
0.0 1.3332 0 -2.0 1e-06 
0.0 1.3333 0 -2.0 1e-06 
0.0 1.3334 0 -2.0 1e-06 
0.0 1.3335 0 -2.0 1e-06 
0.0 1.3336 0 -2.0 1e-06 
0.0 1.3337 0 -2.0 1e-06 
0.0 1.3338 0 -2.0 1e-06 
0.0 1.3339 0 -2.0 1e-06 
0.0 1.334 0 -2.0 1e-06 
0.0 1.3341 0 -2.0 1e-06 
0.0 1.3342 0 -2.0 1e-06 
0.0 1.3343 0 -2.0 1e-06 
0.0 1.3344 0 -2.0 1e-06 
0.0 1.3345 0 -2.0 1e-06 
0.0 1.3346 0 -2.0 1e-06 
0.0 1.3347 0 -2.0 1e-06 
0.0 1.3348 0 -2.0 1e-06 
0.0 1.3349 0 -2.0 1e-06 
0.0 1.335 0 -2.0 1e-06 
0.0 1.3351 0 -2.0 1e-06 
0.0 1.3352 0 -2.0 1e-06 
0.0 1.3353 0 -2.0 1e-06 
0.0 1.3354 0 -2.0 1e-06 
0.0 1.3355 0 -2.0 1e-06 
0.0 1.3356 0 -2.0 1e-06 
0.0 1.3357 0 -2.0 1e-06 
0.0 1.3358 0 -2.0 1e-06 
0.0 1.3359 0 -2.0 1e-06 
0.0 1.336 0 -2.0 1e-06 
0.0 1.3361 0 -2.0 1e-06 
0.0 1.3362 0 -2.0 1e-06 
0.0 1.3363 0 -2.0 1e-06 
0.0 1.3364 0 -2.0 1e-06 
0.0 1.3365 0 -2.0 1e-06 
0.0 1.3366 0 -2.0 1e-06 
0.0 1.3367 0 -2.0 1e-06 
0.0 1.3368 0 -2.0 1e-06 
0.0 1.3369 0 -2.0 1e-06 
0.0 1.337 0 -2.0 1e-06 
0.0 1.3371 0 -2.0 1e-06 
0.0 1.3372 0 -2.0 1e-06 
0.0 1.3373 0 -2.0 1e-06 
0.0 1.3374 0 -2.0 1e-06 
0.0 1.3375 0 -2.0 1e-06 
0.0 1.3376 0 -2.0 1e-06 
0.0 1.3377 0 -2.0 1e-06 
0.0 1.3378 0 -2.0 1e-06 
0.0 1.3379 0 -2.0 1e-06 
0.0 1.338 0 -2.0 1e-06 
0.0 1.3381 0 -2.0 1e-06 
0.0 1.3382 0 -2.0 1e-06 
0.0 1.3383 0 -2.0 1e-06 
0.0 1.3384 0 -2.0 1e-06 
0.0 1.3385 0 -2.0 1e-06 
0.0 1.3386 0 -2.0 1e-06 
0.0 1.3387 0 -2.0 1e-06 
0.0 1.3388 0 -2.0 1e-06 
0.0 1.3389 0 -2.0 1e-06 
0.0 1.339 0 -2.0 1e-06 
0.0 1.3391 0 -2.0 1e-06 
0.0 1.3392 0 -2.0 1e-06 
0.0 1.3393 0 -2.0 1e-06 
0.0 1.3394 0 -2.0 1e-06 
0.0 1.3395 0 -2.0 1e-06 
0.0 1.3396 0 -2.0 1e-06 
0.0 1.3397 0 -2.0 1e-06 
0.0 1.3398 0 -2.0 1e-06 
0.0 1.3399 0 -2.0 1e-06 
0.0 1.34 0 -2.0 1e-06 
0.0 1.3401 0 -2.0 1e-06 
0.0 1.3402 0 -2.0 1e-06 
0.0 1.3403 0 -2.0 1e-06 
0.0 1.3404 0 -2.0 1e-06 
0.0 1.3405 0 -2.0 1e-06 
0.0 1.3406 0 -2.0 1e-06 
0.0 1.3407 0 -2.0 1e-06 
0.0 1.3408 0 -2.0 1e-06 
0.0 1.3409 0 -2.0 1e-06 
0.0 1.341 0 -2.0 1e-06 
0.0 1.3411 0 -2.0 1e-06 
0.0 1.3412 0 -2.0 1e-06 
0.0 1.3413 0 -2.0 1e-06 
0.0 1.3414 0 -2.0 1e-06 
0.0 1.3415 0 -2.0 1e-06 
0.0 1.3416 0 -2.0 1e-06 
0.0 1.3417 0 -2.0 1e-06 
0.0 1.3418 0 -2.0 1e-06 
0.0 1.3419 0 -2.0 1e-06 
0.0 1.342 0 -2.0 1e-06 
0.0 1.3421 0 -2.0 1e-06 
0.0 1.3422 0 -2.0 1e-06 
0.0 1.3423 0 -2.0 1e-06 
0.0 1.3424 0 -2.0 1e-06 
0.0 1.3425 0 -2.0 1e-06 
0.0 1.3426 0 -2.0 1e-06 
0.0 1.3427 0 -2.0 1e-06 
0.0 1.3428 0 -2.0 1e-06 
0.0 1.3429 0 -2.0 1e-06 
0.0 1.343 0 -2.0 1e-06 
0.0 1.3431 0 -2.0 1e-06 
0.0 1.3432 0 -2.0 1e-06 
0.0 1.3433 0 -2.0 1e-06 
0.0 1.3434 0 -2.0 1e-06 
0.0 1.3435 0 -2.0 1e-06 
0.0 1.3436 0 -2.0 1e-06 
0.0 1.3437 0 -2.0 1e-06 
0.0 1.3438 0 -2.0 1e-06 
0.0 1.3439 0 -2.0 1e-06 
0.0 1.344 0 -2.0 1e-06 
0.0 1.3441 0 -2.0 1e-06 
0.0 1.3442 0 -2.0 1e-06 
0.0 1.3443 0 -2.0 1e-06 
0.0 1.3444 0 -2.0 1e-06 
0.0 1.3445 0 -2.0 1e-06 
0.0 1.3446 0 -2.0 1e-06 
0.0 1.3447 0 -2.0 1e-06 
0.0 1.3448 0 -2.0 1e-06 
0.0 1.3449 0 -2.0 1e-06 
0.0 1.345 0 -2.0 1e-06 
0.0 1.3451 0 -2.0 1e-06 
0.0 1.3452 0 -2.0 1e-06 
0.0 1.3453 0 -2.0 1e-06 
0.0 1.3454 0 -2.0 1e-06 
0.0 1.3455 0 -2.0 1e-06 
0.0 1.3456 0 -2.0 1e-06 
0.0 1.3457 0 -2.0 1e-06 
0.0 1.3458 0 -2.0 1e-06 
0.0 1.3459 0 -2.0 1e-06 
0.0 1.346 0 -2.0 1e-06 
0.0 1.3461 0 -2.0 1e-06 
0.0 1.3462 0 -2.0 1e-06 
0.0 1.3463 0 -2.0 1e-06 
0.0 1.3464 0 -2.0 1e-06 
0.0 1.3465 0 -2.0 1e-06 
0.0 1.3466 0 -2.0 1e-06 
0.0 1.3467 0 -2.0 1e-06 
0.0 1.3468 0 -2.0 1e-06 
0.0 1.3469 0 -2.0 1e-06 
0.0 1.347 0 -2.0 1e-06 
0.0 1.3471 0 -2.0 1e-06 
0.0 1.3472 0 -2.0 1e-06 
0.0 1.3473 0 -2.0 1e-06 
0.0 1.3474 0 -2.0 1e-06 
0.0 1.3475 0 -2.0 1e-06 
0.0 1.3476 0 -2.0 1e-06 
0.0 1.3477 0 -2.0 1e-06 
0.0 1.3478 0 -2.0 1e-06 
0.0 1.3479 0 -2.0 1e-06 
0.0 1.348 0 -2.0 1e-06 
0.0 1.3481 0 -2.0 1e-06 
0.0 1.3482 0 -2.0 1e-06 
0.0 1.3483 0 -2.0 1e-06 
0.0 1.3484 0 -2.0 1e-06 
0.0 1.3485 0 -2.0 1e-06 
0.0 1.3486 0 -2.0 1e-06 
0.0 1.3487 0 -2.0 1e-06 
0.0 1.3488 0 -2.0 1e-06 
0.0 1.3489 0 -2.0 1e-06 
0.0 1.349 0 -2.0 1e-06 
0.0 1.3491 0 -2.0 1e-06 
0.0 1.3492 0 -2.0 1e-06 
0.0 1.3493 0 -2.0 1e-06 
0.0 1.3494 0 -2.0 1e-06 
0.0 1.3495 0 -2.0 1e-06 
0.0 1.3496 0 -2.0 1e-06 
0.0 1.3497 0 -2.0 1e-06 
0.0 1.3498 0 -2.0 1e-06 
0.0 1.3499 0 -2.0 1e-06 
0.0 1.35 0 -2.0 1e-06 
0.0 1.3501 0 -2.0 1e-06 
0.0 1.3502 0 -2.0 1e-06 
0.0 1.3503 0 -2.0 1e-06 
0.0 1.3504 0 -2.0 1e-06 
0.0 1.3505 0 -2.0 1e-06 
0.0 1.3506 0 -2.0 1e-06 
0.0 1.3507 0 -2.0 1e-06 
0.0 1.3508 0 -2.0 1e-06 
0.0 1.3509 0 -2.0 1e-06 
0.0 1.351 0 -2.0 1e-06 
0.0 1.3511 0 -2.0 1e-06 
0.0 1.3512 0 -2.0 1e-06 
0.0 1.3513 0 -2.0 1e-06 
0.0 1.3514 0 -2.0 1e-06 
0.0 1.3515 0 -2.0 1e-06 
0.0 1.3516 0 -2.0 1e-06 
0.0 1.3517 0 -2.0 1e-06 
0.0 1.3518 0 -2.0 1e-06 
0.0 1.3519 0 -2.0 1e-06 
0.0 1.352 0 -2.0 1e-06 
0.0 1.3521 0 -2.0 1e-06 
0.0 1.3522 0 -2.0 1e-06 
0.0 1.3523 0 -2.0 1e-06 
0.0 1.3524 0 -2.0 1e-06 
0.0 1.3525 0 -2.0 1e-06 
0.0 1.3526 0 -2.0 1e-06 
0.0 1.3527 0 -2.0 1e-06 
0.0 1.3528 0 -2.0 1e-06 
0.0 1.3529 0 -2.0 1e-06 
0.0 1.353 0 -2.0 1e-06 
0.0 1.3531 0 -2.0 1e-06 
0.0 1.3532 0 -2.0 1e-06 
0.0 1.3533 0 -2.0 1e-06 
0.0 1.3534 0 -2.0 1e-06 
0.0 1.3535 0 -2.0 1e-06 
0.0 1.3536 0 -2.0 1e-06 
0.0 1.3537 0 -2.0 1e-06 
0.0 1.3538 0 -2.0 1e-06 
0.0 1.3539 0 -2.0 1e-06 
0.0 1.354 0 -2.0 1e-06 
0.0 1.3541 0 -2.0 1e-06 
0.0 1.3542 0 -2.0 1e-06 
0.0 1.3543 0 -2.0 1e-06 
0.0 1.3544 0 -2.0 1e-06 
0.0 1.3545 0 -2.0 1e-06 
0.0 1.3546 0 -2.0 1e-06 
0.0 1.3547 0 -2.0 1e-06 
0.0 1.3548 0 -2.0 1e-06 
0.0 1.3549 0 -2.0 1e-06 
0.0 1.355 0 -2.0 1e-06 
0.0 1.3551 0 -2.0 1e-06 
0.0 1.3552 0 -2.0 1e-06 
0.0 1.3553 0 -2.0 1e-06 
0.0 1.3554 0 -2.0 1e-06 
0.0 1.3555 0 -2.0 1e-06 
0.0 1.3556 0 -2.0 1e-06 
0.0 1.3557 0 -2.0 1e-06 
0.0 1.3558 0 -2.0 1e-06 
0.0 1.3559 0 -2.0 1e-06 
0.0 1.356 0 -2.0 1e-06 
0.0 1.3561 0 -2.0 1e-06 
0.0 1.3562 0 -2.0 1e-06 
0.0 1.3563 0 -2.0 1e-06 
0.0 1.3564 0 -2.0 1e-06 
0.0 1.3565 0 -2.0 1e-06 
0.0 1.3566 0 -2.0 1e-06 
0.0 1.3567 0 -2.0 1e-06 
0.0 1.3568 0 -2.0 1e-06 
0.0 1.3569 0 -2.0 1e-06 
0.0 1.357 0 -2.0 1e-06 
0.0 1.3571 0 -2.0 1e-06 
0.0 1.3572 0 -2.0 1e-06 
0.0 1.3573 0 -2.0 1e-06 
0.0 1.3574 0 -2.0 1e-06 
0.0 1.3575 0 -2.0 1e-06 
0.0 1.3576 0 -2.0 1e-06 
0.0 1.3577 0 -2.0 1e-06 
0.0 1.3578 0 -2.0 1e-06 
0.0 1.3579 0 -2.0 1e-06 
0.0 1.358 0 -2.0 1e-06 
0.0 1.3581 0 -2.0 1e-06 
0.0 1.3582 0 -2.0 1e-06 
0.0 1.3583 0 -2.0 1e-06 
0.0 1.3584 0 -2.0 1e-06 
0.0 1.3585 0 -2.0 1e-06 
0.0 1.3586 0 -2.0 1e-06 
0.0 1.3587 0 -2.0 1e-06 
0.0 1.3588 0 -2.0 1e-06 
0.0 1.3589 0 -2.0 1e-06 
0.0 1.359 0 -2.0 1e-06 
0.0 1.3591 0 -2.0 1e-06 
0.0 1.3592 0 -2.0 1e-06 
0.0 1.3593 0 -2.0 1e-06 
0.0 1.3594 0 -2.0 1e-06 
0.0 1.3595 0 -2.0 1e-06 
0.0 1.3596 0 -2.0 1e-06 
0.0 1.3597 0 -2.0 1e-06 
0.0 1.3598 0 -2.0 1e-06 
0.0 1.3599 0 -2.0 1e-06 
0.0 1.36 0 -2.0 1e-06 
0.0 1.3601 0 -2.0 1e-06 
0.0 1.3602 0 -2.0 1e-06 
0.0 1.3603 0 -2.0 1e-06 
0.0 1.3604 0 -2.0 1e-06 
0.0 1.3605 0 -2.0 1e-06 
0.0 1.3606 0 -2.0 1e-06 
0.0 1.3607 0 -2.0 1e-06 
0.0 1.3608 0 -2.0 1e-06 
0.0 1.3609 0 -2.0 1e-06 
0.0 1.361 0 -2.0 1e-06 
0.0 1.3611 0 -2.0 1e-06 
0.0 1.3612 0 -2.0 1e-06 
0.0 1.3613 0 -2.0 1e-06 
0.0 1.3614 0 -2.0 1e-06 
0.0 1.3615 0 -2.0 1e-06 
0.0 1.3616 0 -2.0 1e-06 
0.0 1.3617 0 -2.0 1e-06 
0.0 1.3618 0 -2.0 1e-06 
0.0 1.3619 0 -2.0 1e-06 
0.0 1.362 0 -2.0 1e-06 
0.0 1.3621 0 -2.0 1e-06 
0.0 1.3622 0 -2.0 1e-06 
0.0 1.3623 0 -2.0 1e-06 
0.0 1.3624 0 -2.0 1e-06 
0.0 1.3625 0 -2.0 1e-06 
0.0 1.3626 0 -2.0 1e-06 
0.0 1.3627 0 -2.0 1e-06 
0.0 1.3628 0 -2.0 1e-06 
0.0 1.3629 0 -2.0 1e-06 
0.0 1.363 0 -2.0 1e-06 
0.0 1.3631 0 -2.0 1e-06 
0.0 1.3632 0 -2.0 1e-06 
0.0 1.3633 0 -2.0 1e-06 
0.0 1.3634 0 -2.0 1e-06 
0.0 1.3635 0 -2.0 1e-06 
0.0 1.3636 0 -2.0 1e-06 
0.0 1.3637 0 -2.0 1e-06 
0.0 1.3638 0 -2.0 1e-06 
0.0 1.3639 0 -2.0 1e-06 
0.0 1.364 0 -2.0 1e-06 
0.0 1.3641 0 -2.0 1e-06 
0.0 1.3642 0 -2.0 1e-06 
0.0 1.3643 0 -2.0 1e-06 
0.0 1.3644 0 -2.0 1e-06 
0.0 1.3645 0 -2.0 1e-06 
0.0 1.3646 0 -2.0 1e-06 
0.0 1.3647 0 -2.0 1e-06 
0.0 1.3648 0 -2.0 1e-06 
0.0 1.3649 0 -2.0 1e-06 
0.0 1.365 0 -2.0 1e-06 
0.0 1.3651 0 -2.0 1e-06 
0.0 1.3652 0 -2.0 1e-06 
0.0 1.3653 0 -2.0 1e-06 
0.0 1.3654 0 -2.0 1e-06 
0.0 1.3655 0 -2.0 1e-06 
0.0 1.3656 0 -2.0 1e-06 
0.0 1.3657 0 -2.0 1e-06 
0.0 1.3658 0 -2.0 1e-06 
0.0 1.3659 0 -2.0 1e-06 
0.0 1.366 0 -2.0 1e-06 
0.0 1.3661 0 -2.0 1e-06 
0.0 1.3662 0 -2.0 1e-06 
0.0 1.3663 0 -2.0 1e-06 
0.0 1.3664 0 -2.0 1e-06 
0.0 1.3665 0 -2.0 1e-06 
0.0 1.3666 0 -2.0 1e-06 
0.0 1.3667 0 -2.0 1e-06 
0.0 1.3668 0 -2.0 1e-06 
0.0 1.3669 0 -2.0 1e-06 
0.0 1.367 0 -2.0 1e-06 
0.0 1.3671 0 -2.0 1e-06 
0.0 1.3672 0 -2.0 1e-06 
0.0 1.3673 0 -2.0 1e-06 
0.0 1.3674 0 -2.0 1e-06 
0.0 1.3675 0 -2.0 1e-06 
0.0 1.3676 0 -2.0 1e-06 
0.0 1.3677 0 -2.0 1e-06 
0.0 1.3678 0 -2.0 1e-06 
0.0 1.3679 0 -2.0 1e-06 
0.0 1.368 0 -2.0 1e-06 
0.0 1.3681 0 -2.0 1e-06 
0.0 1.3682 0 -2.0 1e-06 
0.0 1.3683 0 -2.0 1e-06 
0.0 1.3684 0 -2.0 1e-06 
0.0 1.3685 0 -2.0 1e-06 
0.0 1.3686 0 -2.0 1e-06 
0.0 1.3687 0 -2.0 1e-06 
0.0 1.3688 0 -2.0 1e-06 
0.0 1.3689 0 -2.0 1e-06 
0.0 1.369 0 -2.0 1e-06 
0.0 1.3691 0 -2.0 1e-06 
0.0 1.3692 0 -2.0 1e-06 
0.0 1.3693 0 -2.0 1e-06 
0.0 1.3694 0 -2.0 1e-06 
0.0 1.3695 0 -2.0 1e-06 
0.0 1.3696 0 -2.0 1e-06 
0.0 1.3697 0 -2.0 1e-06 
0.0 1.3698 0 -2.0 1e-06 
0.0 1.3699 0 -2.0 1e-06 
0.0 1.37 0 -2.0 1e-06 
0.0 1.3701 0 -2.0 1e-06 
0.0 1.3702 0 -2.0 1e-06 
0.0 1.3703 0 -2.0 1e-06 
0.0 1.3704 0 -2.0 1e-06 
0.0 1.3705 0 -2.0 1e-06 
0.0 1.3706 0 -2.0 1e-06 
0.0 1.3707 0 -2.0 1e-06 
0.0 1.3708 0 -2.0 1e-06 
0.0 1.3709 0 -2.0 1e-06 
0.0 1.371 0 -2.0 1e-06 
0.0 1.3711 0 -2.0 1e-06 
0.0 1.3712 0 -2.0 1e-06 
0.0 1.3713 0 -2.0 1e-06 
0.0 1.3714 0 -2.0 1e-06 
0.0 1.3715 0 -2.0 1e-06 
0.0 1.3716 0 -2.0 1e-06 
0.0 1.3717 0 -2.0 1e-06 
0.0 1.3718 0 -2.0 1e-06 
0.0 1.3719 0 -2.0 1e-06 
0.0 1.372 0 -2.0 1e-06 
0.0 1.3721 0 -2.0 1e-06 
0.0 1.3722 0 -2.0 1e-06 
0.0 1.3723 0 -2.0 1e-06 
0.0 1.3724 0 -2.0 1e-06 
0.0 1.3725 0 -2.0 1e-06 
0.0 1.3726 0 -2.0 1e-06 
0.0 1.3727 0 -2.0 1e-06 
0.0 1.3728 0 -2.0 1e-06 
0.0 1.3729 0 -2.0 1e-06 
0.0 1.373 0 -2.0 1e-06 
0.0 1.3731 0 -2.0 1e-06 
0.0 1.3732 0 -2.0 1e-06 
0.0 1.3733 0 -2.0 1e-06 
0.0 1.3734 0 -2.0 1e-06 
0.0 1.3735 0 -2.0 1e-06 
0.0 1.3736 0 -2.0 1e-06 
0.0 1.3737 0 -2.0 1e-06 
0.0 1.3738 0 -2.0 1e-06 
0.0 1.3739 0 -2.0 1e-06 
0.0 1.374 0 -2.0 1e-06 
0.0 1.3741 0 -2.0 1e-06 
0.0 1.3742 0 -2.0 1e-06 
0.0 1.3743 0 -2.0 1e-06 
0.0 1.3744 0 -2.0 1e-06 
0.0 1.3745 0 -2.0 1e-06 
0.0 1.3746 0 -2.0 1e-06 
0.0 1.3747 0 -2.0 1e-06 
0.0 1.3748 0 -2.0 1e-06 
0.0 1.3749 0 -2.0 1e-06 
0.0 1.375 0 -2.0 1e-06 
0.0 1.3751 0 -2.0 1e-06 
0.0 1.3752 0 -2.0 1e-06 
0.0 1.3753 0 -2.0 1e-06 
0.0 1.3754 0 -2.0 1e-06 
0.0 1.3755 0 -2.0 1e-06 
0.0 1.3756 0 -2.0 1e-06 
0.0 1.3757 0 -2.0 1e-06 
0.0 1.3758 0 -2.0 1e-06 
0.0 1.3759 0 -2.0 1e-06 
0.0 1.376 0 -2.0 1e-06 
0.0 1.3761 0 -2.0 1e-06 
0.0 1.3762 0 -2.0 1e-06 
0.0 1.3763 0 -2.0 1e-06 
0.0 1.3764 0 -2.0 1e-06 
0.0 1.3765 0 -2.0 1e-06 
0.0 1.3766 0 -2.0 1e-06 
0.0 1.3767 0 -2.0 1e-06 
0.0 1.3768 0 -2.0 1e-06 
0.0 1.3769 0 -2.0 1e-06 
0.0 1.377 0 -2.0 1e-06 
0.0 1.3771 0 -2.0 1e-06 
0.0 1.3772 0 -2.0 1e-06 
0.0 1.3773 0 -2.0 1e-06 
0.0 1.3774 0 -2.0 1e-06 
0.0 1.3775 0 -2.0 1e-06 
0.0 1.3776 0 -2.0 1e-06 
0.0 1.3777 0 -2.0 1e-06 
0.0 1.3778 0 -2.0 1e-06 
0.0 1.3779 0 -2.0 1e-06 
0.0 1.378 0 -2.0 1e-06 
0.0 1.3781 0 -2.0 1e-06 
0.0 1.3782 0 -2.0 1e-06 
0.0 1.3783 0 -2.0 1e-06 
0.0 1.3784 0 -2.0 1e-06 
0.0 1.3785 0 -2.0 1e-06 
0.0 1.3786 0 -2.0 1e-06 
0.0 1.3787 0 -2.0 1e-06 
0.0 1.3788 0 -2.0 1e-06 
0.0 1.3789 0 -2.0 1e-06 
0.0 1.379 0 -2.0 1e-06 
0.0 1.3791 0 -2.0 1e-06 
0.0 1.3792 0 -2.0 1e-06 
0.0 1.3793 0 -2.0 1e-06 
0.0 1.3794 0 -2.0 1e-06 
0.0 1.3795 0 -2.0 1e-06 
0.0 1.3796 0 -2.0 1e-06 
0.0 1.3797 0 -2.0 1e-06 
0.0 1.3798 0 -2.0 1e-06 
0.0 1.3799 0 -2.0 1e-06 
0.0 1.38 0 -2.0 1e-06 
0.0 1.3801 0 -2.0 1e-06 
0.0 1.3802 0 -2.0 1e-06 
0.0 1.3803 0 -2.0 1e-06 
0.0 1.3804 0 -2.0 1e-06 
0.0 1.3805 0 -2.0 1e-06 
0.0 1.3806 0 -2.0 1e-06 
0.0 1.3807 0 -2.0 1e-06 
0.0 1.3808 0 -2.0 1e-06 
0.0 1.3809 0 -2.0 1e-06 
0.0 1.381 0 -2.0 1e-06 
0.0 1.3811 0 -2.0 1e-06 
0.0 1.3812 0 -2.0 1e-06 
0.0 1.3813 0 -2.0 1e-06 
0.0 1.3814 0 -2.0 1e-06 
0.0 1.3815 0 -2.0 1e-06 
0.0 1.3816 0 -2.0 1e-06 
0.0 1.3817 0 -2.0 1e-06 
0.0 1.3818 0 -2.0 1e-06 
0.0 1.3819 0 -2.0 1e-06 
0.0 1.382 0 -2.0 1e-06 
0.0 1.3821 0 -2.0 1e-06 
0.0 1.3822 0 -2.0 1e-06 
0.0 1.3823 0 -2.0 1e-06 
0.0 1.3824 0 -2.0 1e-06 
0.0 1.3825 0 -2.0 1e-06 
0.0 1.3826 0 -2.0 1e-06 
0.0 1.3827 0 -2.0 1e-06 
0.0 1.3828 0 -2.0 1e-06 
0.0 1.3829 0 -2.0 1e-06 
0.0 1.383 0 -2.0 1e-06 
0.0 1.3831 0 -2.0 1e-06 
0.0 1.3832 0 -2.0 1e-06 
0.0 1.3833 0 -2.0 1e-06 
0.0 1.3834 0 -2.0 1e-06 
0.0 1.3835 0 -2.0 1e-06 
0.0 1.3836 0 -2.0 1e-06 
0.0 1.3837 0 -2.0 1e-06 
0.0 1.3838 0 -2.0 1e-06 
0.0 1.3839 0 -2.0 1e-06 
0.0 1.384 0 -2.0 1e-06 
0.0 1.3841 0 -2.0 1e-06 
0.0 1.3842 0 -2.0 1e-06 
0.0 1.3843 0 -2.0 1e-06 
0.0 1.3844 0 -2.0 1e-06 
0.0 1.3845 0 -2.0 1e-06 
0.0 1.3846 0 -2.0 1e-06 
0.0 1.3847 0 -2.0 1e-06 
0.0 1.3848 0 -2.0 1e-06 
0.0 1.3849 0 -2.0 1e-06 
0.0 1.385 0 -2.0 1e-06 
0.0 1.3851 0 -2.0 1e-06 
0.0 1.3852 0 -2.0 1e-06 
0.0 1.3853 0 -2.0 1e-06 
0.0 1.3854 0 -2.0 1e-06 
0.0 1.3855 0 -2.0 1e-06 
0.0 1.3856 0 -2.0 1e-06 
0.0 1.3857 0 -2.0 1e-06 
0.0 1.3858 0 -2.0 1e-06 
0.0 1.3859 0 -2.0 1e-06 
0.0 1.386 0 -2.0 1e-06 
0.0 1.3861 0 -2.0 1e-06 
0.0 1.3862 0 -2.0 1e-06 
0.0 1.3863 0 -2.0 1e-06 
0.0 1.3864 0 -2.0 1e-06 
0.0 1.3865 0 -2.0 1e-06 
0.0 1.3866 0 -2.0 1e-06 
0.0 1.3867 0 -2.0 1e-06 
0.0 1.3868 0 -2.0 1e-06 
0.0 1.3869 0 -2.0 1e-06 
0.0 1.387 0 -2.0 1e-06 
0.0 1.3871 0 -2.0 1e-06 
0.0 1.3872 0 -2.0 1e-06 
0.0 1.3873 0 -2.0 1e-06 
0.0 1.3874 0 -2.0 1e-06 
0.0 1.3875 0 -2.0 1e-06 
0.0 1.3876 0 -2.0 1e-06 
0.0 1.3877 0 -2.0 1e-06 
0.0 1.3878 0 -2.0 1e-06 
0.0 1.3879 0 -2.0 1e-06 
0.0 1.388 0 -2.0 1e-06 
0.0 1.3881 0 -2.0 1e-06 
0.0 1.3882 0 -2.0 1e-06 
0.0 1.3883 0 -2.0 1e-06 
0.0 1.3884 0 -2.0 1e-06 
0.0 1.3885 0 -2.0 1e-06 
0.0 1.3886 0 -2.0 1e-06 
0.0 1.3887 0 -2.0 1e-06 
0.0 1.3888 0 -2.0 1e-06 
0.0 1.3889 0 -2.0 1e-06 
0.0 1.389 0 -2.0 1e-06 
0.0 1.3891 0 -2.0 1e-06 
0.0 1.3892 0 -2.0 1e-06 
0.0 1.3893 0 -2.0 1e-06 
0.0 1.3894 0 -2.0 1e-06 
0.0 1.3895 0 -2.0 1e-06 
0.0 1.3896 0 -2.0 1e-06 
0.0 1.3897 0 -2.0 1e-06 
0.0 1.3898 0 -2.0 1e-06 
0.0 1.3899 0 -2.0 1e-06 
0.0 1.39 0 -2.0 1e-06 
0.0 1.3901 0 -2.0 1e-06 
0.0 1.3902 0 -2.0 1e-06 
0.0 1.3903 0 -2.0 1e-06 
0.0 1.3904 0 -2.0 1e-06 
0.0 1.3905 0 -2.0 1e-06 
0.0 1.3906 0 -2.0 1e-06 
0.0 1.3907 0 -2.0 1e-06 
0.0 1.3908 0 -2.0 1e-06 
0.0 1.3909 0 -2.0 1e-06 
0.0 1.391 0 -2.0 1e-06 
0.0 1.3911 0 -2.0 1e-06 
0.0 1.3912 0 -2.0 1e-06 
0.0 1.3913 0 -2.0 1e-06 
0.0 1.3914 0 -2.0 1e-06 
0.0 1.3915 0 -2.0 1e-06 
0.0 1.3916 0 -2.0 1e-06 
0.0 1.3917 0 -2.0 1e-06 
0.0 1.3918 0 -2.0 1e-06 
0.0 1.3919 0 -2.0 1e-06 
0.0 1.392 0 -2.0 1e-06 
0.0 1.3921 0 -2.0 1e-06 
0.0 1.3922 0 -2.0 1e-06 
0.0 1.3923 0 -2.0 1e-06 
0.0 1.3924 0 -2.0 1e-06 
0.0 1.3925 0 -2.0 1e-06 
0.0 1.3926 0 -2.0 1e-06 
0.0 1.3927 0 -2.0 1e-06 
0.0 1.3928 0 -2.0 1e-06 
0.0 1.3929 0 -2.0 1e-06 
0.0 1.393 0 -2.0 1e-06 
0.0 1.3931 0 -2.0 1e-06 
0.0 1.3932 0 -2.0 1e-06 
0.0 1.3933 0 -2.0 1e-06 
0.0 1.3934 0 -2.0 1e-06 
0.0 1.3935 0 -2.0 1e-06 
0.0 1.3936 0 -2.0 1e-06 
0.0 1.3937 0 -2.0 1e-06 
0.0 1.3938 0 -2.0 1e-06 
0.0 1.3939 0 -2.0 1e-06 
0.0 1.394 0 -2.0 1e-06 
0.0 1.3941 0 -2.0 1e-06 
0.0 1.3942 0 -2.0 1e-06 
0.0 1.3943 0 -2.0 1e-06 
0.0 1.3944 0 -2.0 1e-06 
0.0 1.3945 0 -2.0 1e-06 
0.0 1.3946 0 -2.0 1e-06 
0.0 1.3947 0 -2.0 1e-06 
0.0 1.3948 0 -2.0 1e-06 
0.0 1.3949 0 -2.0 1e-06 
0.0 1.395 0 -2.0 1e-06 
0.0 1.3951 0 -2.0 1e-06 
0.0 1.3952 0 -2.0 1e-06 
0.0 1.3953 0 -2.0 1e-06 
0.0 1.3954 0 -2.0 1e-06 
0.0 1.3955 0 -2.0 1e-06 
0.0 1.3956 0 -2.0 1e-06 
0.0 1.3957 0 -2.0 1e-06 
0.0 1.3958 0 -2.0 1e-06 
0.0 1.3959 0 -2.0 1e-06 
0.0 1.396 0 -2.0 1e-06 
0.0 1.3961 0 -2.0 1e-06 
0.0 1.3962 0 -2.0 1e-06 
0.0 1.3963 0 -2.0 1e-06 
0.0 1.3964 0 -2.0 1e-06 
0.0 1.3965 0 -2.0 1e-06 
0.0 1.3966 0 -2.0 1e-06 
0.0 1.3967 0 -2.0 1e-06 
0.0 1.3968 0 -2.0 1e-06 
0.0 1.3969 0 -2.0 1e-06 
0.0 1.397 0 -2.0 1e-06 
0.0 1.3971 0 -2.0 1e-06 
0.0 1.3972 0 -2.0 1e-06 
0.0 1.3973 0 -2.0 1e-06 
0.0 1.3974 0 -2.0 1e-06 
0.0 1.3975 0 -2.0 1e-06 
0.0 1.3976 0 -2.0 1e-06 
0.0 1.3977 0 -2.0 1e-06 
0.0 1.3978 0 -2.0 1e-06 
0.0 1.3979 0 -2.0 1e-06 
0.0 1.398 0 -2.0 1e-06 
0.0 1.3981 0 -2.0 1e-06 
0.0 1.3982 0 -2.0 1e-06 
0.0 1.3983 0 -2.0 1e-06 
0.0 1.3984 0 -2.0 1e-06 
0.0 1.3985 0 -2.0 1e-06 
0.0 1.3986 0 -2.0 1e-06 
0.0 1.3987 0 -2.0 1e-06 
0.0 1.3988 0 -2.0 1e-06 
0.0 1.3989 0 -2.0 1e-06 
0.0 1.399 0 -2.0 1e-06 
0.0 1.3991 0 -2.0 1e-06 
0.0 1.3992 0 -2.0 1e-06 
0.0 1.3993 0 -2.0 1e-06 
0.0 1.3994 0 -2.0 1e-06 
0.0 1.3995 0 -2.0 1e-06 
0.0 1.3996 0 -2.0 1e-06 
0.0 1.3997 0 -2.0 1e-06 
0.0 1.3998 0 -2.0 1e-06 
0.0 1.3999 0 -2.0 1e-06 
0.0 1.4 0 -2.0 1e-06 
0.0 1.4001 0 -2.0 1e-06 
0.0 1.4002 0 -2.0 1e-06 
0.0 1.4003 0 -2.0 1e-06 
0.0 1.4004 0 -2.0 1e-06 
0.0 1.4005 0 -2.0 1e-06 
0.0 1.4006 0 -2.0 1e-06 
0.0 1.4007 0 -2.0 1e-06 
0.0 1.4008 0 -2.0 1e-06 
0.0 1.4009 0 -2.0 1e-06 
0.0 1.401 0 -2.0 1e-06 
0.0 1.4011 0 -2.0 1e-06 
0.0 1.4012 0 -2.0 1e-06 
0.0 1.4013 0 -2.0 1e-06 
0.0 1.4014 0 -2.0 1e-06 
0.0 1.4015 0 -2.0 1e-06 
0.0 1.4016 0 -2.0 1e-06 
0.0 1.4017 0 -2.0 1e-06 
0.0 1.4018 0 -2.0 1e-06 
0.0 1.4019 0 -2.0 1e-06 
0.0 1.402 0 -2.0 1e-06 
0.0 1.4021 0 -2.0 1e-06 
0.0 1.4022 0 -2.0 1e-06 
0.0 1.4023 0 -2.0 1e-06 
0.0 1.4024 0 -2.0 1e-06 
0.0 1.4025 0 -2.0 1e-06 
0.0 1.4026 0 -2.0 1e-06 
0.0 1.4027 0 -2.0 1e-06 
0.0 1.4028 0 -2.0 1e-06 
0.0 1.4029 0 -2.0 1e-06 
0.0 1.403 0 -2.0 1e-06 
0.0 1.4031 0 -2.0 1e-06 
0.0 1.4032 0 -2.0 1e-06 
0.0 1.4033 0 -2.0 1e-06 
0.0 1.4034 0 -2.0 1e-06 
0.0 1.4035 0 -2.0 1e-06 
0.0 1.4036 0 -2.0 1e-06 
0.0 1.4037 0 -2.0 1e-06 
0.0 1.4038 0 -2.0 1e-06 
0.0 1.4039 0 -2.0 1e-06 
0.0 1.404 0 -2.0 1e-06 
0.0 1.4041 0 -2.0 1e-06 
0.0 1.4042 0 -2.0 1e-06 
0.0 1.4043 0 -2.0 1e-06 
0.0 1.4044 0 -2.0 1e-06 
0.0 1.4045 0 -2.0 1e-06 
0.0 1.4046 0 -2.0 1e-06 
0.0 1.4047 0 -2.0 1e-06 
0.0 1.4048 0 -2.0 1e-06 
0.0 1.4049 0 -2.0 1e-06 
0.0 1.405 0 -2.0 1e-06 
0.0 1.4051 0 -2.0 1e-06 
0.0 1.4052 0 -2.0 1e-06 
0.0 1.4053 0 -2.0 1e-06 
0.0 1.4054 0 -2.0 1e-06 
0.0 1.4055 0 -2.0 1e-06 
0.0 1.4056 0 -2.0 1e-06 
0.0 1.4057 0 -2.0 1e-06 
0.0 1.4058 0 -2.0 1e-06 
0.0 1.4059 0 -2.0 1e-06 
0.0 1.406 0 -2.0 1e-06 
0.0 1.4061 0 -2.0 1e-06 
0.0 1.4062 0 -2.0 1e-06 
0.0 1.4063 0 -2.0 1e-06 
0.0 1.4064 0 -2.0 1e-06 
0.0 1.4065 0 -2.0 1e-06 
0.0 1.4066 0 -2.0 1e-06 
0.0 1.4067 0 -2.0 1e-06 
0.0 1.4068 0 -2.0 1e-06 
0.0 1.4069 0 -2.0 1e-06 
0.0 1.407 0 -2.0 1e-06 
0.0 1.4071 0 -2.0 1e-06 
0.0 1.4072 0 -2.0 1e-06 
0.0 1.4073 0 -2.0 1e-06 
0.0 1.4074 0 -2.0 1e-06 
0.0 1.4075 0 -2.0 1e-06 
0.0 1.4076 0 -2.0 1e-06 
0.0 1.4077 0 -2.0 1e-06 
0.0 1.4078 0 -2.0 1e-06 
0.0 1.4079 0 -2.0 1e-06 
0.0 1.408 0 -2.0 1e-06 
0.0 1.4081 0 -2.0 1e-06 
0.0 1.4082 0 -2.0 1e-06 
0.0 1.4083 0 -2.0 1e-06 
0.0 1.4084 0 -2.0 1e-06 
0.0 1.4085 0 -2.0 1e-06 
0.0 1.4086 0 -2.0 1e-06 
0.0 1.4087 0 -2.0 1e-06 
0.0 1.4088 0 -2.0 1e-06 
0.0 1.4089 0 -2.0 1e-06 
0.0 1.409 0 -2.0 1e-06 
0.0 1.4091 0 -2.0 1e-06 
0.0 1.4092 0 -2.0 1e-06 
0.0 1.4093 0 -2.0 1e-06 
0.0 1.4094 0 -2.0 1e-06 
0.0 1.4095 0 -2.0 1e-06 
0.0 1.4096 0 -2.0 1e-06 
0.0 1.4097 0 -2.0 1e-06 
0.0 1.4098 0 -2.0 1e-06 
0.0 1.4099 0 -2.0 1e-06 
0.0 1.41 0 -2.0 1e-06 
0.0 1.4101 0 -2.0 1e-06 
0.0 1.4102 0 -2.0 1e-06 
0.0 1.4103 0 -2.0 1e-06 
0.0 1.4104 0 -2.0 1e-06 
0.0 1.4105 0 -2.0 1e-06 
0.0 1.4106 0 -2.0 1e-06 
0.0 1.4107 0 -2.0 1e-06 
0.0 1.4108 0 -2.0 1e-06 
0.0 1.4109 0 -2.0 1e-06 
0.0 1.411 0 -2.0 1e-06 
0.0 1.4111 0 -2.0 1e-06 
0.0 1.4112 0 -2.0 1e-06 
0.0 1.4113 0 -2.0 1e-06 
0.0 1.4114 0 -2.0 1e-06 
0.0 1.4115 0 -2.0 1e-06 
0.0 1.4116 0 -2.0 1e-06 
0.0 1.4117 0 -2.0 1e-06 
0.0 1.4118 0 -2.0 1e-06 
0.0 1.4119 0 -2.0 1e-06 
0.0 1.412 0 -2.0 1e-06 
0.0 1.4121 0 -2.0 1e-06 
0.0 1.4122 0 -2.0 1e-06 
0.0 1.4123 0 -2.0 1e-06 
0.0 1.4124 0 -2.0 1e-06 
0.0 1.4125 0 -2.0 1e-06 
0.0 1.4126 0 -2.0 1e-06 
0.0 1.4127 0 -2.0 1e-06 
0.0 1.4128 0 -2.0 1e-06 
0.0 1.4129 0 -2.0 1e-06 
0.0 1.413 0 -2.0 1e-06 
0.0 1.4131 0 -2.0 1e-06 
0.0 1.4132 0 -2.0 1e-06 
0.0 1.4133 0 -2.0 1e-06 
0.0 1.4134 0 -2.0 1e-06 
0.0 1.4135 0 -2.0 1e-06 
0.0 1.4136 0 -2.0 1e-06 
0.0 1.4137 0 -2.0 1e-06 
0.0 1.4138 0 -2.0 1e-06 
0.0 1.4139 0 -2.0 1e-06 
0.0 1.414 0 -2.0 1e-06 
0.0 1.4141 0 -2.0 1e-06 
0.0 1.4142 0 -2.0 1e-06 
0.0 1.4143 0 -2.0 1e-06 
0.0 1.4144 0 -2.0 1e-06 
0.0 1.4145 0 -2.0 1e-06 
0.0 1.4146 0 -2.0 1e-06 
0.0 1.4147 0 -2.0 1e-06 
0.0 1.4148 0 -2.0 1e-06 
0.0 1.4149 0 -2.0 1e-06 
0.0 1.415 0 -2.0 1e-06 
0.0 1.4151 0 -2.0 1e-06 
0.0 1.4152 0 -2.0 1e-06 
0.0 1.4153 0 -2.0 1e-06 
0.0 1.4154 0 -2.0 1e-06 
0.0 1.4155 0 -2.0 1e-06 
0.0 1.4156 0 -2.0 1e-06 
0.0 1.4157 0 -2.0 1e-06 
0.0 1.4158 0 -2.0 1e-06 
0.0 1.4159 0 -2.0 1e-06 
0.0 1.416 0 -2.0 1e-06 
0.0 1.4161 0 -2.0 1e-06 
0.0 1.4162 0 -2.0 1e-06 
0.0 1.4163 0 -2.0 1e-06 
0.0 1.4164 0 -2.0 1e-06 
0.0 1.4165 0 -2.0 1e-06 
0.0 1.4166 0 -2.0 1e-06 
0.0 1.4167 0 -2.0 1e-06 
0.0 1.4168 0 -2.0 1e-06 
0.0 1.4169 0 -2.0 1e-06 
0.0 1.417 0 -2.0 1e-06 
0.0 1.4171 0 -2.0 1e-06 
0.0 1.4172 0 -2.0 1e-06 
0.0 1.4173 0 -2.0 1e-06 
0.0 1.4174 0 -2.0 1e-06 
0.0 1.4175 0 -2.0 1e-06 
0.0 1.4176 0 -2.0 1e-06 
0.0 1.4177 0 -2.0 1e-06 
0.0 1.4178 0 -2.0 1e-06 
0.0 1.4179 0 -2.0 1e-06 
0.0 1.418 0 -2.0 1e-06 
0.0 1.4181 0 -2.0 1e-06 
0.0 1.4182 0 -2.0 1e-06 
0.0 1.4183 0 -2.0 1e-06 
0.0 1.4184 0 -2.0 1e-06 
0.0 1.4185 0 -2.0 1e-06 
0.0 1.4186 0 -2.0 1e-06 
0.0 1.4187 0 -2.0 1e-06 
0.0 1.4188 0 -2.0 1e-06 
0.0 1.4189 0 -2.0 1e-06 
0.0 1.419 0 -2.0 1e-06 
0.0 1.4191 0 -2.0 1e-06 
0.0 1.4192 0 -2.0 1e-06 
0.0 1.4193 0 -2.0 1e-06 
0.0 1.4194 0 -2.0 1e-06 
0.0 1.4195 0 -2.0 1e-06 
0.0 1.4196 0 -2.0 1e-06 
0.0 1.4197 0 -2.0 1e-06 
0.0 1.4198 0 -2.0 1e-06 
0.0 1.4199 0 -2.0 1e-06 
0.0 1.42 0 -2.0 1e-06 
0.0 1.4201 0 -2.0 1e-06 
0.0 1.4202 0 -2.0 1e-06 
0.0 1.4203 0 -2.0 1e-06 
0.0 1.4204 0 -2.0 1e-06 
0.0 1.4205 0 -2.0 1e-06 
0.0 1.4206 0 -2.0 1e-06 
0.0 1.4207 0 -2.0 1e-06 
0.0 1.4208 0 -2.0 1e-06 
0.0 1.4209 0 -2.0 1e-06 
0.0 1.421 0 -2.0 1e-06 
0.0 1.4211 0 -2.0 1e-06 
0.0 1.4212 0 -2.0 1e-06 
0.0 1.4213 0 -2.0 1e-06 
0.0 1.4214 0 -2.0 1e-06 
0.0 1.4215 0 -2.0 1e-06 
0.0 1.4216 0 -2.0 1e-06 
0.0 1.4217 0 -2.0 1e-06 
0.0 1.4218 0 -2.0 1e-06 
0.0 1.4219 0 -2.0 1e-06 
0.0 1.422 0 -2.0 1e-06 
0.0 1.4221 0 -2.0 1e-06 
0.0 1.4222 0 -2.0 1e-06 
0.0 1.4223 0 -2.0 1e-06 
0.0 1.4224 0 -2.0 1e-06 
0.0 1.4225 0 -2.0 1e-06 
0.0 1.4226 0 -2.0 1e-06 
0.0 1.4227 0 -2.0 1e-06 
0.0 1.4228 0 -2.0 1e-06 
0.0 1.4229 0 -2.0 1e-06 
0.0 1.423 0 -2.0 1e-06 
0.0 1.4231 0 -2.0 1e-06 
0.0 1.4232 0 -2.0 1e-06 
0.0 1.4233 0 -2.0 1e-06 
0.0 1.4234 0 -2.0 1e-06 
0.0 1.4235 0 -2.0 1e-06 
0.0 1.4236 0 -2.0 1e-06 
0.0 1.4237 0 -2.0 1e-06 
0.0 1.4238 0 -2.0 1e-06 
0.0 1.4239 0 -2.0 1e-06 
0.0 1.424 0 -2.0 1e-06 
0.0 1.4241 0 -2.0 1e-06 
0.0 1.4242 0 -2.0 1e-06 
0.0 1.4243 0 -2.0 1e-06 
0.0 1.4244 0 -2.0 1e-06 
0.0 1.4245 0 -2.0 1e-06 
0.0 1.4246 0 -2.0 1e-06 
0.0 1.4247 0 -2.0 1e-06 
0.0 1.4248 0 -2.0 1e-06 
0.0 1.4249 0 -2.0 1e-06 
0.0 1.425 0 -2.0 1e-06 
0.0 1.4251 0 -2.0 1e-06 
0.0 1.4252 0 -2.0 1e-06 
0.0 1.4253 0 -2.0 1e-06 
0.0 1.4254 0 -2.0 1e-06 
0.0 1.4255 0 -2.0 1e-06 
0.0 1.4256 0 -2.0 1e-06 
0.0 1.4257 0 -2.0 1e-06 
0.0 1.4258 0 -2.0 1e-06 
0.0 1.4259 0 -2.0 1e-06 
0.0 1.426 0 -2.0 1e-06 
0.0 1.4261 0 -2.0 1e-06 
0.0 1.4262 0 -2.0 1e-06 
0.0 1.4263 0 -2.0 1e-06 
0.0 1.4264 0 -2.0 1e-06 
0.0 1.4265 0 -2.0 1e-06 
0.0 1.4266 0 -2.0 1e-06 
0.0 1.4267 0 -2.0 1e-06 
0.0 1.4268 0 -2.0 1e-06 
0.0 1.4269 0 -2.0 1e-06 
0.0 1.427 0 -2.0 1e-06 
0.0 1.4271 0 -2.0 1e-06 
0.0 1.4272 0 -2.0 1e-06 
0.0 1.4273 0 -2.0 1e-06 
0.0 1.4274 0 -2.0 1e-06 
0.0 1.4275 0 -2.0 1e-06 
0.0 1.4276 0 -2.0 1e-06 
0.0 1.4277 0 -2.0 1e-06 
0.0 1.4278 0 -2.0 1e-06 
0.0 1.4279 0 -2.0 1e-06 
0.0 1.428 0 -2.0 1e-06 
0.0 1.4281 0 -2.0 1e-06 
0.0 1.4282 0 -2.0 1e-06 
0.0 1.4283 0 -2.0 1e-06 
0.0 1.4284 0 -2.0 1e-06 
0.0 1.4285 0 -2.0 1e-06 
0.0 1.4286 0 -2.0 1e-06 
0.0 1.4287 0 -2.0 1e-06 
0.0 1.4288 0 -2.0 1e-06 
0.0 1.4289 0 -2.0 1e-06 
0.0 1.429 0 -2.0 1e-06 
0.0 1.4291 0 -2.0 1e-06 
0.0 1.4292 0 -2.0 1e-06 
0.0 1.4293 0 -2.0 1e-06 
0.0 1.4294 0 -2.0 1e-06 
0.0 1.4295 0 -2.0 1e-06 
0.0 1.4296 0 -2.0 1e-06 
0.0 1.4297 0 -2.0 1e-06 
0.0 1.4298 0 -2.0 1e-06 
0.0 1.4299 0 -2.0 1e-06 
0.0 1.43 0 -2.0 1e-06 
0.0 1.4301 0 -2.0 1e-06 
0.0 1.4302 0 -2.0 1e-06 
0.0 1.4303 0 -2.0 1e-06 
0.0 1.4304 0 -2.0 1e-06 
0.0 1.4305 0 -2.0 1e-06 
0.0 1.4306 0 -2.0 1e-06 
0.0 1.4307 0 -2.0 1e-06 
0.0 1.4308 0 -2.0 1e-06 
0.0 1.4309 0 -2.0 1e-06 
0.0 1.431 0 -2.0 1e-06 
0.0 1.4311 0 -2.0 1e-06 
0.0 1.4312 0 -2.0 1e-06 
0.0 1.4313 0 -2.0 1e-06 
0.0 1.4314 0 -2.0 1e-06 
0.0 1.4315 0 -2.0 1e-06 
0.0 1.4316 0 -2.0 1e-06 
0.0 1.4317 0 -2.0 1e-06 
0.0 1.4318 0 -2.0 1e-06 
0.0 1.4319 0 -2.0 1e-06 
0.0 1.432 0 -2.0 1e-06 
0.0 1.4321 0 -2.0 1e-06 
0.0 1.4322 0 -2.0 1e-06 
0.0 1.4323 0 -2.0 1e-06 
0.0 1.4324 0 -2.0 1e-06 
0.0 1.4325 0 -2.0 1e-06 
0.0 1.4326 0 -2.0 1e-06 
0.0 1.4327 0 -2.0 1e-06 
0.0 1.4328 0 -2.0 1e-06 
0.0 1.4329 0 -2.0 1e-06 
0.0 1.433 0 -2.0 1e-06 
0.0 1.4331 0 -2.0 1e-06 
0.0 1.4332 0 -2.0 1e-06 
0.0 1.4333 0 -2.0 1e-06 
0.0 1.4334 0 -2.0 1e-06 
0.0 1.4335 0 -2.0 1e-06 
0.0 1.4336 0 -2.0 1e-06 
0.0 1.4337 0 -2.0 1e-06 
0.0 1.4338 0 -2.0 1e-06 
0.0 1.4339 0 -2.0 1e-06 
0.0 1.434 0 -2.0 1e-06 
0.0 1.4341 0 -2.0 1e-06 
0.0 1.4342 0 -2.0 1e-06 
0.0 1.4343 0 -2.0 1e-06 
0.0 1.4344 0 -2.0 1e-06 
0.0 1.4345 0 -2.0 1e-06 
0.0 1.4346 0 -2.0 1e-06 
0.0 1.4347 0 -2.0 1e-06 
0.0 1.4348 0 -2.0 1e-06 
0.0 1.4349 0 -2.0 1e-06 
0.0 1.435 0 -2.0 1e-06 
0.0 1.4351 0 -2.0 1e-06 
0.0 1.4352 0 -2.0 1e-06 
0.0 1.4353 0 -2.0 1e-06 
0.0 1.4354 0 -2.0 1e-06 
0.0 1.4355 0 -2.0 1e-06 
0.0 1.4356 0 -2.0 1e-06 
0.0 1.4357 0 -2.0 1e-06 
0.0 1.4358 0 -2.0 1e-06 
0.0 1.4359 0 -2.0 1e-06 
0.0 1.436 0 -2.0 1e-06 
0.0 1.4361 0 -2.0 1e-06 
0.0 1.4362 0 -2.0 1e-06 
0.0 1.4363 0 -2.0 1e-06 
0.0 1.4364 0 -2.0 1e-06 
0.0 1.4365 0 -2.0 1e-06 
0.0 1.4366 0 -2.0 1e-06 
0.0 1.4367 0 -2.0 1e-06 
0.0 1.4368 0 -2.0 1e-06 
0.0 1.4369 0 -2.0 1e-06 
0.0 1.437 0 -2.0 1e-06 
0.0 1.4371 0 -2.0 1e-06 
0.0 1.4372 0 -2.0 1e-06 
0.0 1.4373 0 -2.0 1e-06 
0.0 1.4374 0 -2.0 1e-06 
0.0 1.4375 0 -2.0 1e-06 
0.0 1.4376 0 -2.0 1e-06 
0.0 1.4377 0 -2.0 1e-06 
0.0 1.4378 0 -2.0 1e-06 
0.0 1.4379 0 -2.0 1e-06 
0.0 1.438 0 -2.0 1e-06 
0.0 1.4381 0 -2.0 1e-06 
0.0 1.4382 0 -2.0 1e-06 
0.0 1.4383 0 -2.0 1e-06 
0.0 1.4384 0 -2.0 1e-06 
0.0 1.4385 0 -2.0 1e-06 
0.0 1.4386 0 -2.0 1e-06 
0.0 1.4387 0 -2.0 1e-06 
0.0 1.4388 0 -2.0 1e-06 
0.0 1.4389 0 -2.0 1e-06 
0.0 1.439 0 -2.0 1e-06 
0.0 1.4391 0 -2.0 1e-06 
0.0 1.4392 0 -2.0 1e-06 
0.0 1.4393 0 -2.0 1e-06 
0.0 1.4394 0 -2.0 1e-06 
0.0 1.4395 0 -2.0 1e-06 
0.0 1.4396 0 -2.0 1e-06 
0.0 1.4397 0 -2.0 1e-06 
0.0 1.4398 0 -2.0 1e-06 
0.0 1.4399 0 -2.0 1e-06 
0.0 1.44 0 -2.0 1e-06 
0.0 1.4401 0 -2.0 1e-06 
0.0 1.4402 0 -2.0 1e-06 
0.0 1.4403 0 -2.0 1e-06 
0.0 1.4404 0 -2.0 1e-06 
0.0 1.4405 0 -2.0 1e-06 
0.0 1.4406 0 -2.0 1e-06 
0.0 1.4407 0 -2.0 1e-06 
0.0 1.4408 0 -2.0 1e-06 
0.0 1.4409 0 -2.0 1e-06 
0.0 1.441 0 -2.0 1e-06 
0.0 1.4411 0 -2.0 1e-06 
0.0 1.4412 0 -2.0 1e-06 
0.0 1.4413 0 -2.0 1e-06 
0.0 1.4414 0 -2.0 1e-06 
0.0 1.4415 0 -2.0 1e-06 
0.0 1.4416 0 -2.0 1e-06 
0.0 1.4417 0 -2.0 1e-06 
0.0 1.4418 0 -2.0 1e-06 
0.0 1.4419 0 -2.0 1e-06 
0.0 1.442 0 -2.0 1e-06 
0.0 1.4421 0 -2.0 1e-06 
0.0 1.4422 0 -2.0 1e-06 
0.0 1.4423 0 -2.0 1e-06 
0.0 1.4424 0 -2.0 1e-06 
0.0 1.4425 0 -2.0 1e-06 
0.0 1.4426 0 -2.0 1e-06 
0.0 1.4427 0 -2.0 1e-06 
0.0 1.4428 0 -2.0 1e-06 
0.0 1.4429 0 -2.0 1e-06 
0.0 1.443 0 -2.0 1e-06 
0.0 1.4431 0 -2.0 1e-06 
0.0 1.4432 0 -2.0 1e-06 
0.0 1.4433 0 -2.0 1e-06 
0.0 1.4434 0 -2.0 1e-06 
0.0 1.4435 0 -2.0 1e-06 
0.0 1.4436 0 -2.0 1e-06 
0.0 1.4437 0 -2.0 1e-06 
0.0 1.4438 0 -2.0 1e-06 
0.0 1.4439 0 -2.0 1e-06 
0.0 1.444 0 -2.0 1e-06 
0.0 1.4441 0 -2.0 1e-06 
0.0 1.4442 0 -2.0 1e-06 
0.0 1.4443 0 -2.0 1e-06 
0.0 1.4444 0 -2.0 1e-06 
0.0 1.4445 0 -2.0 1e-06 
0.0 1.4446 0 -2.0 1e-06 
0.0 1.4447 0 -2.0 1e-06 
0.0 1.4448 0 -2.0 1e-06 
0.0 1.4449 0 -2.0 1e-06 
0.0 1.445 0 -2.0 1e-06 
0.0 1.4451 0 -2.0 1e-06 
0.0 1.4452 0 -2.0 1e-06 
0.0 1.4453 0 -2.0 1e-06 
0.0 1.4454 0 -2.0 1e-06 
0.0 1.4455 0 -2.0 1e-06 
0.0 1.4456 0 -2.0 1e-06 
0.0 1.4457 0 -2.0 1e-06 
0.0 1.4458 0 -2.0 1e-06 
0.0 1.4459 0 -2.0 1e-06 
0.0 1.446 0 -2.0 1e-06 
0.0 1.4461 0 -2.0 1e-06 
0.0 1.4462 0 -2.0 1e-06 
0.0 1.4463 0 -2.0 1e-06 
0.0 1.4464 0 -2.0 1e-06 
0.0 1.4465 0 -2.0 1e-06 
0.0 1.4466 0 -2.0 1e-06 
0.0 1.4467 0 -2.0 1e-06 
0.0 1.4468 0 -2.0 1e-06 
0.0 1.4469 0 -2.0 1e-06 
0.0 1.447 0 -2.0 1e-06 
0.0 1.4471 0 -2.0 1e-06 
0.0 1.4472 0 -2.0 1e-06 
0.0 1.4473 0 -2.0 1e-06 
0.0 1.4474 0 -2.0 1e-06 
0.0 1.4475 0 -2.0 1e-06 
0.0 1.4476 0 -2.0 1e-06 
0.0 1.4477 0 -2.0 1e-06 
0.0 1.4478 0 -2.0 1e-06 
0.0 1.4479 0 -2.0 1e-06 
0.0 1.448 0 -2.0 1e-06 
0.0 1.4481 0 -2.0 1e-06 
0.0 1.4482 0 -2.0 1e-06 
0.0 1.4483 0 -2.0 1e-06 
0.0 1.4484 0 -2.0 1e-06 
0.0 1.4485 0 -2.0 1e-06 
0.0 1.4486 0 -2.0 1e-06 
0.0 1.4487 0 -2.0 1e-06 
0.0 1.4488 0 -2.0 1e-06 
0.0 1.4489 0 -2.0 1e-06 
0.0 1.449 0 -2.0 1e-06 
0.0 1.4491 0 -2.0 1e-06 
0.0 1.4492 0 -2.0 1e-06 
0.0 1.4493 0 -2.0 1e-06 
0.0 1.4494 0 -2.0 1e-06 
0.0 1.4495 0 -2.0 1e-06 
0.0 1.4496 0 -2.0 1e-06 
0.0 1.4497 0 -2.0 1e-06 
0.0 1.4498 0 -2.0 1e-06 
0.0 1.4499 0 -2.0 1e-06 
0.0 1.45 0 -2.0 1e-06 
0.0 1.4501 0 -2.0 1e-06 
0.0 1.4502 0 -2.0 1e-06 
0.0 1.4503 0 -2.0 1e-06 
0.0 1.4504 0 -2.0 1e-06 
0.0 1.4505 0 -2.0 1e-06 
0.0 1.4506 0 -2.0 1e-06 
0.0 1.4507 0 -2.0 1e-06 
0.0 1.4508 0 -2.0 1e-06 
0.0 1.4509 0 -2.0 1e-06 
0.0 1.451 0 -2.0 1e-06 
0.0 1.4511 0 -2.0 1e-06 
0.0 1.4512 0 -2.0 1e-06 
0.0 1.4513 0 -2.0 1e-06 
0.0 1.4514 0 -2.0 1e-06 
0.0 1.4515 0 -2.0 1e-06 
0.0 1.4516 0 -2.0 1e-06 
0.0 1.4517 0 -2.0 1e-06 
0.0 1.4518 0 -2.0 1e-06 
0.0 1.4519 0 -2.0 1e-06 
0.0 1.452 0 -2.0 1e-06 
0.0 1.4521 0 -2.0 1e-06 
0.0 1.4522 0 -2.0 1e-06 
0.0 1.4523 0 -2.0 1e-06 
0.0 1.4524 0 -2.0 1e-06 
0.0 1.4525 0 -2.0 1e-06 
0.0 1.4526 0 -2.0 1e-06 
0.0 1.4527 0 -2.0 1e-06 
0.0 1.4528 0 -2.0 1e-06 
0.0 1.4529 0 -2.0 1e-06 
0.0 1.453 0 -2.0 1e-06 
0.0 1.4531 0 -2.0 1e-06 
0.0 1.4532 0 -2.0 1e-06 
0.0 1.4533 0 -2.0 1e-06 
0.0 1.4534 0 -2.0 1e-06 
0.0 1.4535 0 -2.0 1e-06 
0.0 1.4536 0 -2.0 1e-06 
0.0 1.4537 0 -2.0 1e-06 
0.0 1.4538 0 -2.0 1e-06 
0.0 1.4539 0 -2.0 1e-06 
0.0 1.454 0 -2.0 1e-06 
0.0 1.4541 0 -2.0 1e-06 
0.0 1.4542 0 -2.0 1e-06 
0.0 1.4543 0 -2.0 1e-06 
0.0 1.4544 0 -2.0 1e-06 
0.0 1.4545 0 -2.0 1e-06 
0.0 1.4546 0 -2.0 1e-06 
0.0 1.4547 0 -2.0 1e-06 
0.0 1.4548 0 -2.0 1e-06 
0.0 1.4549 0 -2.0 1e-06 
0.0 1.455 0 -2.0 1e-06 
0.0 1.4551 0 -2.0 1e-06 
0.0 1.4552 0 -2.0 1e-06 
0.0 1.4553 0 -2.0 1e-06 
0.0 1.4554 0 -2.0 1e-06 
0.0 1.4555 0 -2.0 1e-06 
0.0 1.4556 0 -2.0 1e-06 
0.0 1.4557 0 -2.0 1e-06 
0.0 1.4558 0 -2.0 1e-06 
0.0 1.4559 0 -2.0 1e-06 
0.0 1.456 0 -2.0 1e-06 
0.0 1.4561 0 -2.0 1e-06 
0.0 1.4562 0 -2.0 1e-06 
0.0 1.4563 0 -2.0 1e-06 
0.0 1.4564 0 -2.0 1e-06 
0.0 1.4565 0 -2.0 1e-06 
0.0 1.4566 0 -2.0 1e-06 
0.0 1.4567 0 -2.0 1e-06 
0.0 1.4568 0 -2.0 1e-06 
0.0 1.4569 0 -2.0 1e-06 
0.0 1.457 0 -2.0 1e-06 
0.0 1.4571 0 -2.0 1e-06 
0.0 1.4572 0 -2.0 1e-06 
0.0 1.4573 0 -2.0 1e-06 
0.0 1.4574 0 -2.0 1e-06 
0.0 1.4575 0 -2.0 1e-06 
0.0 1.4576 0 -2.0 1e-06 
0.0 1.4577 0 -2.0 1e-06 
0.0 1.4578 0 -2.0 1e-06 
0.0 1.4579 0 -2.0 1e-06 
0.0 1.458 0 -2.0 1e-06 
0.0 1.4581 0 -2.0 1e-06 
0.0 1.4582 0 -2.0 1e-06 
0.0 1.4583 0 -2.0 1e-06 
0.0 1.4584 0 -2.0 1e-06 
0.0 1.4585 0 -2.0 1e-06 
0.0 1.4586 0 -2.0 1e-06 
0.0 1.4587 0 -2.0 1e-06 
0.0 1.4588 0 -2.0 1e-06 
0.0 1.4589 0 -2.0 1e-06 
0.0 1.459 0 -2.0 1e-06 
0.0 1.4591 0 -2.0 1e-06 
0.0 1.4592 0 -2.0 1e-06 
0.0 1.4593 0 -2.0 1e-06 
0.0 1.4594 0 -2.0 1e-06 
0.0 1.4595 0 -2.0 1e-06 
0.0 1.4596 0 -2.0 1e-06 
0.0 1.4597 0 -2.0 1e-06 
0.0 1.4598 0 -2.0 1e-06 
0.0 1.4599 0 -2.0 1e-06 
0.0 1.46 0 -2.0 1e-06 
0.0 1.4601 0 -2.0 1e-06 
0.0 1.4602 0 -2.0 1e-06 
0.0 1.4603 0 -2.0 1e-06 
0.0 1.4604 0 -2.0 1e-06 
0.0 1.4605 0 -2.0 1e-06 
0.0 1.4606 0 -2.0 1e-06 
0.0 1.4607 0 -2.0 1e-06 
0.0 1.4608 0 -2.0 1e-06 
0.0 1.4609 0 -2.0 1e-06 
0.0 1.461 0 -2.0 1e-06 
0.0 1.4611 0 -2.0 1e-06 
0.0 1.4612 0 -2.0 1e-06 
0.0 1.4613 0 -2.0 1e-06 
0.0 1.4614 0 -2.0 1e-06 
0.0 1.4615 0 -2.0 1e-06 
0.0 1.4616 0 -2.0 1e-06 
0.0 1.4617 0 -2.0 1e-06 
0.0 1.4618 0 -2.0 1e-06 
0.0 1.4619 0 -2.0 1e-06 
0.0 1.462 0 -2.0 1e-06 
0.0 1.4621 0 -2.0 1e-06 
0.0 1.4622 0 -2.0 1e-06 
0.0 1.4623 0 -2.0 1e-06 
0.0 1.4624 0 -2.0 1e-06 
0.0 1.4625 0 -2.0 1e-06 
0.0 1.4626 0 -2.0 1e-06 
0.0 1.4627 0 -2.0 1e-06 
0.0 1.4628 0 -2.0 1e-06 
0.0 1.4629 0 -2.0 1e-06 
0.0 1.463 0 -2.0 1e-06 
0.0 1.4631 0 -2.0 1e-06 
0.0 1.4632 0 -2.0 1e-06 
0.0 1.4633 0 -2.0 1e-06 
0.0 1.4634 0 -2.0 1e-06 
0.0 1.4635 0 -2.0 1e-06 
0.0 1.4636 0 -2.0 1e-06 
0.0 1.4637 0 -2.0 1e-06 
0.0 1.4638 0 -2.0 1e-06 
0.0 1.4639 0 -2.0 1e-06 
0.0 1.464 0 -2.0 1e-06 
0.0 1.4641 0 -2.0 1e-06 
0.0 1.4642 0 -2.0 1e-06 
0.0 1.4643 0 -2.0 1e-06 
0.0 1.4644 0 -2.0 1e-06 
0.0 1.4645 0 -2.0 1e-06 
0.0 1.4646 0 -2.0 1e-06 
0.0 1.4647 0 -2.0 1e-06 
0.0 1.4648 0 -2.0 1e-06 
0.0 1.4649 0 -2.0 1e-06 
0.0 1.465 0 -2.0 1e-06 
0.0 1.4651 0 -2.0 1e-06 
0.0 1.4652 0 -2.0 1e-06 
0.0 1.4653 0 -2.0 1e-06 
0.0 1.4654 0 -2.0 1e-06 
0.0 1.4655 0 -2.0 1e-06 
0.0 1.4656 0 -2.0 1e-06 
0.0 1.4657 0 -2.0 1e-06 
0.0 1.4658 0 -2.0 1e-06 
0.0 1.4659 0 -2.0 1e-06 
0.0 1.466 0 -2.0 1e-06 
0.0 1.4661 0 -2.0 1e-06 
0.0 1.4662 0 -2.0 1e-06 
0.0 1.4663 0 -2.0 1e-06 
0.0 1.4664 0 -2.0 1e-06 
0.0 1.4665 0 -2.0 1e-06 
0.0 1.4666 0 -2.0 1e-06 
0.0 1.4667 0 -2.0 1e-06 
0.0 1.4668 0 -2.0 1e-06 
0.0 1.4669 0 -2.0 1e-06 
0.0 1.467 0 -2.0 1e-06 
0.0 1.4671 0 -2.0 1e-06 
0.0 1.4672 0 -2.0 1e-06 
0.0 1.4673 0 -2.0 1e-06 
0.0 1.4674 0 -2.0 1e-06 
0.0 1.4675 0 -2.0 1e-06 
0.0 1.4676 0 -2.0 1e-06 
0.0 1.4677 0 -2.0 1e-06 
0.0 1.4678 0 -2.0 1e-06 
0.0 1.4679 0 -2.0 1e-06 
0.0 1.468 0 -2.0 1e-06 
0.0 1.4681 0 -2.0 1e-06 
0.0 1.4682 0 -2.0 1e-06 
0.0 1.4683 0 -2.0 1e-06 
0.0 1.4684 0 -2.0 1e-06 
0.0 1.4685 0 -2.0 1e-06 
0.0 1.4686 0 -2.0 1e-06 
0.0 1.4687 0 -2.0 1e-06 
0.0 1.4688 0 -2.0 1e-06 
0.0 1.4689 0 -2.0 1e-06 
0.0 1.469 0 -2.0 1e-06 
0.0 1.4691 0 -2.0 1e-06 
0.0 1.4692 0 -2.0 1e-06 
0.0 1.4693 0 -2.0 1e-06 
0.0 1.4694 0 -2.0 1e-06 
0.0 1.4695 0 -2.0 1e-06 
0.0 1.4696 0 -2.0 1e-06 
0.0 1.4697 0 -2.0 1e-06 
0.0 1.4698 0 -2.0 1e-06 
0.0 1.4699 0 -2.0 1e-06 
0.0 1.47 0 -2.0 1e-06 
0.0 1.4701 0 -2.0 1e-06 
0.0 1.4702 0 -2.0 1e-06 
0.0 1.4703 0 -2.0 1e-06 
0.0 1.4704 0 -2.0 1e-06 
0.0 1.4705 0 -2.0 1e-06 
0.0 1.4706 0 -2.0 1e-06 
0.0 1.4707 0 -2.0 1e-06 
0.0 1.4708 0 -2.0 1e-06 
0.0 1.4709 0 -2.0 1e-06 
0.0 1.471 0 -2.0 1e-06 
0.0 1.4711 0 -2.0 1e-06 
0.0 1.4712 0 -2.0 1e-06 
0.0 1.4713 0 -2.0 1e-06 
0.0 1.4714 0 -2.0 1e-06 
0.0 1.4715 0 -2.0 1e-06 
0.0 1.4716 0 -2.0 1e-06 
0.0 1.4717 0 -2.0 1e-06 
0.0 1.4718 0 -2.0 1e-06 
0.0 1.4719 0 -2.0 1e-06 
0.0 1.472 0 -2.0 1e-06 
0.0 1.4721 0 -2.0 1e-06 
0.0 1.4722 0 -2.0 1e-06 
0.0 1.4723 0 -2.0 1e-06 
0.0 1.4724 0 -2.0 1e-06 
0.0 1.4725 0 -2.0 1e-06 
0.0 1.4726 0 -2.0 1e-06 
0.0 1.4727 0 -2.0 1e-06 
0.0 1.4728 0 -2.0 1e-06 
0.0 1.4729 0 -2.0 1e-06 
0.0 1.473 0 -2.0 1e-06 
0.0 1.4731 0 -2.0 1e-06 
0.0 1.4732 0 -2.0 1e-06 
0.0 1.4733 0 -2.0 1e-06 
0.0 1.4734 0 -2.0 1e-06 
0.0 1.4735 0 -2.0 1e-06 
0.0 1.4736 0 -2.0 1e-06 
0.0 1.4737 0 -2.0 1e-06 
0.0 1.4738 0 -2.0 1e-06 
0.0 1.4739 0 -2.0 1e-06 
0.0 1.474 0 -2.0 1e-06 
0.0 1.4741 0 -2.0 1e-06 
0.0 1.4742 0 -2.0 1e-06 
0.0 1.4743 0 -2.0 1e-06 
0.0 1.4744 0 -2.0 1e-06 
0.0 1.4745 0 -2.0 1e-06 
0.0 1.4746 0 -2.0 1e-06 
0.0 1.4747 0 -2.0 1e-06 
0.0 1.4748 0 -2.0 1e-06 
0.0 1.4749 0 -2.0 1e-06 
0.0 1.475 0 -2.0 1e-06 
0.0 1.4751 0 -2.0 1e-06 
0.0 1.4752 0 -2.0 1e-06 
0.0 1.4753 0 -2.0 1e-06 
0.0 1.4754 0 -2.0 1e-06 
0.0 1.4755 0 -2.0 1e-06 
0.0 1.4756 0 -2.0 1e-06 
0.0 1.4757 0 -2.0 1e-06 
0.0 1.4758 0 -2.0 1e-06 
0.0 1.4759 0 -2.0 1e-06 
0.0 1.476 0 -2.0 1e-06 
0.0 1.4761 0 -2.0 1e-06 
0.0 1.4762 0 -2.0 1e-06 
0.0 1.4763 0 -2.0 1e-06 
0.0 1.4764 0 -2.0 1e-06 
0.0 1.4765 0 -2.0 1e-06 
0.0 1.4766 0 -2.0 1e-06 
0.0 1.4767 0 -2.0 1e-06 
0.0 1.4768 0 -2.0 1e-06 
0.0 1.4769 0 -2.0 1e-06 
0.0 1.477 0 -2.0 1e-06 
0.0 1.4771 0 -2.0 1e-06 
0.0 1.4772 0 -2.0 1e-06 
0.0 1.4773 0 -2.0 1e-06 
0.0 1.4774 0 -2.0 1e-06 
0.0 1.4775 0 -2.0 1e-06 
0.0 1.4776 0 -2.0 1e-06 
0.0 1.4777 0 -2.0 1e-06 
0.0 1.4778 0 -2.0 1e-06 
0.0 1.4779 0 -2.0 1e-06 
0.0 1.478 0 -2.0 1e-06 
0.0 1.4781 0 -2.0 1e-06 
0.0 1.4782 0 -2.0 1e-06 
0.0 1.4783 0 -2.0 1e-06 
0.0 1.4784 0 -2.0 1e-06 
0.0 1.4785 0 -2.0 1e-06 
0.0 1.4786 0 -2.0 1e-06 
0.0 1.4787 0 -2.0 1e-06 
0.0 1.4788 0 -2.0 1e-06 
0.0 1.4789 0 -2.0 1e-06 
0.0 1.479 0 -2.0 1e-06 
0.0 1.4791 0 -2.0 1e-06 
0.0 1.4792 0 -2.0 1e-06 
0.0 1.4793 0 -2.0 1e-06 
0.0 1.4794 0 -2.0 1e-06 
0.0 1.4795 0 -2.0 1e-06 
0.0 1.4796 0 -2.0 1e-06 
0.0 1.4797 0 -2.0 1e-06 
0.0 1.4798 0 -2.0 1e-06 
0.0 1.4799 0 -2.0 1e-06 
0.0 1.48 0 -2.0 1e-06 
0.0 1.4801 0 -2.0 1e-06 
0.0 1.4802 0 -2.0 1e-06 
0.0 1.4803 0 -2.0 1e-06 
0.0 1.4804 0 -2.0 1e-06 
0.0 1.4805 0 -2.0 1e-06 
0.0 1.4806 0 -2.0 1e-06 
0.0 1.4807 0 -2.0 1e-06 
0.0 1.4808 0 -2.0 1e-06 
0.0 1.4809 0 -2.0 1e-06 
0.0 1.481 0 -2.0 1e-06 
0.0 1.4811 0 -2.0 1e-06 
0.0 1.4812 0 -2.0 1e-06 
0.0 1.4813 0 -2.0 1e-06 
0.0 1.4814 0 -2.0 1e-06 
0.0 1.4815 0 -2.0 1e-06 
0.0 1.4816 0 -2.0 1e-06 
0.0 1.4817 0 -2.0 1e-06 
0.0 1.4818 0 -2.0 1e-06 
0.0 1.4819 0 -2.0 1e-06 
0.0 1.482 0 -2.0 1e-06 
0.0 1.4821 0 -2.0 1e-06 
0.0 1.4822 0 -2.0 1e-06 
0.0 1.4823 0 -2.0 1e-06 
0.0 1.4824 0 -2.0 1e-06 
0.0 1.4825 0 -2.0 1e-06 
0.0 1.4826 0 -2.0 1e-06 
0.0 1.4827 0 -2.0 1e-06 
0.0 1.4828 0 -2.0 1e-06 
0.0 1.4829 0 -2.0 1e-06 
0.0 1.483 0 -2.0 1e-06 
0.0 1.4831 0 -2.0 1e-06 
0.0 1.4832 0 -2.0 1e-06 
0.0 1.4833 0 -2.0 1e-06 
0.0 1.4834 0 -2.0 1e-06 
0.0 1.4835 0 -2.0 1e-06 
0.0 1.4836 0 -2.0 1e-06 
0.0 1.4837 0 -2.0 1e-06 
0.0 1.4838 0 -2.0 1e-06 
0.0 1.4839 0 -2.0 1e-06 
0.0 1.484 0 -2.0 1e-06 
0.0 1.4841 0 -2.0 1e-06 
0.0 1.4842 0 -2.0 1e-06 
0.0 1.4843 0 -2.0 1e-06 
0.0 1.4844 0 -2.0 1e-06 
0.0 1.4845 0 -2.0 1e-06 
0.0 1.4846 0 -2.0 1e-06 
0.0 1.4847 0 -2.0 1e-06 
0.0 1.4848 0 -2.0 1e-06 
0.0 1.4849 0 -2.0 1e-06 
0.0 1.485 0 -2.0 1e-06 
0.0 1.4851 0 -2.0 1e-06 
0.0 1.4852 0 -2.0 1e-06 
0.0 1.4853 0 -2.0 1e-06 
0.0 1.4854 0 -2.0 1e-06 
0.0 1.4855 0 -2.0 1e-06 
0.0 1.4856 0 -2.0 1e-06 
0.0 1.4857 0 -2.0 1e-06 
0.0 1.4858 0 -2.0 1e-06 
0.0 1.4859 0 -2.0 1e-06 
0.0 1.486 0 -2.0 1e-06 
0.0 1.4861 0 -2.0 1e-06 
0.0 1.4862 0 -2.0 1e-06 
0.0 1.4863 0 -2.0 1e-06 
0.0 1.4864 0 -2.0 1e-06 
0.0 1.4865 0 -2.0 1e-06 
0.0 1.4866 0 -2.0 1e-06 
0.0 1.4867 0 -2.0 1e-06 
0.0 1.4868 0 -2.0 1e-06 
0.0 1.4869 0 -2.0 1e-06 
0.0 1.487 0 -2.0 1e-06 
0.0 1.4871 0 -2.0 1e-06 
0.0 1.4872 0 -2.0 1e-06 
0.0 1.4873 0 -2.0 1e-06 
0.0 1.4874 0 -2.0 1e-06 
0.0 1.4875 0 -2.0 1e-06 
0.0 1.4876 0 -2.0 1e-06 
0.0 1.4877 0 -2.0 1e-06 
0.0 1.4878 0 -2.0 1e-06 
0.0 1.4879 0 -2.0 1e-06 
0.0 1.488 0 -2.0 1e-06 
0.0 1.4881 0 -2.0 1e-06 
0.0 1.4882 0 -2.0 1e-06 
0.0 1.4883 0 -2.0 1e-06 
0.0 1.4884 0 -2.0 1e-06 
0.0 1.4885 0 -2.0 1e-06 
0.0 1.4886 0 -2.0 1e-06 
0.0 1.4887 0 -2.0 1e-06 
0.0 1.4888 0 -2.0 1e-06 
0.0 1.4889 0 -2.0 1e-06 
0.0 1.489 0 -2.0 1e-06 
0.0 1.4891 0 -2.0 1e-06 
0.0 1.4892 0 -2.0 1e-06 
0.0 1.4893 0 -2.0 1e-06 
0.0 1.4894 0 -2.0 1e-06 
0.0 1.4895 0 -2.0 1e-06 
0.0 1.4896 0 -2.0 1e-06 
0.0 1.4897 0 -2.0 1e-06 
0.0 1.4898 0 -2.0 1e-06 
0.0 1.4899 0 -2.0 1e-06 
0.0 1.49 0 -2.0 1e-06 
0.0 1.4901 0 -2.0 1e-06 
0.0 1.4902 0 -2.0 1e-06 
0.0 1.4903 0 -2.0 1e-06 
0.0 1.4904 0 -2.0 1e-06 
0.0 1.4905 0 -2.0 1e-06 
0.0 1.4906 0 -2.0 1e-06 
0.0 1.4907 0 -2.0 1e-06 
0.0 1.4908 0 -2.0 1e-06 
0.0 1.4909 0 -2.0 1e-06 
0.0 1.491 0 -2.0 1e-06 
0.0 1.4911 0 -2.0 1e-06 
0.0 1.4912 0 -2.0 1e-06 
0.0 1.4913 0 -2.0 1e-06 
0.0 1.4914 0 -2.0 1e-06 
0.0 1.4915 0 -2.0 1e-06 
0.0 1.4916 0 -2.0 1e-06 
0.0 1.4917 0 -2.0 1e-06 
0.0 1.4918 0 -2.0 1e-06 
0.0 1.4919 0 -2.0 1e-06 
0.0 1.492 0 -2.0 1e-06 
0.0 1.4921 0 -2.0 1e-06 
0.0 1.4922 0 -2.0 1e-06 
0.0 1.4923 0 -2.0 1e-06 
0.0 1.4924 0 -2.0 1e-06 
0.0 1.4925 0 -2.0 1e-06 
0.0 1.4926 0 -2.0 1e-06 
0.0 1.4927 0 -2.0 1e-06 
0.0 1.4928 0 -2.0 1e-06 
0.0 1.4929 0 -2.0 1e-06 
0.0 1.493 0 -2.0 1e-06 
0.0 1.4931 0 -2.0 1e-06 
0.0 1.4932 0 -2.0 1e-06 
0.0 1.4933 0 -2.0 1e-06 
0.0 1.4934 0 -2.0 1e-06 
0.0 1.4935 0 -2.0 1e-06 
0.0 1.4936 0 -2.0 1e-06 
0.0 1.4937 0 -2.0 1e-06 
0.0 1.4938 0 -2.0 1e-06 
0.0 1.4939 0 -2.0 1e-06 
0.0 1.494 0 -2.0 1e-06 
0.0 1.4941 0 -2.0 1e-06 
0.0 1.4942 0 -2.0 1e-06 
0.0 1.4943 0 -2.0 1e-06 
0.0 1.4944 0 -2.0 1e-06 
0.0 1.4945 0 -2.0 1e-06 
0.0 1.4946 0 -2.0 1e-06 
0.0 1.4947 0 -2.0 1e-06 
0.0 1.4948 0 -2.0 1e-06 
0.0 1.4949 0 -2.0 1e-06 
0.0 1.495 0 -2.0 1e-06 
0.0 1.4951 0 -2.0 1e-06 
0.0 1.4952 0 -2.0 1e-06 
0.0 1.4953 0 -2.0 1e-06 
0.0 1.4954 0 -2.0 1e-06 
0.0 1.4955 0 -2.0 1e-06 
0.0 1.4956 0 -2.0 1e-06 
0.0 1.4957 0 -2.0 1e-06 
0.0 1.4958 0 -2.0 1e-06 
0.0 1.4959 0 -2.0 1e-06 
0.0 1.496 0 -2.0 1e-06 
0.0 1.4961 0 -2.0 1e-06 
0.0 1.4962 0 -2.0 1e-06 
0.0 1.4963 0 -2.0 1e-06 
0.0 1.4964 0 -2.0 1e-06 
0.0 1.4965 0 -2.0 1e-06 
0.0 1.4966 0 -2.0 1e-06 
0.0 1.4967 0 -2.0 1e-06 
0.0 1.4968 0 -2.0 1e-06 
0.0 1.4969 0 -2.0 1e-06 
0.0 1.497 0 -2.0 1e-06 
0.0 1.4971 0 -2.0 1e-06 
0.0 1.4972 0 -2.0 1e-06 
0.0 1.4973 0 -2.0 1e-06 
0.0 1.4974 0 -2.0 1e-06 
0.0 1.4975 0 -2.0 1e-06 
0.0 1.4976 0 -2.0 1e-06 
0.0 1.4977 0 -2.0 1e-06 
0.0 1.4978 0 -2.0 1e-06 
0.0 1.4979 0 -2.0 1e-06 
0.0 1.498 0 -2.0 1e-06 
0.0 1.4981 0 -2.0 1e-06 
0.0 1.4982 0 -2.0 1e-06 
0.0 1.4983 0 -2.0 1e-06 
0.0 1.4984 0 -2.0 1e-06 
0.0 1.4985 0 -2.0 1e-06 
0.0 1.4986 0 -2.0 1e-06 
0.0 1.4987 0 -2.0 1e-06 
0.0 1.4988 0 -2.0 1e-06 
0.0 1.4989 0 -2.0 1e-06 
0.0 1.499 0 -2.0 1e-06 
0.0 1.4991 0 -2.0 1e-06 
0.0 1.4992 0 -2.0 1e-06 
0.0 1.4993 0 -2.0 1e-06 
0.0 1.4994 0 -2.0 1e-06 
0.0 1.4995 0 -2.0 1e-06 
0.0 1.4996 0 -2.0 1e-06 
0.0 1.4997 0 -2.0 1e-06 
0.0 1.4998 0 -2.0 1e-06 
0.0 1.4999 0 -2.0 1e-06 
0.0 -1.5 0 2.0 1e-06 
0.0 -1.4999 0 2.0 1e-06 
0.0 -1.4998 0 2.0 1e-06 
0.0 -1.4997 0 2.0 1e-06 
0.0 -1.4996 0 2.0 1e-06 
0.0 -1.4995 0 2.0 1e-06 
0.0 -1.4994 0 2.0 1e-06 
0.0 -1.4993 0 2.0 1e-06 
0.0 -1.4992 0 2.0 1e-06 
0.0 -1.4991 0 2.0 1e-06 
0.0 -1.499 0 2.0 1e-06 
0.0 -1.4989 0 2.0 1e-06 
0.0 -1.4988 0 2.0 1e-06 
0.0 -1.4987 0 2.0 1e-06 
0.0 -1.4986 0 2.0 1e-06 
0.0 -1.4985 0 2.0 1e-06 
0.0 -1.4984 0 2.0 1e-06 
0.0 -1.4983 0 2.0 1e-06 
0.0 -1.4982 0 2.0 1e-06 
0.0 -1.4981 0 2.0 1e-06 
0.0 -1.498 0 2.0 1e-06 
0.0 -1.4979 0 2.0 1e-06 
0.0 -1.4978 0 2.0 1e-06 
0.0 -1.4977 0 2.0 1e-06 
0.0 -1.4976 0 2.0 1e-06 
0.0 -1.4975 0 2.0 1e-06 
0.0 -1.4974 0 2.0 1e-06 
0.0 -1.4973 0 2.0 1e-06 
0.0 -1.4972 0 2.0 1e-06 
0.0 -1.4971 0 2.0 1e-06 
0.0 -1.497 0 2.0 1e-06 
0.0 -1.4969 0 2.0 1e-06 
0.0 -1.4968 0 2.0 1e-06 
0.0 -1.4967 0 2.0 1e-06 
0.0 -1.4966 0 2.0 1e-06 
0.0 -1.4965 0 2.0 1e-06 
0.0 -1.4964 0 2.0 1e-06 
0.0 -1.4963 0 2.0 1e-06 
0.0 -1.4962 0 2.0 1e-06 
0.0 -1.4961 0 2.0 1e-06 
0.0 -1.496 0 2.0 1e-06 
0.0 -1.4959 0 2.0 1e-06 
0.0 -1.4958 0 2.0 1e-06 
0.0 -1.4957 0 2.0 1e-06 
0.0 -1.4956 0 2.0 1e-06 
0.0 -1.4955 0 2.0 1e-06 
0.0 -1.4954 0 2.0 1e-06 
0.0 -1.4953 0 2.0 1e-06 
0.0 -1.4952 0 2.0 1e-06 
0.0 -1.4951 0 2.0 1e-06 
0.0 -1.495 0 2.0 1e-06 
0.0 -1.4949 0 2.0 1e-06 
0.0 -1.4948 0 2.0 1e-06 
0.0 -1.4947 0 2.0 1e-06 
0.0 -1.4946 0 2.0 1e-06 
0.0 -1.4945 0 2.0 1e-06 
0.0 -1.4944 0 2.0 1e-06 
0.0 -1.4943 0 2.0 1e-06 
0.0 -1.4942 0 2.0 1e-06 
0.0 -1.4941 0 2.0 1e-06 
0.0 -1.494 0 2.0 1e-06 
0.0 -1.4939 0 2.0 1e-06 
0.0 -1.4938 0 2.0 1e-06 
0.0 -1.4937 0 2.0 1e-06 
0.0 -1.4936 0 2.0 1e-06 
0.0 -1.4935 0 2.0 1e-06 
0.0 -1.4934 0 2.0 1e-06 
0.0 -1.4933 0 2.0 1e-06 
0.0 -1.4932 0 2.0 1e-06 
0.0 -1.4931 0 2.0 1e-06 
0.0 -1.493 0 2.0 1e-06 
0.0 -1.4929 0 2.0 1e-06 
0.0 -1.4928 0 2.0 1e-06 
0.0 -1.4927 0 2.0 1e-06 
0.0 -1.4926 0 2.0 1e-06 
0.0 -1.4925 0 2.0 1e-06 
0.0 -1.4924 0 2.0 1e-06 
0.0 -1.4923 0 2.0 1e-06 
0.0 -1.4922 0 2.0 1e-06 
0.0 -1.4921 0 2.0 1e-06 
0.0 -1.492 0 2.0 1e-06 
0.0 -1.4919 0 2.0 1e-06 
0.0 -1.4918 0 2.0 1e-06 
0.0 -1.4917 0 2.0 1e-06 
0.0 -1.4916 0 2.0 1e-06 
0.0 -1.4915 0 2.0 1e-06 
0.0 -1.4914 0 2.0 1e-06 
0.0 -1.4913 0 2.0 1e-06 
0.0 -1.4912 0 2.0 1e-06 
0.0 -1.4911 0 2.0 1e-06 
0.0 -1.491 0 2.0 1e-06 
0.0 -1.4909 0 2.0 1e-06 
0.0 -1.4908 0 2.0 1e-06 
0.0 -1.4907 0 2.0 1e-06 
0.0 -1.4906 0 2.0 1e-06 
0.0 -1.4905 0 2.0 1e-06 
0.0 -1.4904 0 2.0 1e-06 
0.0 -1.4903 0 2.0 1e-06 
0.0 -1.4902 0 2.0 1e-06 
0.0 -1.4901 0 2.0 1e-06 
0.0 -1.49 0 2.0 1e-06 
0.0 -1.4899 0 2.0 1e-06 
0.0 -1.4898 0 2.0 1e-06 
0.0 -1.4897 0 2.0 1e-06 
0.0 -1.4896 0 2.0 1e-06 
0.0 -1.4895 0 2.0 1e-06 
0.0 -1.4894 0 2.0 1e-06 
0.0 -1.4893 0 2.0 1e-06 
0.0 -1.4892 0 2.0 1e-06 
0.0 -1.4891 0 2.0 1e-06 
0.0 -1.489 0 2.0 1e-06 
0.0 -1.4889 0 2.0 1e-06 
0.0 -1.4888 0 2.0 1e-06 
0.0 -1.4887 0 2.0 1e-06 
0.0 -1.4886 0 2.0 1e-06 
0.0 -1.4885 0 2.0 1e-06 
0.0 -1.4884 0 2.0 1e-06 
0.0 -1.4883 0 2.0 1e-06 
0.0 -1.4882 0 2.0 1e-06 
0.0 -1.4881 0 2.0 1e-06 
0.0 -1.488 0 2.0 1e-06 
0.0 -1.4879 0 2.0 1e-06 
0.0 -1.4878 0 2.0 1e-06 
0.0 -1.4877 0 2.0 1e-06 
0.0 -1.4876 0 2.0 1e-06 
0.0 -1.4875 0 2.0 1e-06 
0.0 -1.4874 0 2.0 1e-06 
0.0 -1.4873 0 2.0 1e-06 
0.0 -1.4872 0 2.0 1e-06 
0.0 -1.4871 0 2.0 1e-06 
0.0 -1.487 0 2.0 1e-06 
0.0 -1.4869 0 2.0 1e-06 
0.0 -1.4868 0 2.0 1e-06 
0.0 -1.4867 0 2.0 1e-06 
0.0 -1.4866 0 2.0 1e-06 
0.0 -1.4865 0 2.0 1e-06 
0.0 -1.4864 0 2.0 1e-06 
0.0 -1.4863 0 2.0 1e-06 
0.0 -1.4862 0 2.0 1e-06 
0.0 -1.4861 0 2.0 1e-06 
0.0 -1.486 0 2.0 1e-06 
0.0 -1.4859 0 2.0 1e-06 
0.0 -1.4858 0 2.0 1e-06 
0.0 -1.4857 0 2.0 1e-06 
0.0 -1.4856 0 2.0 1e-06 
0.0 -1.4855 0 2.0 1e-06 
0.0 -1.4854 0 2.0 1e-06 
0.0 -1.4853 0 2.0 1e-06 
0.0 -1.4852 0 2.0 1e-06 
0.0 -1.4851 0 2.0 1e-06 
0.0 -1.485 0 2.0 1e-06 
0.0 -1.4849 0 2.0 1e-06 
0.0 -1.4848 0 2.0 1e-06 
0.0 -1.4847 0 2.0 1e-06 
0.0 -1.4846 0 2.0 1e-06 
0.0 -1.4845 0 2.0 1e-06 
0.0 -1.4844 0 2.0 1e-06 
0.0 -1.4843 0 2.0 1e-06 
0.0 -1.4842 0 2.0 1e-06 
0.0 -1.4841 0 2.0 1e-06 
0.0 -1.484 0 2.0 1e-06 
0.0 -1.4839 0 2.0 1e-06 
0.0 -1.4838 0 2.0 1e-06 
0.0 -1.4837 0 2.0 1e-06 
0.0 -1.4836 0 2.0 1e-06 
0.0 -1.4835 0 2.0 1e-06 
0.0 -1.4834 0 2.0 1e-06 
0.0 -1.4833 0 2.0 1e-06 
0.0 -1.4832 0 2.0 1e-06 
0.0 -1.4831 0 2.0 1e-06 
0.0 -1.483 0 2.0 1e-06 
0.0 -1.4829 0 2.0 1e-06 
0.0 -1.4828 0 2.0 1e-06 
0.0 -1.4827 0 2.0 1e-06 
0.0 -1.4826 0 2.0 1e-06 
0.0 -1.4825 0 2.0 1e-06 
0.0 -1.4824 0 2.0 1e-06 
0.0 -1.4823 0 2.0 1e-06 
0.0 -1.4822 0 2.0 1e-06 
0.0 -1.4821 0 2.0 1e-06 
0.0 -1.482 0 2.0 1e-06 
0.0 -1.4819 0 2.0 1e-06 
0.0 -1.4818 0 2.0 1e-06 
0.0 -1.4817 0 2.0 1e-06 
0.0 -1.4816 0 2.0 1e-06 
0.0 -1.4815 0 2.0 1e-06 
0.0 -1.4814 0 2.0 1e-06 
0.0 -1.4813 0 2.0 1e-06 
0.0 -1.4812 0 2.0 1e-06 
0.0 -1.4811 0 2.0 1e-06 
0.0 -1.481 0 2.0 1e-06 
0.0 -1.4809 0 2.0 1e-06 
0.0 -1.4808 0 2.0 1e-06 
0.0 -1.4807 0 2.0 1e-06 
0.0 -1.4806 0 2.0 1e-06 
0.0 -1.4805 0 2.0 1e-06 
0.0 -1.4804 0 2.0 1e-06 
0.0 -1.4803 0 2.0 1e-06 
0.0 -1.4802 0 2.0 1e-06 
0.0 -1.4801 0 2.0 1e-06 
0.0 -1.48 0 2.0 1e-06 
0.0 -1.4799 0 2.0 1e-06 
0.0 -1.4798 0 2.0 1e-06 
0.0 -1.4797 0 2.0 1e-06 
0.0 -1.4796 0 2.0 1e-06 
0.0 -1.4795 0 2.0 1e-06 
0.0 -1.4794 0 2.0 1e-06 
0.0 -1.4793 0 2.0 1e-06 
0.0 -1.4792 0 2.0 1e-06 
0.0 -1.4791 0 2.0 1e-06 
0.0 -1.479 0 2.0 1e-06 
0.0 -1.4789 0 2.0 1e-06 
0.0 -1.4788 0 2.0 1e-06 
0.0 -1.4787 0 2.0 1e-06 
0.0 -1.4786 0 2.0 1e-06 
0.0 -1.4785 0 2.0 1e-06 
0.0 -1.4784 0 2.0 1e-06 
0.0 -1.4783 0 2.0 1e-06 
0.0 -1.4782 0 2.0 1e-06 
0.0 -1.4781 0 2.0 1e-06 
0.0 -1.478 0 2.0 1e-06 
0.0 -1.4779 0 2.0 1e-06 
0.0 -1.4778 0 2.0 1e-06 
0.0 -1.4777 0 2.0 1e-06 
0.0 -1.4776 0 2.0 1e-06 
0.0 -1.4775 0 2.0 1e-06 
0.0 -1.4774 0 2.0 1e-06 
0.0 -1.4773 0 2.0 1e-06 
0.0 -1.4772 0 2.0 1e-06 
0.0 -1.4771 0 2.0 1e-06 
0.0 -1.477 0 2.0 1e-06 
0.0 -1.4769 0 2.0 1e-06 
0.0 -1.4768 0 2.0 1e-06 
0.0 -1.4767 0 2.0 1e-06 
0.0 -1.4766 0 2.0 1e-06 
0.0 -1.4765 0 2.0 1e-06 
0.0 -1.4764 0 2.0 1e-06 
0.0 -1.4763 0 2.0 1e-06 
0.0 -1.4762 0 2.0 1e-06 
0.0 -1.4761 0 2.0 1e-06 
0.0 -1.476 0 2.0 1e-06 
0.0 -1.4759 0 2.0 1e-06 
0.0 -1.4758 0 2.0 1e-06 
0.0 -1.4757 0 2.0 1e-06 
0.0 -1.4756 0 2.0 1e-06 
0.0 -1.4755 0 2.0 1e-06 
0.0 -1.4754 0 2.0 1e-06 
0.0 -1.4753 0 2.0 1e-06 
0.0 -1.4752 0 2.0 1e-06 
0.0 -1.4751 0 2.0 1e-06 
0.0 -1.475 0 2.0 1e-06 
0.0 -1.4749 0 2.0 1e-06 
0.0 -1.4748 0 2.0 1e-06 
0.0 -1.4747 0 2.0 1e-06 
0.0 -1.4746 0 2.0 1e-06 
0.0 -1.4745 0 2.0 1e-06 
0.0 -1.4744 0 2.0 1e-06 
0.0 -1.4743 0 2.0 1e-06 
0.0 -1.4742 0 2.0 1e-06 
0.0 -1.4741 0 2.0 1e-06 
0.0 -1.474 0 2.0 1e-06 
0.0 -1.4739 0 2.0 1e-06 
0.0 -1.4738 0 2.0 1e-06 
0.0 -1.4737 0 2.0 1e-06 
0.0 -1.4736 0 2.0 1e-06 
0.0 -1.4735 0 2.0 1e-06 
0.0 -1.4734 0 2.0 1e-06 
0.0 -1.4733 0 2.0 1e-06 
0.0 -1.4732 0 2.0 1e-06 
0.0 -1.4731 0 2.0 1e-06 
0.0 -1.473 0 2.0 1e-06 
0.0 -1.4729 0 2.0 1e-06 
0.0 -1.4728 0 2.0 1e-06 
0.0 -1.4727 0 2.0 1e-06 
0.0 -1.4726 0 2.0 1e-06 
0.0 -1.4725 0 2.0 1e-06 
0.0 -1.4724 0 2.0 1e-06 
0.0 -1.4723 0 2.0 1e-06 
0.0 -1.4722 0 2.0 1e-06 
0.0 -1.4721 0 2.0 1e-06 
0.0 -1.472 0 2.0 1e-06 
0.0 -1.4719 0 2.0 1e-06 
0.0 -1.4718 0 2.0 1e-06 
0.0 -1.4717 0 2.0 1e-06 
0.0 -1.4716 0 2.0 1e-06 
0.0 -1.4715 0 2.0 1e-06 
0.0 -1.4714 0 2.0 1e-06 
0.0 -1.4713 0 2.0 1e-06 
0.0 -1.4712 0 2.0 1e-06 
0.0 -1.4711 0 2.0 1e-06 
0.0 -1.471 0 2.0 1e-06 
0.0 -1.4709 0 2.0 1e-06 
0.0 -1.4708 0 2.0 1e-06 
0.0 -1.4707 0 2.0 1e-06 
0.0 -1.4706 0 2.0 1e-06 
0.0 -1.4705 0 2.0 1e-06 
0.0 -1.4704 0 2.0 1e-06 
0.0 -1.4703 0 2.0 1e-06 
0.0 -1.4702 0 2.0 1e-06 
0.0 -1.4701 0 2.0 1e-06 
0.0 -1.47 0 2.0 1e-06 
0.0 -1.4699 0 2.0 1e-06 
0.0 -1.4698 0 2.0 1e-06 
0.0 -1.4697 0 2.0 1e-06 
0.0 -1.4696 0 2.0 1e-06 
0.0 -1.4695 0 2.0 1e-06 
0.0 -1.4694 0 2.0 1e-06 
0.0 -1.4693 0 2.0 1e-06 
0.0 -1.4692 0 2.0 1e-06 
0.0 -1.4691 0 2.0 1e-06 
0.0 -1.469 0 2.0 1e-06 
0.0 -1.4689 0 2.0 1e-06 
0.0 -1.4688 0 2.0 1e-06 
0.0 -1.4687 0 2.0 1e-06 
0.0 -1.4686 0 2.0 1e-06 
0.0 -1.4685 0 2.0 1e-06 
0.0 -1.4684 0 2.0 1e-06 
0.0 -1.4683 0 2.0 1e-06 
0.0 -1.4682 0 2.0 1e-06 
0.0 -1.4681 0 2.0 1e-06 
0.0 -1.468 0 2.0 1e-06 
0.0 -1.4679 0 2.0 1e-06 
0.0 -1.4678 0 2.0 1e-06 
0.0 -1.4677 0 2.0 1e-06 
0.0 -1.4676 0 2.0 1e-06 
0.0 -1.4675 0 2.0 1e-06 
0.0 -1.4674 0 2.0 1e-06 
0.0 -1.4673 0 2.0 1e-06 
0.0 -1.4672 0 2.0 1e-06 
0.0 -1.4671 0 2.0 1e-06 
0.0 -1.467 0 2.0 1e-06 
0.0 -1.4669 0 2.0 1e-06 
0.0 -1.4668 0 2.0 1e-06 
0.0 -1.4667 0 2.0 1e-06 
0.0 -1.4666 0 2.0 1e-06 
0.0 -1.4665 0 2.0 1e-06 
0.0 -1.4664 0 2.0 1e-06 
0.0 -1.4663 0 2.0 1e-06 
0.0 -1.4662 0 2.0 1e-06 
0.0 -1.4661 0 2.0 1e-06 
0.0 -1.466 0 2.0 1e-06 
0.0 -1.4659 0 2.0 1e-06 
0.0 -1.4658 0 2.0 1e-06 
0.0 -1.4657 0 2.0 1e-06 
0.0 -1.4656 0 2.0 1e-06 
0.0 -1.4655 0 2.0 1e-06 
0.0 -1.4654 0 2.0 1e-06 
0.0 -1.4653 0 2.0 1e-06 
0.0 -1.4652 0 2.0 1e-06 
0.0 -1.4651 0 2.0 1e-06 
0.0 -1.465 0 2.0 1e-06 
0.0 -1.4649 0 2.0 1e-06 
0.0 -1.4648 0 2.0 1e-06 
0.0 -1.4647 0 2.0 1e-06 
0.0 -1.4646 0 2.0 1e-06 
0.0 -1.4645 0 2.0 1e-06 
0.0 -1.4644 0 2.0 1e-06 
0.0 -1.4643 0 2.0 1e-06 
0.0 -1.4642 0 2.0 1e-06 
0.0 -1.4641 0 2.0 1e-06 
0.0 -1.464 0 2.0 1e-06 
0.0 -1.4639 0 2.0 1e-06 
0.0 -1.4638 0 2.0 1e-06 
0.0 -1.4637 0 2.0 1e-06 
0.0 -1.4636 0 2.0 1e-06 
0.0 -1.4635 0 2.0 1e-06 
0.0 -1.4634 0 2.0 1e-06 
0.0 -1.4633 0 2.0 1e-06 
0.0 -1.4632 0 2.0 1e-06 
0.0 -1.4631 0 2.0 1e-06 
0.0 -1.463 0 2.0 1e-06 
0.0 -1.4629 0 2.0 1e-06 
0.0 -1.4628 0 2.0 1e-06 
0.0 -1.4627 0 2.0 1e-06 
0.0 -1.4626 0 2.0 1e-06 
0.0 -1.4625 0 2.0 1e-06 
0.0 -1.4624 0 2.0 1e-06 
0.0 -1.4623 0 2.0 1e-06 
0.0 -1.4622 0 2.0 1e-06 
0.0 -1.4621 0 2.0 1e-06 
0.0 -1.462 0 2.0 1e-06 
0.0 -1.4619 0 2.0 1e-06 
0.0 -1.4618 0 2.0 1e-06 
0.0 -1.4617 0 2.0 1e-06 
0.0 -1.4616 0 2.0 1e-06 
0.0 -1.4615 0 2.0 1e-06 
0.0 -1.4614 0 2.0 1e-06 
0.0 -1.4613 0 2.0 1e-06 
0.0 -1.4612 0 2.0 1e-06 
0.0 -1.4611 0 2.0 1e-06 
0.0 -1.461 0 2.0 1e-06 
0.0 -1.4609 0 2.0 1e-06 
0.0 -1.4608 0 2.0 1e-06 
0.0 -1.4607 0 2.0 1e-06 
0.0 -1.4606 0 2.0 1e-06 
0.0 -1.4605 0 2.0 1e-06 
0.0 -1.4604 0 2.0 1e-06 
0.0 -1.4603 0 2.0 1e-06 
0.0 -1.4602 0 2.0 1e-06 
0.0 -1.4601 0 2.0 1e-06 
0.0 -1.46 0 2.0 1e-06 
0.0 -1.4599 0 2.0 1e-06 
0.0 -1.4598 0 2.0 1e-06 
0.0 -1.4597 0 2.0 1e-06 
0.0 -1.4596 0 2.0 1e-06 
0.0 -1.4595 0 2.0 1e-06 
0.0 -1.4594 0 2.0 1e-06 
0.0 -1.4593 0 2.0 1e-06 
0.0 -1.4592 0 2.0 1e-06 
0.0 -1.4591 0 2.0 1e-06 
0.0 -1.459 0 2.0 1e-06 
0.0 -1.4589 0 2.0 1e-06 
0.0 -1.4588 0 2.0 1e-06 
0.0 -1.4587 0 2.0 1e-06 
0.0 -1.4586 0 2.0 1e-06 
0.0 -1.4585 0 2.0 1e-06 
0.0 -1.4584 0 2.0 1e-06 
0.0 -1.4583 0 2.0 1e-06 
0.0 -1.4582 0 2.0 1e-06 
0.0 -1.4581 0 2.0 1e-06 
0.0 -1.458 0 2.0 1e-06 
0.0 -1.4579 0 2.0 1e-06 
0.0 -1.4578 0 2.0 1e-06 
0.0 -1.4577 0 2.0 1e-06 
0.0 -1.4576 0 2.0 1e-06 
0.0 -1.4575 0 2.0 1e-06 
0.0 -1.4574 0 2.0 1e-06 
0.0 -1.4573 0 2.0 1e-06 
0.0 -1.4572 0 2.0 1e-06 
0.0 -1.4571 0 2.0 1e-06 
0.0 -1.457 0 2.0 1e-06 
0.0 -1.4569 0 2.0 1e-06 
0.0 -1.4568 0 2.0 1e-06 
0.0 -1.4567 0 2.0 1e-06 
0.0 -1.4566 0 2.0 1e-06 
0.0 -1.4565 0 2.0 1e-06 
0.0 -1.4564 0 2.0 1e-06 
0.0 -1.4563 0 2.0 1e-06 
0.0 -1.4562 0 2.0 1e-06 
0.0 -1.4561 0 2.0 1e-06 
0.0 -1.456 0 2.0 1e-06 
0.0 -1.4559 0 2.0 1e-06 
0.0 -1.4558 0 2.0 1e-06 
0.0 -1.4557 0 2.0 1e-06 
0.0 -1.4556 0 2.0 1e-06 
0.0 -1.4555 0 2.0 1e-06 
0.0 -1.4554 0 2.0 1e-06 
0.0 -1.4553 0 2.0 1e-06 
0.0 -1.4552 0 2.0 1e-06 
0.0 -1.4551 0 2.0 1e-06 
0.0 -1.455 0 2.0 1e-06 
0.0 -1.4549 0 2.0 1e-06 
0.0 -1.4548 0 2.0 1e-06 
0.0 -1.4547 0 2.0 1e-06 
0.0 -1.4546 0 2.0 1e-06 
0.0 -1.4545 0 2.0 1e-06 
0.0 -1.4544 0 2.0 1e-06 
0.0 -1.4543 0 2.0 1e-06 
0.0 -1.4542 0 2.0 1e-06 
0.0 -1.4541 0 2.0 1e-06 
0.0 -1.454 0 2.0 1e-06 
0.0 -1.4539 0 2.0 1e-06 
0.0 -1.4538 0 2.0 1e-06 
0.0 -1.4537 0 2.0 1e-06 
0.0 -1.4536 0 2.0 1e-06 
0.0 -1.4535 0 2.0 1e-06 
0.0 -1.4534 0 2.0 1e-06 
0.0 -1.4533 0 2.0 1e-06 
0.0 -1.4532 0 2.0 1e-06 
0.0 -1.4531 0 2.0 1e-06 
0.0 -1.453 0 2.0 1e-06 
0.0 -1.4529 0 2.0 1e-06 
0.0 -1.4528 0 2.0 1e-06 
0.0 -1.4527 0 2.0 1e-06 
0.0 -1.4526 0 2.0 1e-06 
0.0 -1.4525 0 2.0 1e-06 
0.0 -1.4524 0 2.0 1e-06 
0.0 -1.4523 0 2.0 1e-06 
0.0 -1.4522 0 2.0 1e-06 
0.0 -1.4521 0 2.0 1e-06 
0.0 -1.452 0 2.0 1e-06 
0.0 -1.4519 0 2.0 1e-06 
0.0 -1.4518 0 2.0 1e-06 
0.0 -1.4517 0 2.0 1e-06 
0.0 -1.4516 0 2.0 1e-06 
0.0 -1.4515 0 2.0 1e-06 
0.0 -1.4514 0 2.0 1e-06 
0.0 -1.4513 0 2.0 1e-06 
0.0 -1.4512 0 2.0 1e-06 
0.0 -1.4511 0 2.0 1e-06 
0.0 -1.451 0 2.0 1e-06 
0.0 -1.4509 0 2.0 1e-06 
0.0 -1.4508 0 2.0 1e-06 
0.0 -1.4507 0 2.0 1e-06 
0.0 -1.4506 0 2.0 1e-06 
0.0 -1.4505 0 2.0 1e-06 
0.0 -1.4504 0 2.0 1e-06 
0.0 -1.4503 0 2.0 1e-06 
0.0 -1.4502 0 2.0 1e-06 
0.0 -1.4501 0 2.0 1e-06 
0.0 -1.45 0 2.0 1e-06 
0.0 -1.4499 0 2.0 1e-06 
0.0 -1.4498 0 2.0 1e-06 
0.0 -1.4497 0 2.0 1e-06 
0.0 -1.4496 0 2.0 1e-06 
0.0 -1.4495 0 2.0 1e-06 
0.0 -1.4494 0 2.0 1e-06 
0.0 -1.4493 0 2.0 1e-06 
0.0 -1.4492 0 2.0 1e-06 
0.0 -1.4491 0 2.0 1e-06 
0.0 -1.449 0 2.0 1e-06 
0.0 -1.4489 0 2.0 1e-06 
0.0 -1.4488 0 2.0 1e-06 
0.0 -1.4487 0 2.0 1e-06 
0.0 -1.4486 0 2.0 1e-06 
0.0 -1.4485 0 2.0 1e-06 
0.0 -1.4484 0 2.0 1e-06 
0.0 -1.4483 0 2.0 1e-06 
0.0 -1.4482 0 2.0 1e-06 
0.0 -1.4481 0 2.0 1e-06 
0.0 -1.448 0 2.0 1e-06 
0.0 -1.4479 0 2.0 1e-06 
0.0 -1.4478 0 2.0 1e-06 
0.0 -1.4477 0 2.0 1e-06 
0.0 -1.4476 0 2.0 1e-06 
0.0 -1.4475 0 2.0 1e-06 
0.0 -1.4474 0 2.0 1e-06 
0.0 -1.4473 0 2.0 1e-06 
0.0 -1.4472 0 2.0 1e-06 
0.0 -1.4471 0 2.0 1e-06 
0.0 -1.447 0 2.0 1e-06 
0.0 -1.4469 0 2.0 1e-06 
0.0 -1.4468 0 2.0 1e-06 
0.0 -1.4467 0 2.0 1e-06 
0.0 -1.4466 0 2.0 1e-06 
0.0 -1.4465 0 2.0 1e-06 
0.0 -1.4464 0 2.0 1e-06 
0.0 -1.4463 0 2.0 1e-06 
0.0 -1.4462 0 2.0 1e-06 
0.0 -1.4461 0 2.0 1e-06 
0.0 -1.446 0 2.0 1e-06 
0.0 -1.4459 0 2.0 1e-06 
0.0 -1.4458 0 2.0 1e-06 
0.0 -1.4457 0 2.0 1e-06 
0.0 -1.4456 0 2.0 1e-06 
0.0 -1.4455 0 2.0 1e-06 
0.0 -1.4454 0 2.0 1e-06 
0.0 -1.4453 0 2.0 1e-06 
0.0 -1.4452 0 2.0 1e-06 
0.0 -1.4451 0 2.0 1e-06 
0.0 -1.445 0 2.0 1e-06 
0.0 -1.4449 0 2.0 1e-06 
0.0 -1.4448 0 2.0 1e-06 
0.0 -1.4447 0 2.0 1e-06 
0.0 -1.4446 0 2.0 1e-06 
0.0 -1.4445 0 2.0 1e-06 
0.0 -1.4444 0 2.0 1e-06 
0.0 -1.4443 0 2.0 1e-06 
0.0 -1.4442 0 2.0 1e-06 
0.0 -1.4441 0 2.0 1e-06 
0.0 -1.444 0 2.0 1e-06 
0.0 -1.4439 0 2.0 1e-06 
0.0 -1.4438 0 2.0 1e-06 
0.0 -1.4437 0 2.0 1e-06 
0.0 -1.4436 0 2.0 1e-06 
0.0 -1.4435 0 2.0 1e-06 
0.0 -1.4434 0 2.0 1e-06 
0.0 -1.4433 0 2.0 1e-06 
0.0 -1.4432 0 2.0 1e-06 
0.0 -1.4431 0 2.0 1e-06 
0.0 -1.443 0 2.0 1e-06 
0.0 -1.4429 0 2.0 1e-06 
0.0 -1.4428 0 2.0 1e-06 
0.0 -1.4427 0 2.0 1e-06 
0.0 -1.4426 0 2.0 1e-06 
0.0 -1.4425 0 2.0 1e-06 
0.0 -1.4424 0 2.0 1e-06 
0.0 -1.4423 0 2.0 1e-06 
0.0 -1.4422 0 2.0 1e-06 
0.0 -1.4421 0 2.0 1e-06 
0.0 -1.442 0 2.0 1e-06 
0.0 -1.4419 0 2.0 1e-06 
0.0 -1.4418 0 2.0 1e-06 
0.0 -1.4417 0 2.0 1e-06 
0.0 -1.4416 0 2.0 1e-06 
0.0 -1.4415 0 2.0 1e-06 
0.0 -1.4414 0 2.0 1e-06 
0.0 -1.4413 0 2.0 1e-06 
0.0 -1.4412 0 2.0 1e-06 
0.0 -1.4411 0 2.0 1e-06 
0.0 -1.441 0 2.0 1e-06 
0.0 -1.4409 0 2.0 1e-06 
0.0 -1.4408 0 2.0 1e-06 
0.0 -1.4407 0 2.0 1e-06 
0.0 -1.4406 0 2.0 1e-06 
0.0 -1.4405 0 2.0 1e-06 
0.0 -1.4404 0 2.0 1e-06 
0.0 -1.4403 0 2.0 1e-06 
0.0 -1.4402 0 2.0 1e-06 
0.0 -1.4401 0 2.0 1e-06 
0.0 -1.44 0 2.0 1e-06 
0.0 -1.4399 0 2.0 1e-06 
0.0 -1.4398 0 2.0 1e-06 
0.0 -1.4397 0 2.0 1e-06 
0.0 -1.4396 0 2.0 1e-06 
0.0 -1.4395 0 2.0 1e-06 
0.0 -1.4394 0 2.0 1e-06 
0.0 -1.4393 0 2.0 1e-06 
0.0 -1.4392 0 2.0 1e-06 
0.0 -1.4391 0 2.0 1e-06 
0.0 -1.439 0 2.0 1e-06 
0.0 -1.4389 0 2.0 1e-06 
0.0 -1.4388 0 2.0 1e-06 
0.0 -1.4387 0 2.0 1e-06 
0.0 -1.4386 0 2.0 1e-06 
0.0 -1.4385 0 2.0 1e-06 
0.0 -1.4384 0 2.0 1e-06 
0.0 -1.4383 0 2.0 1e-06 
0.0 -1.4382 0 2.0 1e-06 
0.0 -1.4381 0 2.0 1e-06 
0.0 -1.438 0 2.0 1e-06 
0.0 -1.4379 0 2.0 1e-06 
0.0 -1.4378 0 2.0 1e-06 
0.0 -1.4377 0 2.0 1e-06 
0.0 -1.4376 0 2.0 1e-06 
0.0 -1.4375 0 2.0 1e-06 
0.0 -1.4374 0 2.0 1e-06 
0.0 -1.4373 0 2.0 1e-06 
0.0 -1.4372 0 2.0 1e-06 
0.0 -1.4371 0 2.0 1e-06 
0.0 -1.437 0 2.0 1e-06 
0.0 -1.4369 0 2.0 1e-06 
0.0 -1.4368 0 2.0 1e-06 
0.0 -1.4367 0 2.0 1e-06 
0.0 -1.4366 0 2.0 1e-06 
0.0 -1.4365 0 2.0 1e-06 
0.0 -1.4364 0 2.0 1e-06 
0.0 -1.4363 0 2.0 1e-06 
0.0 -1.4362 0 2.0 1e-06 
0.0 -1.4361 0 2.0 1e-06 
0.0 -1.436 0 2.0 1e-06 
0.0 -1.4359 0 2.0 1e-06 
0.0 -1.4358 0 2.0 1e-06 
0.0 -1.4357 0 2.0 1e-06 
0.0 -1.4356 0 2.0 1e-06 
0.0 -1.4355 0 2.0 1e-06 
0.0 -1.4354 0 2.0 1e-06 
0.0 -1.4353 0 2.0 1e-06 
0.0 -1.4352 0 2.0 1e-06 
0.0 -1.4351 0 2.0 1e-06 
0.0 -1.435 0 2.0 1e-06 
0.0 -1.4349 0 2.0 1e-06 
0.0 -1.4348 0 2.0 1e-06 
0.0 -1.4347 0 2.0 1e-06 
0.0 -1.4346 0 2.0 1e-06 
0.0 -1.4345 0 2.0 1e-06 
0.0 -1.4344 0 2.0 1e-06 
0.0 -1.4343 0 2.0 1e-06 
0.0 -1.4342 0 2.0 1e-06 
0.0 -1.4341 0 2.0 1e-06 
0.0 -1.434 0 2.0 1e-06 
0.0 -1.4339 0 2.0 1e-06 
0.0 -1.4338 0 2.0 1e-06 
0.0 -1.4337 0 2.0 1e-06 
0.0 -1.4336 0 2.0 1e-06 
0.0 -1.4335 0 2.0 1e-06 
0.0 -1.4334 0 2.0 1e-06 
0.0 -1.4333 0 2.0 1e-06 
0.0 -1.4332 0 2.0 1e-06 
0.0 -1.4331 0 2.0 1e-06 
0.0 -1.433 0 2.0 1e-06 
0.0 -1.4329 0 2.0 1e-06 
0.0 -1.4328 0 2.0 1e-06 
0.0 -1.4327 0 2.0 1e-06 
0.0 -1.4326 0 2.0 1e-06 
0.0 -1.4325 0 2.0 1e-06 
0.0 -1.4324 0 2.0 1e-06 
0.0 -1.4323 0 2.0 1e-06 
0.0 -1.4322 0 2.0 1e-06 
0.0 -1.4321 0 2.0 1e-06 
0.0 -1.432 0 2.0 1e-06 
0.0 -1.4319 0 2.0 1e-06 
0.0 -1.4318 0 2.0 1e-06 
0.0 -1.4317 0 2.0 1e-06 
0.0 -1.4316 0 2.0 1e-06 
0.0 -1.4315 0 2.0 1e-06 
0.0 -1.4314 0 2.0 1e-06 
0.0 -1.4313 0 2.0 1e-06 
0.0 -1.4312 0 2.0 1e-06 
0.0 -1.4311 0 2.0 1e-06 
0.0 -1.431 0 2.0 1e-06 
0.0 -1.4309 0 2.0 1e-06 
0.0 -1.4308 0 2.0 1e-06 
0.0 -1.4307 0 2.0 1e-06 
0.0 -1.4306 0 2.0 1e-06 
0.0 -1.4305 0 2.0 1e-06 
0.0 -1.4304 0 2.0 1e-06 
0.0 -1.4303 0 2.0 1e-06 
0.0 -1.4302 0 2.0 1e-06 
0.0 -1.4301 0 2.0 1e-06 
0.0 -1.43 0 2.0 1e-06 
0.0 -1.4299 0 2.0 1e-06 
0.0 -1.4298 0 2.0 1e-06 
0.0 -1.4297 0 2.0 1e-06 
0.0 -1.4296 0 2.0 1e-06 
0.0 -1.4295 0 2.0 1e-06 
0.0 -1.4294 0 2.0 1e-06 
0.0 -1.4293 0 2.0 1e-06 
0.0 -1.4292 0 2.0 1e-06 
0.0 -1.4291 0 2.0 1e-06 
0.0 -1.429 0 2.0 1e-06 
0.0 -1.4289 0 2.0 1e-06 
0.0 -1.4288 0 2.0 1e-06 
0.0 -1.4287 0 2.0 1e-06 
0.0 -1.4286 0 2.0 1e-06 
0.0 -1.4285 0 2.0 1e-06 
0.0 -1.4284 0 2.0 1e-06 
0.0 -1.4283 0 2.0 1e-06 
0.0 -1.4282 0 2.0 1e-06 
0.0 -1.4281 0 2.0 1e-06 
0.0 -1.428 0 2.0 1e-06 
0.0 -1.4279 0 2.0 1e-06 
0.0 -1.4278 0 2.0 1e-06 
0.0 -1.4277 0 2.0 1e-06 
0.0 -1.4276 0 2.0 1e-06 
0.0 -1.4275 0 2.0 1e-06 
0.0 -1.4274 0 2.0 1e-06 
0.0 -1.4273 0 2.0 1e-06 
0.0 -1.4272 0 2.0 1e-06 
0.0 -1.4271 0 2.0 1e-06 
0.0 -1.427 0 2.0 1e-06 
0.0 -1.4269 0 2.0 1e-06 
0.0 -1.4268 0 2.0 1e-06 
0.0 -1.4267 0 2.0 1e-06 
0.0 -1.4266 0 2.0 1e-06 
0.0 -1.4265 0 2.0 1e-06 
0.0 -1.4264 0 2.0 1e-06 
0.0 -1.4263 0 2.0 1e-06 
0.0 -1.4262 0 2.0 1e-06 
0.0 -1.4261 0 2.0 1e-06 
0.0 -1.426 0 2.0 1e-06 
0.0 -1.4259 0 2.0 1e-06 
0.0 -1.4258 0 2.0 1e-06 
0.0 -1.4257 0 2.0 1e-06 
0.0 -1.4256 0 2.0 1e-06 
0.0 -1.4255 0 2.0 1e-06 
0.0 -1.4254 0 2.0 1e-06 
0.0 -1.4253 0 2.0 1e-06 
0.0 -1.4252 0 2.0 1e-06 
0.0 -1.4251 0 2.0 1e-06 
0.0 -1.425 0 2.0 1e-06 
0.0 -1.4249 0 2.0 1e-06 
0.0 -1.4248 0 2.0 1e-06 
0.0 -1.4247 0 2.0 1e-06 
0.0 -1.4246 0 2.0 1e-06 
0.0 -1.4245 0 2.0 1e-06 
0.0 -1.4244 0 2.0 1e-06 
0.0 -1.4243 0 2.0 1e-06 
0.0 -1.4242 0 2.0 1e-06 
0.0 -1.4241 0 2.0 1e-06 
0.0 -1.424 0 2.0 1e-06 
0.0 -1.4239 0 2.0 1e-06 
0.0 -1.4238 0 2.0 1e-06 
0.0 -1.4237 0 2.0 1e-06 
0.0 -1.4236 0 2.0 1e-06 
0.0 -1.4235 0 2.0 1e-06 
0.0 -1.4234 0 2.0 1e-06 
0.0 -1.4233 0 2.0 1e-06 
0.0 -1.4232 0 2.0 1e-06 
0.0 -1.4231 0 2.0 1e-06 
0.0 -1.423 0 2.0 1e-06 
0.0 -1.4229 0 2.0 1e-06 
0.0 -1.4228 0 2.0 1e-06 
0.0 -1.4227 0 2.0 1e-06 
0.0 -1.4226 0 2.0 1e-06 
0.0 -1.4225 0 2.0 1e-06 
0.0 -1.4224 0 2.0 1e-06 
0.0 -1.4223 0 2.0 1e-06 
0.0 -1.4222 0 2.0 1e-06 
0.0 -1.4221 0 2.0 1e-06 
0.0 -1.422 0 2.0 1e-06 
0.0 -1.4219 0 2.0 1e-06 
0.0 -1.4218 0 2.0 1e-06 
0.0 -1.4217 0 2.0 1e-06 
0.0 -1.4216 0 2.0 1e-06 
0.0 -1.4215 0 2.0 1e-06 
0.0 -1.4214 0 2.0 1e-06 
0.0 -1.4213 0 2.0 1e-06 
0.0 -1.4212 0 2.0 1e-06 
0.0 -1.4211 0 2.0 1e-06 
0.0 -1.421 0 2.0 1e-06 
0.0 -1.4209 0 2.0 1e-06 
0.0 -1.4208 0 2.0 1e-06 
0.0 -1.4207 0 2.0 1e-06 
0.0 -1.4206 0 2.0 1e-06 
0.0 -1.4205 0 2.0 1e-06 
0.0 -1.4204 0 2.0 1e-06 
0.0 -1.4203 0 2.0 1e-06 
0.0 -1.4202 0 2.0 1e-06 
0.0 -1.4201 0 2.0 1e-06 
0.0 -1.42 0 2.0 1e-06 
0.0 -1.4199 0 2.0 1e-06 
0.0 -1.4198 0 2.0 1e-06 
0.0 -1.4197 0 2.0 1e-06 
0.0 -1.4196 0 2.0 1e-06 
0.0 -1.4195 0 2.0 1e-06 
0.0 -1.4194 0 2.0 1e-06 
0.0 -1.4193 0 2.0 1e-06 
0.0 -1.4192 0 2.0 1e-06 
0.0 -1.4191 0 2.0 1e-06 
0.0 -1.419 0 2.0 1e-06 
0.0 -1.4189 0 2.0 1e-06 
0.0 -1.4188 0 2.0 1e-06 
0.0 -1.4187 0 2.0 1e-06 
0.0 -1.4186 0 2.0 1e-06 
0.0 -1.4185 0 2.0 1e-06 
0.0 -1.4184 0 2.0 1e-06 
0.0 -1.4183 0 2.0 1e-06 
0.0 -1.4182 0 2.0 1e-06 
0.0 -1.4181 0 2.0 1e-06 
0.0 -1.418 0 2.0 1e-06 
0.0 -1.4179 0 2.0 1e-06 
0.0 -1.4178 0 2.0 1e-06 
0.0 -1.4177 0 2.0 1e-06 
0.0 -1.4176 0 2.0 1e-06 
0.0 -1.4175 0 2.0 1e-06 
0.0 -1.4174 0 2.0 1e-06 
0.0 -1.4173 0 2.0 1e-06 
0.0 -1.4172 0 2.0 1e-06 
0.0 -1.4171 0 2.0 1e-06 
0.0 -1.417 0 2.0 1e-06 
0.0 -1.4169 0 2.0 1e-06 
0.0 -1.4168 0 2.0 1e-06 
0.0 -1.4167 0 2.0 1e-06 
0.0 -1.4166 0 2.0 1e-06 
0.0 -1.4165 0 2.0 1e-06 
0.0 -1.4164 0 2.0 1e-06 
0.0 -1.4163 0 2.0 1e-06 
0.0 -1.4162 0 2.0 1e-06 
0.0 -1.4161 0 2.0 1e-06 
0.0 -1.416 0 2.0 1e-06 
0.0 -1.4159 0 2.0 1e-06 
0.0 -1.4158 0 2.0 1e-06 
0.0 -1.4157 0 2.0 1e-06 
0.0 -1.4156 0 2.0 1e-06 
0.0 -1.4155 0 2.0 1e-06 
0.0 -1.4154 0 2.0 1e-06 
0.0 -1.4153 0 2.0 1e-06 
0.0 -1.4152 0 2.0 1e-06 
0.0 -1.4151 0 2.0 1e-06 
0.0 -1.415 0 2.0 1e-06 
0.0 -1.4149 0 2.0 1e-06 
0.0 -1.4148 0 2.0 1e-06 
0.0 -1.4147 0 2.0 1e-06 
0.0 -1.4146 0 2.0 1e-06 
0.0 -1.4145 0 2.0 1e-06 
0.0 -1.4144 0 2.0 1e-06 
0.0 -1.4143 0 2.0 1e-06 
0.0 -1.4142 0 2.0 1e-06 
0.0 -1.4141 0 2.0 1e-06 
0.0 -1.414 0 2.0 1e-06 
0.0 -1.4139 0 2.0 1e-06 
0.0 -1.4138 0 2.0 1e-06 
0.0 -1.4137 0 2.0 1e-06 
0.0 -1.4136 0 2.0 1e-06 
0.0 -1.4135 0 2.0 1e-06 
0.0 -1.4134 0 2.0 1e-06 
0.0 -1.4133 0 2.0 1e-06 
0.0 -1.4132 0 2.0 1e-06 
0.0 -1.4131 0 2.0 1e-06 
0.0 -1.413 0 2.0 1e-06 
0.0 -1.4129 0 2.0 1e-06 
0.0 -1.4128 0 2.0 1e-06 
0.0 -1.4127 0 2.0 1e-06 
0.0 -1.4126 0 2.0 1e-06 
0.0 -1.4125 0 2.0 1e-06 
0.0 -1.4124 0 2.0 1e-06 
0.0 -1.4123 0 2.0 1e-06 
0.0 -1.4122 0 2.0 1e-06 
0.0 -1.4121 0 2.0 1e-06 
0.0 -1.412 0 2.0 1e-06 
0.0 -1.4119 0 2.0 1e-06 
0.0 -1.4118 0 2.0 1e-06 
0.0 -1.4117 0 2.0 1e-06 
0.0 -1.4116 0 2.0 1e-06 
0.0 -1.4115 0 2.0 1e-06 
0.0 -1.4114 0 2.0 1e-06 
0.0 -1.4113 0 2.0 1e-06 
0.0 -1.4112 0 2.0 1e-06 
0.0 -1.4111 0 2.0 1e-06 
0.0 -1.411 0 2.0 1e-06 
0.0 -1.4109 0 2.0 1e-06 
0.0 -1.4108 0 2.0 1e-06 
0.0 -1.4107 0 2.0 1e-06 
0.0 -1.4106 0 2.0 1e-06 
0.0 -1.4105 0 2.0 1e-06 
0.0 -1.4104 0 2.0 1e-06 
0.0 -1.4103 0 2.0 1e-06 
0.0 -1.4102 0 2.0 1e-06 
0.0 -1.4101 0 2.0 1e-06 
0.0 -1.41 0 2.0 1e-06 
0.0 -1.4099 0 2.0 1e-06 
0.0 -1.4098 0 2.0 1e-06 
0.0 -1.4097 0 2.0 1e-06 
0.0 -1.4096 0 2.0 1e-06 
0.0 -1.4095 0 2.0 1e-06 
0.0 -1.4094 0 2.0 1e-06 
0.0 -1.4093 0 2.0 1e-06 
0.0 -1.4092 0 2.0 1e-06 
0.0 -1.4091 0 2.0 1e-06 
0.0 -1.409 0 2.0 1e-06 
0.0 -1.4089 0 2.0 1e-06 
0.0 -1.4088 0 2.0 1e-06 
0.0 -1.4087 0 2.0 1e-06 
0.0 -1.4086 0 2.0 1e-06 
0.0 -1.4085 0 2.0 1e-06 
0.0 -1.4084 0 2.0 1e-06 
0.0 -1.4083 0 2.0 1e-06 
0.0 -1.4082 0 2.0 1e-06 
0.0 -1.4081 0 2.0 1e-06 
0.0 -1.408 0 2.0 1e-06 
0.0 -1.4079 0 2.0 1e-06 
0.0 -1.4078 0 2.0 1e-06 
0.0 -1.4077 0 2.0 1e-06 
0.0 -1.4076 0 2.0 1e-06 
0.0 -1.4075 0 2.0 1e-06 
0.0 -1.4074 0 2.0 1e-06 
0.0 -1.4073 0 2.0 1e-06 
0.0 -1.4072 0 2.0 1e-06 
0.0 -1.4071 0 2.0 1e-06 
0.0 -1.407 0 2.0 1e-06 
0.0 -1.4069 0 2.0 1e-06 
0.0 -1.4068 0 2.0 1e-06 
0.0 -1.4067 0 2.0 1e-06 
0.0 -1.4066 0 2.0 1e-06 
0.0 -1.4065 0 2.0 1e-06 
0.0 -1.4064 0 2.0 1e-06 
0.0 -1.4063 0 2.0 1e-06 
0.0 -1.4062 0 2.0 1e-06 
0.0 -1.4061 0 2.0 1e-06 
0.0 -1.406 0 2.0 1e-06 
0.0 -1.4059 0 2.0 1e-06 
0.0 -1.4058 0 2.0 1e-06 
0.0 -1.4057 0 2.0 1e-06 
0.0 -1.4056 0 2.0 1e-06 
0.0 -1.4055 0 2.0 1e-06 
0.0 -1.4054 0 2.0 1e-06 
0.0 -1.4053 0 2.0 1e-06 
0.0 -1.4052 0 2.0 1e-06 
0.0 -1.4051 0 2.0 1e-06 
0.0 -1.405 0 2.0 1e-06 
0.0 -1.4049 0 2.0 1e-06 
0.0 -1.4048 0 2.0 1e-06 
0.0 -1.4047 0 2.0 1e-06 
0.0 -1.4046 0 2.0 1e-06 
0.0 -1.4045 0 2.0 1e-06 
0.0 -1.4044 0 2.0 1e-06 
0.0 -1.4043 0 2.0 1e-06 
0.0 -1.4042 0 2.0 1e-06 
0.0 -1.4041 0 2.0 1e-06 
0.0 -1.404 0 2.0 1e-06 
0.0 -1.4039 0 2.0 1e-06 
0.0 -1.4038 0 2.0 1e-06 
0.0 -1.4037 0 2.0 1e-06 
0.0 -1.4036 0 2.0 1e-06 
0.0 -1.4035 0 2.0 1e-06 
0.0 -1.4034 0 2.0 1e-06 
0.0 -1.4033 0 2.0 1e-06 
0.0 -1.4032 0 2.0 1e-06 
0.0 -1.4031 0 2.0 1e-06 
0.0 -1.403 0 2.0 1e-06 
0.0 -1.4029 0 2.0 1e-06 
0.0 -1.4028 0 2.0 1e-06 
0.0 -1.4027 0 2.0 1e-06 
0.0 -1.4026 0 2.0 1e-06 
0.0 -1.4025 0 2.0 1e-06 
0.0 -1.4024 0 2.0 1e-06 
0.0 -1.4023 0 2.0 1e-06 
0.0 -1.4022 0 2.0 1e-06 
0.0 -1.4021 0 2.0 1e-06 
0.0 -1.402 0 2.0 1e-06 
0.0 -1.4019 0 2.0 1e-06 
0.0 -1.4018 0 2.0 1e-06 
0.0 -1.4017 0 2.0 1e-06 
0.0 -1.4016 0 2.0 1e-06 
0.0 -1.4015 0 2.0 1e-06 
0.0 -1.4014 0 2.0 1e-06 
0.0 -1.4013 0 2.0 1e-06 
0.0 -1.4012 0 2.0 1e-06 
0.0 -1.4011 0 2.0 1e-06 
0.0 -1.401 0 2.0 1e-06 
0.0 -1.4009 0 2.0 1e-06 
0.0 -1.4008 0 2.0 1e-06 
0.0 -1.4007 0 2.0 1e-06 
0.0 -1.4006 0 2.0 1e-06 
0.0 -1.4005 0 2.0 1e-06 
0.0 -1.4004 0 2.0 1e-06 
0.0 -1.4003 0 2.0 1e-06 
0.0 -1.4002 0 2.0 1e-06 
0.0 -1.4001 0 2.0 1e-06 
0.0 -1.4 0 2.0 1e-06 
0.0 -1.3999 0 2.0 1e-06 
0.0 -1.3998 0 2.0 1e-06 
0.0 -1.3997 0 2.0 1e-06 
0.0 -1.3996 0 2.0 1e-06 
0.0 -1.3995 0 2.0 1e-06 
0.0 -1.3994 0 2.0 1e-06 
0.0 -1.3993 0 2.0 1e-06 
0.0 -1.3992 0 2.0 1e-06 
0.0 -1.3991 0 2.0 1e-06 
0.0 -1.399 0 2.0 1e-06 
0.0 -1.3989 0 2.0 1e-06 
0.0 -1.3988 0 2.0 1e-06 
0.0 -1.3987 0 2.0 1e-06 
0.0 -1.3986 0 2.0 1e-06 
0.0 -1.3985 0 2.0 1e-06 
0.0 -1.3984 0 2.0 1e-06 
0.0 -1.3983 0 2.0 1e-06 
0.0 -1.3982 0 2.0 1e-06 
0.0 -1.3981 0 2.0 1e-06 
0.0 -1.398 0 2.0 1e-06 
0.0 -1.3979 0 2.0 1e-06 
0.0 -1.3978 0 2.0 1e-06 
0.0 -1.3977 0 2.0 1e-06 
0.0 -1.3976 0 2.0 1e-06 
0.0 -1.3975 0 2.0 1e-06 
0.0 -1.3974 0 2.0 1e-06 
0.0 -1.3973 0 2.0 1e-06 
0.0 -1.3972 0 2.0 1e-06 
0.0 -1.3971 0 2.0 1e-06 
0.0 -1.397 0 2.0 1e-06 
0.0 -1.3969 0 2.0 1e-06 
0.0 -1.3968 0 2.0 1e-06 
0.0 -1.3967 0 2.0 1e-06 
0.0 -1.3966 0 2.0 1e-06 
0.0 -1.3965 0 2.0 1e-06 
0.0 -1.3964 0 2.0 1e-06 
0.0 -1.3963 0 2.0 1e-06 
0.0 -1.3962 0 2.0 1e-06 
0.0 -1.3961 0 2.0 1e-06 
0.0 -1.396 0 2.0 1e-06 
0.0 -1.3959 0 2.0 1e-06 
0.0 -1.3958 0 2.0 1e-06 
0.0 -1.3957 0 2.0 1e-06 
0.0 -1.3956 0 2.0 1e-06 
0.0 -1.3955 0 2.0 1e-06 
0.0 -1.3954 0 2.0 1e-06 
0.0 -1.3953 0 2.0 1e-06 
0.0 -1.3952 0 2.0 1e-06 
0.0 -1.3951 0 2.0 1e-06 
0.0 -1.395 0 2.0 1e-06 
0.0 -1.3949 0 2.0 1e-06 
0.0 -1.3948 0 2.0 1e-06 
0.0 -1.3947 0 2.0 1e-06 
0.0 -1.3946 0 2.0 1e-06 
0.0 -1.3945 0 2.0 1e-06 
0.0 -1.3944 0 2.0 1e-06 
0.0 -1.3943 0 2.0 1e-06 
0.0 -1.3942 0 2.0 1e-06 
0.0 -1.3941 0 2.0 1e-06 
0.0 -1.394 0 2.0 1e-06 
0.0 -1.3939 0 2.0 1e-06 
0.0 -1.3938 0 2.0 1e-06 
0.0 -1.3937 0 2.0 1e-06 
0.0 -1.3936 0 2.0 1e-06 
0.0 -1.3935 0 2.0 1e-06 
0.0 -1.3934 0 2.0 1e-06 
0.0 -1.3933 0 2.0 1e-06 
0.0 -1.3932 0 2.0 1e-06 
0.0 -1.3931 0 2.0 1e-06 
0.0 -1.393 0 2.0 1e-06 
0.0 -1.3929 0 2.0 1e-06 
0.0 -1.3928 0 2.0 1e-06 
0.0 -1.3927 0 2.0 1e-06 
0.0 -1.3926 0 2.0 1e-06 
0.0 -1.3925 0 2.0 1e-06 
0.0 -1.3924 0 2.0 1e-06 
0.0 -1.3923 0 2.0 1e-06 
0.0 -1.3922 0 2.0 1e-06 
0.0 -1.3921 0 2.0 1e-06 
0.0 -1.392 0 2.0 1e-06 
0.0 -1.3919 0 2.0 1e-06 
0.0 -1.3918 0 2.0 1e-06 
0.0 -1.3917 0 2.0 1e-06 
0.0 -1.3916 0 2.0 1e-06 
0.0 -1.3915 0 2.0 1e-06 
0.0 -1.3914 0 2.0 1e-06 
0.0 -1.3913 0 2.0 1e-06 
0.0 -1.3912 0 2.0 1e-06 
0.0 -1.3911 0 2.0 1e-06 
0.0 -1.391 0 2.0 1e-06 
0.0 -1.3909 0 2.0 1e-06 
0.0 -1.3908 0 2.0 1e-06 
0.0 -1.3907 0 2.0 1e-06 
0.0 -1.3906 0 2.0 1e-06 
0.0 -1.3905 0 2.0 1e-06 
0.0 -1.3904 0 2.0 1e-06 
0.0 -1.3903 0 2.0 1e-06 
0.0 -1.3902 0 2.0 1e-06 
0.0 -1.3901 0 2.0 1e-06 
0.0 -1.39 0 2.0 1e-06 
0.0 -1.3899 0 2.0 1e-06 
0.0 -1.3898 0 2.0 1e-06 
0.0 -1.3897 0 2.0 1e-06 
0.0 -1.3896 0 2.0 1e-06 
0.0 -1.3895 0 2.0 1e-06 
0.0 -1.3894 0 2.0 1e-06 
0.0 -1.3893 0 2.0 1e-06 
0.0 -1.3892 0 2.0 1e-06 
0.0 -1.3891 0 2.0 1e-06 
0.0 -1.389 0 2.0 1e-06 
0.0 -1.3889 0 2.0 1e-06 
0.0 -1.3888 0 2.0 1e-06 
0.0 -1.3887 0 2.0 1e-06 
0.0 -1.3886 0 2.0 1e-06 
0.0 -1.3885 0 2.0 1e-06 
0.0 -1.3884 0 2.0 1e-06 
0.0 -1.3883 0 2.0 1e-06 
0.0 -1.3882 0 2.0 1e-06 
0.0 -1.3881 0 2.0 1e-06 
0.0 -1.388 0 2.0 1e-06 
0.0 -1.3879 0 2.0 1e-06 
0.0 -1.3878 0 2.0 1e-06 
0.0 -1.3877 0 2.0 1e-06 
0.0 -1.3876 0 2.0 1e-06 
0.0 -1.3875 0 2.0 1e-06 
0.0 -1.3874 0 2.0 1e-06 
0.0 -1.3873 0 2.0 1e-06 
0.0 -1.3872 0 2.0 1e-06 
0.0 -1.3871 0 2.0 1e-06 
0.0 -1.387 0 2.0 1e-06 
0.0 -1.3869 0 2.0 1e-06 
0.0 -1.3868 0 2.0 1e-06 
0.0 -1.3867 0 2.0 1e-06 
0.0 -1.3866 0 2.0 1e-06 
0.0 -1.3865 0 2.0 1e-06 
0.0 -1.3864 0 2.0 1e-06 
0.0 -1.3863 0 2.0 1e-06 
0.0 -1.3862 0 2.0 1e-06 
0.0 -1.3861 0 2.0 1e-06 
0.0 -1.386 0 2.0 1e-06 
0.0 -1.3859 0 2.0 1e-06 
0.0 -1.3858 0 2.0 1e-06 
0.0 -1.3857 0 2.0 1e-06 
0.0 -1.3856 0 2.0 1e-06 
0.0 -1.3855 0 2.0 1e-06 
0.0 -1.3854 0 2.0 1e-06 
0.0 -1.3853 0 2.0 1e-06 
0.0 -1.3852 0 2.0 1e-06 
0.0 -1.3851 0 2.0 1e-06 
0.0 -1.385 0 2.0 1e-06 
0.0 -1.3849 0 2.0 1e-06 
0.0 -1.3848 0 2.0 1e-06 
0.0 -1.3847 0 2.0 1e-06 
0.0 -1.3846 0 2.0 1e-06 
0.0 -1.3845 0 2.0 1e-06 
0.0 -1.3844 0 2.0 1e-06 
0.0 -1.3843 0 2.0 1e-06 
0.0 -1.3842 0 2.0 1e-06 
0.0 -1.3841 0 2.0 1e-06 
0.0 -1.384 0 2.0 1e-06 
0.0 -1.3839 0 2.0 1e-06 
0.0 -1.3838 0 2.0 1e-06 
0.0 -1.3837 0 2.0 1e-06 
0.0 -1.3836 0 2.0 1e-06 
0.0 -1.3835 0 2.0 1e-06 
0.0 -1.3834 0 2.0 1e-06 
0.0 -1.3833 0 2.0 1e-06 
0.0 -1.3832 0 2.0 1e-06 
0.0 -1.3831 0 2.0 1e-06 
0.0 -1.383 0 2.0 1e-06 
0.0 -1.3829 0 2.0 1e-06 
0.0 -1.3828 0 2.0 1e-06 
0.0 -1.3827 0 2.0 1e-06 
0.0 -1.3826 0 2.0 1e-06 
0.0 -1.3825 0 2.0 1e-06 
0.0 -1.3824 0 2.0 1e-06 
0.0 -1.3823 0 2.0 1e-06 
0.0 -1.3822 0 2.0 1e-06 
0.0 -1.3821 0 2.0 1e-06 
0.0 -1.382 0 2.0 1e-06 
0.0 -1.3819 0 2.0 1e-06 
0.0 -1.3818 0 2.0 1e-06 
0.0 -1.3817 0 2.0 1e-06 
0.0 -1.3816 0 2.0 1e-06 
0.0 -1.3815 0 2.0 1e-06 
0.0 -1.3814 0 2.0 1e-06 
0.0 -1.3813 0 2.0 1e-06 
0.0 -1.3812 0 2.0 1e-06 
0.0 -1.3811 0 2.0 1e-06 
0.0 -1.381 0 2.0 1e-06 
0.0 -1.3809 0 2.0 1e-06 
0.0 -1.3808 0 2.0 1e-06 
0.0 -1.3807 0 2.0 1e-06 
0.0 -1.3806 0 2.0 1e-06 
0.0 -1.3805 0 2.0 1e-06 
0.0 -1.3804 0 2.0 1e-06 
0.0 -1.3803 0 2.0 1e-06 
0.0 -1.3802 0 2.0 1e-06 
0.0 -1.3801 0 2.0 1e-06 
0.0 -1.38 0 2.0 1e-06 
0.0 -1.3799 0 2.0 1e-06 
0.0 -1.3798 0 2.0 1e-06 
0.0 -1.3797 0 2.0 1e-06 
0.0 -1.3796 0 2.0 1e-06 
0.0 -1.3795 0 2.0 1e-06 
0.0 -1.3794 0 2.0 1e-06 
0.0 -1.3793 0 2.0 1e-06 
0.0 -1.3792 0 2.0 1e-06 
0.0 -1.3791 0 2.0 1e-06 
0.0 -1.379 0 2.0 1e-06 
0.0 -1.3789 0 2.0 1e-06 
0.0 -1.3788 0 2.0 1e-06 
0.0 -1.3787 0 2.0 1e-06 
0.0 -1.3786 0 2.0 1e-06 
0.0 -1.3785 0 2.0 1e-06 
0.0 -1.3784 0 2.0 1e-06 
0.0 -1.3783 0 2.0 1e-06 
0.0 -1.3782 0 2.0 1e-06 
0.0 -1.3781 0 2.0 1e-06 
0.0 -1.378 0 2.0 1e-06 
0.0 -1.3779 0 2.0 1e-06 
0.0 -1.3778 0 2.0 1e-06 
0.0 -1.3777 0 2.0 1e-06 
0.0 -1.3776 0 2.0 1e-06 
0.0 -1.3775 0 2.0 1e-06 
0.0 -1.3774 0 2.0 1e-06 
0.0 -1.3773 0 2.0 1e-06 
0.0 -1.3772 0 2.0 1e-06 
0.0 -1.3771 0 2.0 1e-06 
0.0 -1.377 0 2.0 1e-06 
0.0 -1.3769 0 2.0 1e-06 
0.0 -1.3768 0 2.0 1e-06 
0.0 -1.3767 0 2.0 1e-06 
0.0 -1.3766 0 2.0 1e-06 
0.0 -1.3765 0 2.0 1e-06 
0.0 -1.3764 0 2.0 1e-06 
0.0 -1.3763 0 2.0 1e-06 
0.0 -1.3762 0 2.0 1e-06 
0.0 -1.3761 0 2.0 1e-06 
0.0 -1.376 0 2.0 1e-06 
0.0 -1.3759 0 2.0 1e-06 
0.0 -1.3758 0 2.0 1e-06 
0.0 -1.3757 0 2.0 1e-06 
0.0 -1.3756 0 2.0 1e-06 
0.0 -1.3755 0 2.0 1e-06 
0.0 -1.3754 0 2.0 1e-06 
0.0 -1.3753 0 2.0 1e-06 
0.0 -1.3752 0 2.0 1e-06 
0.0 -1.3751 0 2.0 1e-06 
0.0 -1.375 0 2.0 1e-06 
0.0 -1.3749 0 2.0 1e-06 
0.0 -1.3748 0 2.0 1e-06 
0.0 -1.3747 0 2.0 1e-06 
0.0 -1.3746 0 2.0 1e-06 
0.0 -1.3745 0 2.0 1e-06 
0.0 -1.3744 0 2.0 1e-06 
0.0 -1.3743 0 2.0 1e-06 
0.0 -1.3742 0 2.0 1e-06 
0.0 -1.3741 0 2.0 1e-06 
0.0 -1.374 0 2.0 1e-06 
0.0 -1.3739 0 2.0 1e-06 
0.0 -1.3738 0 2.0 1e-06 
0.0 -1.3737 0 2.0 1e-06 
0.0 -1.3736 0 2.0 1e-06 
0.0 -1.3735 0 2.0 1e-06 
0.0 -1.3734 0 2.0 1e-06 
0.0 -1.3733 0 2.0 1e-06 
0.0 -1.3732 0 2.0 1e-06 
0.0 -1.3731 0 2.0 1e-06 
0.0 -1.373 0 2.0 1e-06 
0.0 -1.3729 0 2.0 1e-06 
0.0 -1.3728 0 2.0 1e-06 
0.0 -1.3727 0 2.0 1e-06 
0.0 -1.3726 0 2.0 1e-06 
0.0 -1.3725 0 2.0 1e-06 
0.0 -1.3724 0 2.0 1e-06 
0.0 -1.3723 0 2.0 1e-06 
0.0 -1.3722 0 2.0 1e-06 
0.0 -1.3721 0 2.0 1e-06 
0.0 -1.372 0 2.0 1e-06 
0.0 -1.3719 0 2.0 1e-06 
0.0 -1.3718 0 2.0 1e-06 
0.0 -1.3717 0 2.0 1e-06 
0.0 -1.3716 0 2.0 1e-06 
0.0 -1.3715 0 2.0 1e-06 
0.0 -1.3714 0 2.0 1e-06 
0.0 -1.3713 0 2.0 1e-06 
0.0 -1.3712 0 2.0 1e-06 
0.0 -1.3711 0 2.0 1e-06 
0.0 -1.371 0 2.0 1e-06 
0.0 -1.3709 0 2.0 1e-06 
0.0 -1.3708 0 2.0 1e-06 
0.0 -1.3707 0 2.0 1e-06 
0.0 -1.3706 0 2.0 1e-06 
0.0 -1.3705 0 2.0 1e-06 
0.0 -1.3704 0 2.0 1e-06 
0.0 -1.3703 0 2.0 1e-06 
0.0 -1.3702 0 2.0 1e-06 
0.0 -1.3701 0 2.0 1e-06 
0.0 -1.37 0 2.0 1e-06 
0.0 -1.3699 0 2.0 1e-06 
0.0 -1.3698 0 2.0 1e-06 
0.0 -1.3697 0 2.0 1e-06 
0.0 -1.3696 0 2.0 1e-06 
0.0 -1.3695 0 2.0 1e-06 
0.0 -1.3694 0 2.0 1e-06 
0.0 -1.3693 0 2.0 1e-06 
0.0 -1.3692 0 2.0 1e-06 
0.0 -1.3691 0 2.0 1e-06 
0.0 -1.369 0 2.0 1e-06 
0.0 -1.3689 0 2.0 1e-06 
0.0 -1.3688 0 2.0 1e-06 
0.0 -1.3687 0 2.0 1e-06 
0.0 -1.3686 0 2.0 1e-06 
0.0 -1.3685 0 2.0 1e-06 
0.0 -1.3684 0 2.0 1e-06 
0.0 -1.3683 0 2.0 1e-06 
0.0 -1.3682 0 2.0 1e-06 
0.0 -1.3681 0 2.0 1e-06 
0.0 -1.368 0 2.0 1e-06 
0.0 -1.3679 0 2.0 1e-06 
0.0 -1.3678 0 2.0 1e-06 
0.0 -1.3677 0 2.0 1e-06 
0.0 -1.3676 0 2.0 1e-06 
0.0 -1.3675 0 2.0 1e-06 
0.0 -1.3674 0 2.0 1e-06 
0.0 -1.3673 0 2.0 1e-06 
0.0 -1.3672 0 2.0 1e-06 
0.0 -1.3671 0 2.0 1e-06 
0.0 -1.367 0 2.0 1e-06 
0.0 -1.3669 0 2.0 1e-06 
0.0 -1.3668 0 2.0 1e-06 
0.0 -1.3667 0 2.0 1e-06 
0.0 -1.3666 0 2.0 1e-06 
0.0 -1.3665 0 2.0 1e-06 
0.0 -1.3664 0 2.0 1e-06 
0.0 -1.3663 0 2.0 1e-06 
0.0 -1.3662 0 2.0 1e-06 
0.0 -1.3661 0 2.0 1e-06 
0.0 -1.366 0 2.0 1e-06 
0.0 -1.3659 0 2.0 1e-06 
0.0 -1.3658 0 2.0 1e-06 
0.0 -1.3657 0 2.0 1e-06 
0.0 -1.3656 0 2.0 1e-06 
0.0 -1.3655 0 2.0 1e-06 
0.0 -1.3654 0 2.0 1e-06 
0.0 -1.3653 0 2.0 1e-06 
0.0 -1.3652 0 2.0 1e-06 
0.0 -1.3651 0 2.0 1e-06 
0.0 -1.365 0 2.0 1e-06 
0.0 -1.3649 0 2.0 1e-06 
0.0 -1.3648 0 2.0 1e-06 
0.0 -1.3647 0 2.0 1e-06 
0.0 -1.3646 0 2.0 1e-06 
0.0 -1.3645 0 2.0 1e-06 
0.0 -1.3644 0 2.0 1e-06 
0.0 -1.3643 0 2.0 1e-06 
0.0 -1.3642 0 2.0 1e-06 
0.0 -1.3641 0 2.0 1e-06 
0.0 -1.364 0 2.0 1e-06 
0.0 -1.3639 0 2.0 1e-06 
0.0 -1.3638 0 2.0 1e-06 
0.0 -1.3637 0 2.0 1e-06 
0.0 -1.3636 0 2.0 1e-06 
0.0 -1.3635 0 2.0 1e-06 
0.0 -1.3634 0 2.0 1e-06 
0.0 -1.3633 0 2.0 1e-06 
0.0 -1.3632 0 2.0 1e-06 
0.0 -1.3631 0 2.0 1e-06 
0.0 -1.363 0 2.0 1e-06 
0.0 -1.3629 0 2.0 1e-06 
0.0 -1.3628 0 2.0 1e-06 
0.0 -1.3627 0 2.0 1e-06 
0.0 -1.3626 0 2.0 1e-06 
0.0 -1.3625 0 2.0 1e-06 
0.0 -1.3624 0 2.0 1e-06 
0.0 -1.3623 0 2.0 1e-06 
0.0 -1.3622 0 2.0 1e-06 
0.0 -1.3621 0 2.0 1e-06 
0.0 -1.362 0 2.0 1e-06 
0.0 -1.3619 0 2.0 1e-06 
0.0 -1.3618 0 2.0 1e-06 
0.0 -1.3617 0 2.0 1e-06 
0.0 -1.3616 0 2.0 1e-06 
0.0 -1.3615 0 2.0 1e-06 
0.0 -1.3614 0 2.0 1e-06 
0.0 -1.3613 0 2.0 1e-06 
0.0 -1.3612 0 2.0 1e-06 
0.0 -1.3611 0 2.0 1e-06 
0.0 -1.361 0 2.0 1e-06 
0.0 -1.3609 0 2.0 1e-06 
0.0 -1.3608 0 2.0 1e-06 
0.0 -1.3607 0 2.0 1e-06 
0.0 -1.3606 0 2.0 1e-06 
0.0 -1.3605 0 2.0 1e-06 
0.0 -1.3604 0 2.0 1e-06 
0.0 -1.3603 0 2.0 1e-06 
0.0 -1.3602 0 2.0 1e-06 
0.0 -1.3601 0 2.0 1e-06 
0.0 -1.36 0 2.0 1e-06 
0.0 -1.3599 0 2.0 1e-06 
0.0 -1.3598 0 2.0 1e-06 
0.0 -1.3597 0 2.0 1e-06 
0.0 -1.3596 0 2.0 1e-06 
0.0 -1.3595 0 2.0 1e-06 
0.0 -1.3594 0 2.0 1e-06 
0.0 -1.3593 0 2.0 1e-06 
0.0 -1.3592 0 2.0 1e-06 
0.0 -1.3591 0 2.0 1e-06 
0.0 -1.359 0 2.0 1e-06 
0.0 -1.3589 0 2.0 1e-06 
0.0 -1.3588 0 2.0 1e-06 
0.0 -1.3587 0 2.0 1e-06 
0.0 -1.3586 0 2.0 1e-06 
0.0 -1.3585 0 2.0 1e-06 
0.0 -1.3584 0 2.0 1e-06 
0.0 -1.3583 0 2.0 1e-06 
0.0 -1.3582 0 2.0 1e-06 
0.0 -1.3581 0 2.0 1e-06 
0.0 -1.358 0 2.0 1e-06 
0.0 -1.3579 0 2.0 1e-06 
0.0 -1.3578 0 2.0 1e-06 
0.0 -1.3577 0 2.0 1e-06 
0.0 -1.3576 0 2.0 1e-06 
0.0 -1.3575 0 2.0 1e-06 
0.0 -1.3574 0 2.0 1e-06 
0.0 -1.3573 0 2.0 1e-06 
0.0 -1.3572 0 2.0 1e-06 
0.0 -1.3571 0 2.0 1e-06 
0.0 -1.357 0 2.0 1e-06 
0.0 -1.3569 0 2.0 1e-06 
0.0 -1.3568 0 2.0 1e-06 
0.0 -1.3567 0 2.0 1e-06 
0.0 -1.3566 0 2.0 1e-06 
0.0 -1.3565 0 2.0 1e-06 
0.0 -1.3564 0 2.0 1e-06 
0.0 -1.3563 0 2.0 1e-06 
0.0 -1.3562 0 2.0 1e-06 
0.0 -1.3561 0 2.0 1e-06 
0.0 -1.356 0 2.0 1e-06 
0.0 -1.3559 0 2.0 1e-06 
0.0 -1.3558 0 2.0 1e-06 
0.0 -1.3557 0 2.0 1e-06 
0.0 -1.3556 0 2.0 1e-06 
0.0 -1.3555 0 2.0 1e-06 
0.0 -1.3554 0 2.0 1e-06 
0.0 -1.3553 0 2.0 1e-06 
0.0 -1.3552 0 2.0 1e-06 
0.0 -1.3551 0 2.0 1e-06 
0.0 -1.355 0 2.0 1e-06 
0.0 -1.3549 0 2.0 1e-06 
0.0 -1.3548 0 2.0 1e-06 
0.0 -1.3547 0 2.0 1e-06 
0.0 -1.3546 0 2.0 1e-06 
0.0 -1.3545 0 2.0 1e-06 
0.0 -1.3544 0 2.0 1e-06 
0.0 -1.3543 0 2.0 1e-06 
0.0 -1.3542 0 2.0 1e-06 
0.0 -1.3541 0 2.0 1e-06 
0.0 -1.354 0 2.0 1e-06 
0.0 -1.3539 0 2.0 1e-06 
0.0 -1.3538 0 2.0 1e-06 
0.0 -1.3537 0 2.0 1e-06 
0.0 -1.3536 0 2.0 1e-06 
0.0 -1.3535 0 2.0 1e-06 
0.0 -1.3534 0 2.0 1e-06 
0.0 -1.3533 0 2.0 1e-06 
0.0 -1.3532 0 2.0 1e-06 
0.0 -1.3531 0 2.0 1e-06 
0.0 -1.353 0 2.0 1e-06 
0.0 -1.3529 0 2.0 1e-06 
0.0 -1.3528 0 2.0 1e-06 
0.0 -1.3527 0 2.0 1e-06 
0.0 -1.3526 0 2.0 1e-06 
0.0 -1.3525 0 2.0 1e-06 
0.0 -1.3524 0 2.0 1e-06 
0.0 -1.3523 0 2.0 1e-06 
0.0 -1.3522 0 2.0 1e-06 
0.0 -1.3521 0 2.0 1e-06 
0.0 -1.352 0 2.0 1e-06 
0.0 -1.3519 0 2.0 1e-06 
0.0 -1.3518 0 2.0 1e-06 
0.0 -1.3517 0 2.0 1e-06 
0.0 -1.3516 0 2.0 1e-06 
0.0 -1.3515 0 2.0 1e-06 
0.0 -1.3514 0 2.0 1e-06 
0.0 -1.3513 0 2.0 1e-06 
0.0 -1.3512 0 2.0 1e-06 
0.0 -1.3511 0 2.0 1e-06 
0.0 -1.351 0 2.0 1e-06 
0.0 -1.3509 0 2.0 1e-06 
0.0 -1.3508 0 2.0 1e-06 
0.0 -1.3507 0 2.0 1e-06 
0.0 -1.3506 0 2.0 1e-06 
0.0 -1.3505 0 2.0 1e-06 
0.0 -1.3504 0 2.0 1e-06 
0.0 -1.3503 0 2.0 1e-06 
0.0 -1.3502 0 2.0 1e-06 
0.0 -1.3501 0 2.0 1e-06 
0.0 -1.35 0 2.0 1e-06 
0.0 -1.3499 0 2.0 1e-06 
0.0 -1.3498 0 2.0 1e-06 
0.0 -1.3497 0 2.0 1e-06 
0.0 -1.3496 0 2.0 1e-06 
0.0 -1.3495 0 2.0 1e-06 
0.0 -1.3494 0 2.0 1e-06 
0.0 -1.3493 0 2.0 1e-06 
0.0 -1.3492 0 2.0 1e-06 
0.0 -1.3491 0 2.0 1e-06 
0.0 -1.349 0 2.0 1e-06 
0.0 -1.3489 0 2.0 1e-06 
0.0 -1.3488 0 2.0 1e-06 
0.0 -1.3487 0 2.0 1e-06 
0.0 -1.3486 0 2.0 1e-06 
0.0 -1.3485 0 2.0 1e-06 
0.0 -1.3484 0 2.0 1e-06 
0.0 -1.3483 0 2.0 1e-06 
0.0 -1.3482 0 2.0 1e-06 
0.0 -1.3481 0 2.0 1e-06 
0.0 -1.348 0 2.0 1e-06 
0.0 -1.3479 0 2.0 1e-06 
0.0 -1.3478 0 2.0 1e-06 
0.0 -1.3477 0 2.0 1e-06 
0.0 -1.3476 0 2.0 1e-06 
0.0 -1.3475 0 2.0 1e-06 
0.0 -1.3474 0 2.0 1e-06 
0.0 -1.3473 0 2.0 1e-06 
0.0 -1.3472 0 2.0 1e-06 
0.0 -1.3471 0 2.0 1e-06 
0.0 -1.347 0 2.0 1e-06 
0.0 -1.3469 0 2.0 1e-06 
0.0 -1.3468 0 2.0 1e-06 
0.0 -1.3467 0 2.0 1e-06 
0.0 -1.3466 0 2.0 1e-06 
0.0 -1.3465 0 2.0 1e-06 
0.0 -1.3464 0 2.0 1e-06 
0.0 -1.3463 0 2.0 1e-06 
0.0 -1.3462 0 2.0 1e-06 
0.0 -1.3461 0 2.0 1e-06 
0.0 -1.346 0 2.0 1e-06 
0.0 -1.3459 0 2.0 1e-06 
0.0 -1.3458 0 2.0 1e-06 
0.0 -1.3457 0 2.0 1e-06 
0.0 -1.3456 0 2.0 1e-06 
0.0 -1.3455 0 2.0 1e-06 
0.0 -1.3454 0 2.0 1e-06 
0.0 -1.3453 0 2.0 1e-06 
0.0 -1.3452 0 2.0 1e-06 
0.0 -1.3451 0 2.0 1e-06 
0.0 -1.345 0 2.0 1e-06 
0.0 -1.3449 0 2.0 1e-06 
0.0 -1.3448 0 2.0 1e-06 
0.0 -1.3447 0 2.0 1e-06 
0.0 -1.3446 0 2.0 1e-06 
0.0 -1.3445 0 2.0 1e-06 
0.0 -1.3444 0 2.0 1e-06 
0.0 -1.3443 0 2.0 1e-06 
0.0 -1.3442 0 2.0 1e-06 
0.0 -1.3441 0 2.0 1e-06 
0.0 -1.344 0 2.0 1e-06 
0.0 -1.3439 0 2.0 1e-06 
0.0 -1.3438 0 2.0 1e-06 
0.0 -1.3437 0 2.0 1e-06 
0.0 -1.3436 0 2.0 1e-06 
0.0 -1.3435 0 2.0 1e-06 
0.0 -1.3434 0 2.0 1e-06 
0.0 -1.3433 0 2.0 1e-06 
0.0 -1.3432 0 2.0 1e-06 
0.0 -1.3431 0 2.0 1e-06 
0.0 -1.343 0 2.0 1e-06 
0.0 -1.3429 0 2.0 1e-06 
0.0 -1.3428 0 2.0 1e-06 
0.0 -1.3427 0 2.0 1e-06 
0.0 -1.3426 0 2.0 1e-06 
0.0 -1.3425 0 2.0 1e-06 
0.0 -1.3424 0 2.0 1e-06 
0.0 -1.3423 0 2.0 1e-06 
0.0 -1.3422 0 2.0 1e-06 
0.0 -1.3421 0 2.0 1e-06 
0.0 -1.342 0 2.0 1e-06 
0.0 -1.3419 0 2.0 1e-06 
0.0 -1.3418 0 2.0 1e-06 
0.0 -1.3417 0 2.0 1e-06 
0.0 -1.3416 0 2.0 1e-06 
0.0 -1.3415 0 2.0 1e-06 
0.0 -1.3414 0 2.0 1e-06 
0.0 -1.3413 0 2.0 1e-06 
0.0 -1.3412 0 2.0 1e-06 
0.0 -1.3411 0 2.0 1e-06 
0.0 -1.341 0 2.0 1e-06 
0.0 -1.3409 0 2.0 1e-06 
0.0 -1.3408 0 2.0 1e-06 
0.0 -1.3407 0 2.0 1e-06 
0.0 -1.3406 0 2.0 1e-06 
0.0 -1.3405 0 2.0 1e-06 
0.0 -1.3404 0 2.0 1e-06 
0.0 -1.3403 0 2.0 1e-06 
0.0 -1.3402 0 2.0 1e-06 
0.0 -1.3401 0 2.0 1e-06 
0.0 -1.34 0 2.0 1e-06 
0.0 -1.3399 0 2.0 1e-06 
0.0 -1.3398 0 2.0 1e-06 
0.0 -1.3397 0 2.0 1e-06 
0.0 -1.3396 0 2.0 1e-06 
0.0 -1.3395 0 2.0 1e-06 
0.0 -1.3394 0 2.0 1e-06 
0.0 -1.3393 0 2.0 1e-06 
0.0 -1.3392 0 2.0 1e-06 
0.0 -1.3391 0 2.0 1e-06 
0.0 -1.339 0 2.0 1e-06 
0.0 -1.3389 0 2.0 1e-06 
0.0 -1.3388 0 2.0 1e-06 
0.0 -1.3387 0 2.0 1e-06 
0.0 -1.3386 0 2.0 1e-06 
0.0 -1.3385 0 2.0 1e-06 
0.0 -1.3384 0 2.0 1e-06 
0.0 -1.3383 0 2.0 1e-06 
0.0 -1.3382 0 2.0 1e-06 
0.0 -1.3381 0 2.0 1e-06 
0.0 -1.338 0 2.0 1e-06 
0.0 -1.3379 0 2.0 1e-06 
0.0 -1.3378 0 2.0 1e-06 
0.0 -1.3377 0 2.0 1e-06 
0.0 -1.3376 0 2.0 1e-06 
0.0 -1.3375 0 2.0 1e-06 
0.0 -1.3374 0 2.0 1e-06 
0.0 -1.3373 0 2.0 1e-06 
0.0 -1.3372 0 2.0 1e-06 
0.0 -1.3371 0 2.0 1e-06 
0.0 -1.337 0 2.0 1e-06 
0.0 -1.3369 0 2.0 1e-06 
0.0 -1.3368 0 2.0 1e-06 
0.0 -1.3367 0 2.0 1e-06 
0.0 -1.3366 0 2.0 1e-06 
0.0 -1.3365 0 2.0 1e-06 
0.0 -1.3364 0 2.0 1e-06 
0.0 -1.3363 0 2.0 1e-06 
0.0 -1.3362 0 2.0 1e-06 
0.0 -1.3361 0 2.0 1e-06 
0.0 -1.336 0 2.0 1e-06 
0.0 -1.3359 0 2.0 1e-06 
0.0 -1.3358 0 2.0 1e-06 
0.0 -1.3357 0 2.0 1e-06 
0.0 -1.3356 0 2.0 1e-06 
0.0 -1.3355 0 2.0 1e-06 
0.0 -1.3354 0 2.0 1e-06 
0.0 -1.3353 0 2.0 1e-06 
0.0 -1.3352 0 2.0 1e-06 
0.0 -1.3351 0 2.0 1e-06 
0.0 -1.335 0 2.0 1e-06 
0.0 -1.3349 0 2.0 1e-06 
0.0 -1.3348 0 2.0 1e-06 
0.0 -1.3347 0 2.0 1e-06 
0.0 -1.3346 0 2.0 1e-06 
0.0 -1.3345 0 2.0 1e-06 
0.0 -1.3344 0 2.0 1e-06 
0.0 -1.3343 0 2.0 1e-06 
0.0 -1.3342 0 2.0 1e-06 
0.0 -1.3341 0 2.0 1e-06 
0.0 -1.334 0 2.0 1e-06 
0.0 -1.3339 0 2.0 1e-06 
0.0 -1.3338 0 2.0 1e-06 
0.0 -1.3337 0 2.0 1e-06 
0.0 -1.3336 0 2.0 1e-06 
0.0 -1.3335 0 2.0 1e-06 
0.0 -1.3334 0 2.0 1e-06 
0.0 -1.3333 0 2.0 1e-06 
0.0 -1.3332 0 2.0 1e-06 
0.0 -1.3331 0 2.0 1e-06 
0.0 -1.333 0 2.0 1e-06 
0.0 -1.3329 0 2.0 1e-06 
0.0 -1.3328 0 2.0 1e-06 
0.0 -1.3327 0 2.0 1e-06 
0.0 -1.3326 0 2.0 1e-06 
0.0 -1.3325 0 2.0 1e-06 
0.0 -1.3324 0 2.0 1e-06 
0.0 -1.3323 0 2.0 1e-06 
0.0 -1.3322 0 2.0 1e-06 
0.0 -1.3321 0 2.0 1e-06 
0.0 -1.332 0 2.0 1e-06 
0.0 -1.3319 0 2.0 1e-06 
0.0 -1.3318 0 2.0 1e-06 
0.0 -1.3317 0 2.0 1e-06 
0.0 -1.3316 0 2.0 1e-06 
0.0 -1.3315 0 2.0 1e-06 
0.0 -1.3314 0 2.0 1e-06 
0.0 -1.3313 0 2.0 1e-06 
0.0 -1.3312 0 2.0 1e-06 
0.0 -1.3311 0 2.0 1e-06 
0.0 -1.331 0 2.0 1e-06 
0.0 -1.3309 0 2.0 1e-06 
0.0 -1.3308 0 2.0 1e-06 
0.0 -1.3307 0 2.0 1e-06 
0.0 -1.3306 0 2.0 1e-06 
0.0 -1.3305 0 2.0 1e-06 
0.0 -1.3304 0 2.0 1e-06 
0.0 -1.3303 0 2.0 1e-06 
0.0 -1.3302 0 2.0 1e-06 
0.0 -1.3301 0 2.0 1e-06 
0.0 -1.33 0 2.0 1e-06 
0.0 -1.3299 0 2.0 1e-06 
0.0 -1.3298 0 2.0 1e-06 
0.0 -1.3297 0 2.0 1e-06 
0.0 -1.3296 0 2.0 1e-06 
0.0 -1.3295 0 2.0 1e-06 
0.0 -1.3294 0 2.0 1e-06 
0.0 -1.3293 0 2.0 1e-06 
0.0 -1.3292 0 2.0 1e-06 
0.0 -1.3291 0 2.0 1e-06 
0.0 -1.329 0 2.0 1e-06 
0.0 -1.3289 0 2.0 1e-06 
0.0 -1.3288 0 2.0 1e-06 
0.0 -1.3287 0 2.0 1e-06 
0.0 -1.3286 0 2.0 1e-06 
0.0 -1.3285 0 2.0 1e-06 
0.0 -1.3284 0 2.0 1e-06 
0.0 -1.3283 0 2.0 1e-06 
0.0 -1.3282 0 2.0 1e-06 
0.0 -1.3281 0 2.0 1e-06 
0.0 -1.328 0 2.0 1e-06 
0.0 -1.3279 0 2.0 1e-06 
0.0 -1.3278 0 2.0 1e-06 
0.0 -1.3277 0 2.0 1e-06 
0.0 -1.3276 0 2.0 1e-06 
0.0 -1.3275 0 2.0 1e-06 
0.0 -1.3274 0 2.0 1e-06 
0.0 -1.3273 0 2.0 1e-06 
0.0 -1.3272 0 2.0 1e-06 
0.0 -1.3271 0 2.0 1e-06 
0.0 -1.327 0 2.0 1e-06 
0.0 -1.3269 0 2.0 1e-06 
0.0 -1.3268 0 2.0 1e-06 
0.0 -1.3267 0 2.0 1e-06 
0.0 -1.3266 0 2.0 1e-06 
0.0 -1.3265 0 2.0 1e-06 
0.0 -1.3264 0 2.0 1e-06 
0.0 -1.3263 0 2.0 1e-06 
0.0 -1.3262 0 2.0 1e-06 
0.0 -1.3261 0 2.0 1e-06 
0.0 -1.326 0 2.0 1e-06 
0.0 -1.3259 0 2.0 1e-06 
0.0 -1.3258 0 2.0 1e-06 
0.0 -1.3257 0 2.0 1e-06 
0.0 -1.3256 0 2.0 1e-06 
0.0 -1.3255 0 2.0 1e-06 
0.0 -1.3254 0 2.0 1e-06 
0.0 -1.3253 0 2.0 1e-06 
0.0 -1.3252 0 2.0 1e-06 
0.0 -1.3251 0 2.0 1e-06 
0.0 -1.325 0 2.0 1e-06 
0.0 -1.3249 0 2.0 1e-06 
0.0 -1.3248 0 2.0 1e-06 
0.0 -1.3247 0 2.0 1e-06 
0.0 -1.3246 0 2.0 1e-06 
0.0 -1.3245 0 2.0 1e-06 
0.0 -1.3244 0 2.0 1e-06 
0.0 -1.3243 0 2.0 1e-06 
0.0 -1.3242 0 2.0 1e-06 
0.0 -1.3241 0 2.0 1e-06 
0.0 -1.324 0 2.0 1e-06 
0.0 -1.3239 0 2.0 1e-06 
0.0 -1.3238 0 2.0 1e-06 
0.0 -1.3237 0 2.0 1e-06 
0.0 -1.3236 0 2.0 1e-06 
0.0 -1.3235 0 2.0 1e-06 
0.0 -1.3234 0 2.0 1e-06 
0.0 -1.3233 0 2.0 1e-06 
0.0 -1.3232 0 2.0 1e-06 
0.0 -1.3231 0 2.0 1e-06 
0.0 -1.323 0 2.0 1e-06 
0.0 -1.3229 0 2.0 1e-06 
0.0 -1.3228 0 2.0 1e-06 
0.0 -1.3227 0 2.0 1e-06 
0.0 -1.3226 0 2.0 1e-06 
0.0 -1.3225 0 2.0 1e-06 
0.0 -1.3224 0 2.0 1e-06 
0.0 -1.3223 0 2.0 1e-06 
0.0 -1.3222 0 2.0 1e-06 
0.0 -1.3221 0 2.0 1e-06 
0.0 -1.322 0 2.0 1e-06 
0.0 -1.3219 0 2.0 1e-06 
0.0 -1.3218 0 2.0 1e-06 
0.0 -1.3217 0 2.0 1e-06 
0.0 -1.3216 0 2.0 1e-06 
0.0 -1.3215 0 2.0 1e-06 
0.0 -1.3214 0 2.0 1e-06 
0.0 -1.3213 0 2.0 1e-06 
0.0 -1.3212 0 2.0 1e-06 
0.0 -1.3211 0 2.0 1e-06 
0.0 -1.321 0 2.0 1e-06 
0.0 -1.3209 0 2.0 1e-06 
0.0 -1.3208 0 2.0 1e-06 
0.0 -1.3207 0 2.0 1e-06 
0.0 -1.3206 0 2.0 1e-06 
0.0 -1.3205 0 2.0 1e-06 
0.0 -1.3204 0 2.0 1e-06 
0.0 -1.3203 0 2.0 1e-06 
0.0 -1.3202 0 2.0 1e-06 
0.0 -1.3201 0 2.0 1e-06 
0.0 -1.32 0 2.0 1e-06 
0.0 -1.3199 0 2.0 1e-06 
0.0 -1.3198 0 2.0 1e-06 
0.0 -1.3197 0 2.0 1e-06 
0.0 -1.3196 0 2.0 1e-06 
0.0 -1.3195 0 2.0 1e-06 
0.0 -1.3194 0 2.0 1e-06 
0.0 -1.3193 0 2.0 1e-06 
0.0 -1.3192 0 2.0 1e-06 
0.0 -1.3191 0 2.0 1e-06 
0.0 -1.319 0 2.0 1e-06 
0.0 -1.3189 0 2.0 1e-06 
0.0 -1.3188 0 2.0 1e-06 
0.0 -1.3187 0 2.0 1e-06 
0.0 -1.3186 0 2.0 1e-06 
0.0 -1.3185 0 2.0 1e-06 
0.0 -1.3184 0 2.0 1e-06 
0.0 -1.3183 0 2.0 1e-06 
0.0 -1.3182 0 2.0 1e-06 
0.0 -1.3181 0 2.0 1e-06 
0.0 -1.318 0 2.0 1e-06 
0.0 -1.3179 0 2.0 1e-06 
0.0 -1.3178 0 2.0 1e-06 
0.0 -1.3177 0 2.0 1e-06 
0.0 -1.3176 0 2.0 1e-06 
0.0 -1.3175 0 2.0 1e-06 
0.0 -1.3174 0 2.0 1e-06 
0.0 -1.3173 0 2.0 1e-06 
0.0 -1.3172 0 2.0 1e-06 
0.0 -1.3171 0 2.0 1e-06 
0.0 -1.317 0 2.0 1e-06 
0.0 -1.3169 0 2.0 1e-06 
0.0 -1.3168 0 2.0 1e-06 
0.0 -1.3167 0 2.0 1e-06 
0.0 -1.3166 0 2.0 1e-06 
0.0 -1.3165 0 2.0 1e-06 
0.0 -1.3164 0 2.0 1e-06 
0.0 -1.3163 0 2.0 1e-06 
0.0 -1.3162 0 2.0 1e-06 
0.0 -1.3161 0 2.0 1e-06 
0.0 -1.316 0 2.0 1e-06 
0.0 -1.3159 0 2.0 1e-06 
0.0 -1.3158 0 2.0 1e-06 
0.0 -1.3157 0 2.0 1e-06 
0.0 -1.3156 0 2.0 1e-06 
0.0 -1.3155 0 2.0 1e-06 
0.0 -1.3154 0 2.0 1e-06 
0.0 -1.3153 0 2.0 1e-06 
0.0 -1.3152 0 2.0 1e-06 
0.0 -1.3151 0 2.0 1e-06 
0.0 -1.315 0 2.0 1e-06 
0.0 -1.3149 0 2.0 1e-06 
0.0 -1.3148 0 2.0 1e-06 
0.0 -1.3147 0 2.0 1e-06 
0.0 -1.3146 0 2.0 1e-06 
0.0 -1.3145 0 2.0 1e-06 
0.0 -1.3144 0 2.0 1e-06 
0.0 -1.3143 0 2.0 1e-06 
0.0 -1.3142 0 2.0 1e-06 
0.0 -1.3141 0 2.0 1e-06 
0.0 -1.314 0 2.0 1e-06 
0.0 -1.3139 0 2.0 1e-06 
0.0 -1.3138 0 2.0 1e-06 
0.0 -1.3137 0 2.0 1e-06 
0.0 -1.3136 0 2.0 1e-06 
0.0 -1.3135 0 2.0 1e-06 
0.0 -1.3134 0 2.0 1e-06 
0.0 -1.3133 0 2.0 1e-06 
0.0 -1.3132 0 2.0 1e-06 
0.0 -1.3131 0 2.0 1e-06 
0.0 -1.313 0 2.0 1e-06 
0.0 -1.3129 0 2.0 1e-06 
0.0 -1.3128 0 2.0 1e-06 
0.0 -1.3127 0 2.0 1e-06 
0.0 -1.3126 0 2.0 1e-06 
0.0 -1.3125 0 2.0 1e-06 
0.0 -1.3124 0 2.0 1e-06 
0.0 -1.3123 0 2.0 1e-06 
0.0 -1.3122 0 2.0 1e-06 
0.0 -1.3121 0 2.0 1e-06 
0.0 -1.312 0 2.0 1e-06 
0.0 -1.3119 0 2.0 1e-06 
0.0 -1.3118 0 2.0 1e-06 
0.0 -1.3117 0 2.0 1e-06 
0.0 -1.3116 0 2.0 1e-06 
0.0 -1.3115 0 2.0 1e-06 
0.0 -1.3114 0 2.0 1e-06 
0.0 -1.3113 0 2.0 1e-06 
0.0 -1.3112 0 2.0 1e-06 
0.0 -1.3111 0 2.0 1e-06 
0.0 -1.311 0 2.0 1e-06 
0.0 -1.3109 0 2.0 1e-06 
0.0 -1.3108 0 2.0 1e-06 
0.0 -1.3107 0 2.0 1e-06 
0.0 -1.3106 0 2.0 1e-06 
0.0 -1.3105 0 2.0 1e-06 
0.0 -1.3104 0 2.0 1e-06 
0.0 -1.3103 0 2.0 1e-06 
0.0 -1.3102 0 2.0 1e-06 
0.0 -1.3101 0 2.0 1e-06 
0.0 -1.31 0 2.0 1e-06 
0.0 -1.3099 0 2.0 1e-06 
0.0 -1.3098 0 2.0 1e-06 
0.0 -1.3097 0 2.0 1e-06 
0.0 -1.3096 0 2.0 1e-06 
0.0 -1.3095 0 2.0 1e-06 
0.0 -1.3094 0 2.0 1e-06 
0.0 -1.3093 0 2.0 1e-06 
0.0 -1.3092 0 2.0 1e-06 
0.0 -1.3091 0 2.0 1e-06 
0.0 -1.309 0 2.0 1e-06 
0.0 -1.3089 0 2.0 1e-06 
0.0 -1.3088 0 2.0 1e-06 
0.0 -1.3087 0 2.0 1e-06 
0.0 -1.3086 0 2.0 1e-06 
0.0 -1.3085 0 2.0 1e-06 
0.0 -1.3084 0 2.0 1e-06 
0.0 -1.3083 0 2.0 1e-06 
0.0 -1.3082 0 2.0 1e-06 
0.0 -1.3081 0 2.0 1e-06 
0.0 -1.308 0 2.0 1e-06 
0.0 -1.3079 0 2.0 1e-06 
0.0 -1.3078 0 2.0 1e-06 
0.0 -1.3077 0 2.0 1e-06 
0.0 -1.3076 0 2.0 1e-06 
0.0 -1.3075 0 2.0 1e-06 
0.0 -1.3074 0 2.0 1e-06 
0.0 -1.3073 0 2.0 1e-06 
0.0 -1.3072 0 2.0 1e-06 
0.0 -1.3071 0 2.0 1e-06 
0.0 -1.307 0 2.0 1e-06 
0.0 -1.3069 0 2.0 1e-06 
0.0 -1.3068 0 2.0 1e-06 
0.0 -1.3067 0 2.0 1e-06 
0.0 -1.3066 0 2.0 1e-06 
0.0 -1.3065 0 2.0 1e-06 
0.0 -1.3064 0 2.0 1e-06 
0.0 -1.3063 0 2.0 1e-06 
0.0 -1.3062 0 2.0 1e-06 
0.0 -1.3061 0 2.0 1e-06 
0.0 -1.306 0 2.0 1e-06 
0.0 -1.3059 0 2.0 1e-06 
0.0 -1.3058 0 2.0 1e-06 
0.0 -1.3057 0 2.0 1e-06 
0.0 -1.3056 0 2.0 1e-06 
0.0 -1.3055 0 2.0 1e-06 
0.0 -1.3054 0 2.0 1e-06 
0.0 -1.3053 0 2.0 1e-06 
0.0 -1.3052 0 2.0 1e-06 
0.0 -1.3051 0 2.0 1e-06 
0.0 -1.305 0 2.0 1e-06 
0.0 -1.3049 0 2.0 1e-06 
0.0 -1.3048 0 2.0 1e-06 
0.0 -1.3047 0 2.0 1e-06 
0.0 -1.3046 0 2.0 1e-06 
0.0 -1.3045 0 2.0 1e-06 
0.0 -1.3044 0 2.0 1e-06 
0.0 -1.3043 0 2.0 1e-06 
0.0 -1.3042 0 2.0 1e-06 
0.0 -1.3041 0 2.0 1e-06 
0.0 -1.304 0 2.0 1e-06 
0.0 -1.3039 0 2.0 1e-06 
0.0 -1.3038 0 2.0 1e-06 
0.0 -1.3037 0 2.0 1e-06 
0.0 -1.3036 0 2.0 1e-06 
0.0 -1.3035 0 2.0 1e-06 
0.0 -1.3034 0 2.0 1e-06 
0.0 -1.3033 0 2.0 1e-06 
0.0 -1.3032 0 2.0 1e-06 
0.0 -1.3031 0 2.0 1e-06 
0.0 -1.303 0 2.0 1e-06 
0.0 -1.3029 0 2.0 1e-06 
0.0 -1.3028 0 2.0 1e-06 
0.0 -1.3027 0 2.0 1e-06 
0.0 -1.3026 0 2.0 1e-06 
0.0 -1.3025 0 2.0 1e-06 
0.0 -1.3024 0 2.0 1e-06 
0.0 -1.3023 0 2.0 1e-06 
0.0 -1.3022 0 2.0 1e-06 
0.0 -1.3021 0 2.0 1e-06 
0.0 -1.302 0 2.0 1e-06 
0.0 -1.3019 0 2.0 1e-06 
0.0 -1.3018 0 2.0 1e-06 
0.0 -1.3017 0 2.0 1e-06 
0.0 -1.3016 0 2.0 1e-06 
0.0 -1.3015 0 2.0 1e-06 
0.0 -1.3014 0 2.0 1e-06 
0.0 -1.3013 0 2.0 1e-06 
0.0 -1.3012 0 2.0 1e-06 
0.0 -1.3011 0 2.0 1e-06 
0.0 -1.301 0 2.0 1e-06 
0.0 -1.3009 0 2.0 1e-06 
0.0 -1.3008 0 2.0 1e-06 
0.0 -1.3007 0 2.0 1e-06 
0.0 -1.3006 0 2.0 1e-06 
0.0 -1.3005 0 2.0 1e-06 
0.0 -1.3004 0 2.0 1e-06 
0.0 -1.3003 0 2.0 1e-06 
0.0 -1.3002 0 2.0 1e-06 
0.0 -1.3001 0 2.0 1e-06 
0.0 -1.3 0 2.0 1e-06 
0.0 -1.2999 0 2.0 1e-06 
0.0 -1.2998 0 2.0 1e-06 
0.0 -1.2997 0 2.0 1e-06 
0.0 -1.2996 0 2.0 1e-06 
0.0 -1.2995 0 2.0 1e-06 
0.0 -1.2994 0 2.0 1e-06 
0.0 -1.2993 0 2.0 1e-06 
0.0 -1.2992 0 2.0 1e-06 
0.0 -1.2991 0 2.0 1e-06 
0.0 -1.299 0 2.0 1e-06 
0.0 -1.2989 0 2.0 1e-06 
0.0 -1.2988 0 2.0 1e-06 
0.0 -1.2987 0 2.0 1e-06 
0.0 -1.2986 0 2.0 1e-06 
0.0 -1.2985 0 2.0 1e-06 
0.0 -1.2984 0 2.0 1e-06 
0.0 -1.2983 0 2.0 1e-06 
0.0 -1.2982 0 2.0 1e-06 
0.0 -1.2981 0 2.0 1e-06 
0.0 -1.298 0 2.0 1e-06 
0.0 -1.2979 0 2.0 1e-06 
0.0 -1.2978 0 2.0 1e-06 
0.0 -1.2977 0 2.0 1e-06 
0.0 -1.2976 0 2.0 1e-06 
0.0 -1.2975 0 2.0 1e-06 
0.0 -1.2974 0 2.0 1e-06 
0.0 -1.2973 0 2.0 1e-06 
0.0 -1.2972 0 2.0 1e-06 
0.0 -1.2971 0 2.0 1e-06 
0.0 -1.297 0 2.0 1e-06 
0.0 -1.2969 0 2.0 1e-06 
0.0 -1.2968 0 2.0 1e-06 
0.0 -1.2967 0 2.0 1e-06 
0.0 -1.2966 0 2.0 1e-06 
0.0 -1.2965 0 2.0 1e-06 
0.0 -1.2964 0 2.0 1e-06 
0.0 -1.2963 0 2.0 1e-06 
0.0 -1.2962 0 2.0 1e-06 
0.0 -1.2961 0 2.0 1e-06 
0.0 -1.296 0 2.0 1e-06 
0.0 -1.2959 0 2.0 1e-06 
0.0 -1.2958 0 2.0 1e-06 
0.0 -1.2957 0 2.0 1e-06 
0.0 -1.2956 0 2.0 1e-06 
0.0 -1.2955 0 2.0 1e-06 
0.0 -1.2954 0 2.0 1e-06 
0.0 -1.2953 0 2.0 1e-06 
0.0 -1.2952 0 2.0 1e-06 
0.0 -1.2951 0 2.0 1e-06 
0.0 -1.295 0 2.0 1e-06 
0.0 -1.2949 0 2.0 1e-06 
0.0 -1.2948 0 2.0 1e-06 
0.0 -1.2947 0 2.0 1e-06 
0.0 -1.2946 0 2.0 1e-06 
0.0 -1.2945 0 2.0 1e-06 
0.0 -1.2944 0 2.0 1e-06 
0.0 -1.2943 0 2.0 1e-06 
0.0 -1.2942 0 2.0 1e-06 
0.0 -1.2941 0 2.0 1e-06 
0.0 -1.294 0 2.0 1e-06 
0.0 -1.2939 0 2.0 1e-06 
0.0 -1.2938 0 2.0 1e-06 
0.0 -1.2937 0 2.0 1e-06 
0.0 -1.2936 0 2.0 1e-06 
0.0 -1.2935 0 2.0 1e-06 
0.0 -1.2934 0 2.0 1e-06 
0.0 -1.2933 0 2.0 1e-06 
0.0 -1.2932 0 2.0 1e-06 
0.0 -1.2931 0 2.0 1e-06 
0.0 -1.293 0 2.0 1e-06 
0.0 -1.2929 0 2.0 1e-06 
0.0 -1.2928 0 2.0 1e-06 
0.0 -1.2927 0 2.0 1e-06 
0.0 -1.2926 0 2.0 1e-06 
0.0 -1.2925 0 2.0 1e-06 
0.0 -1.2924 0 2.0 1e-06 
0.0 -1.2923 0 2.0 1e-06 
0.0 -1.2922 0 2.0 1e-06 
0.0 -1.2921 0 2.0 1e-06 
0.0 -1.292 0 2.0 1e-06 
0.0 -1.2919 0 2.0 1e-06 
0.0 -1.2918 0 2.0 1e-06 
0.0 -1.2917 0 2.0 1e-06 
0.0 -1.2916 0 2.0 1e-06 
0.0 -1.2915 0 2.0 1e-06 
0.0 -1.2914 0 2.0 1e-06 
0.0 -1.2913 0 2.0 1e-06 
0.0 -1.2912 0 2.0 1e-06 
0.0 -1.2911 0 2.0 1e-06 
0.0 -1.291 0 2.0 1e-06 
0.0 -1.2909 0 2.0 1e-06 
0.0 -1.2908 0 2.0 1e-06 
0.0 -1.2907 0 2.0 1e-06 
0.0 -1.2906 0 2.0 1e-06 
0.0 -1.2905 0 2.0 1e-06 
0.0 -1.2904 0 2.0 1e-06 
0.0 -1.2903 0 2.0 1e-06 
0.0 -1.2902 0 2.0 1e-06 
0.0 -1.2901 0 2.0 1e-06 
0.0 -1.29 0 2.0 1e-06 
0.0 -1.2899 0 2.0 1e-06 
0.0 -1.2898 0 2.0 1e-06 
0.0 -1.2897 0 2.0 1e-06 
0.0 -1.2896 0 2.0 1e-06 
0.0 -1.2895 0 2.0 1e-06 
0.0 -1.2894 0 2.0 1e-06 
0.0 -1.2893 0 2.0 1e-06 
0.0 -1.2892 0 2.0 1e-06 
0.0 -1.2891 0 2.0 1e-06 
0.0 -1.289 0 2.0 1e-06 
0.0 -1.2889 0 2.0 1e-06 
0.0 -1.2888 0 2.0 1e-06 
0.0 -1.2887 0 2.0 1e-06 
0.0 -1.2886 0 2.0 1e-06 
0.0 -1.2885 0 2.0 1e-06 
0.0 -1.2884 0 2.0 1e-06 
0.0 -1.2883 0 2.0 1e-06 
0.0 -1.2882 0 2.0 1e-06 
0.0 -1.2881 0 2.0 1e-06 
0.0 -1.288 0 2.0 1e-06 
0.0 -1.2879 0 2.0 1e-06 
0.0 -1.2878 0 2.0 1e-06 
0.0 -1.2877 0 2.0 1e-06 
0.0 -1.2876 0 2.0 1e-06 
0.0 -1.2875 0 2.0 1e-06 
0.0 -1.2874 0 2.0 1e-06 
0.0 -1.2873 0 2.0 1e-06 
0.0 -1.2872 0 2.0 1e-06 
0.0 -1.2871 0 2.0 1e-06 
0.0 -1.287 0 2.0 1e-06 
0.0 -1.2869 0 2.0 1e-06 
0.0 -1.2868 0 2.0 1e-06 
0.0 -1.2867 0 2.0 1e-06 
0.0 -1.2866 0 2.0 1e-06 
0.0 -1.2865 0 2.0 1e-06 
0.0 -1.2864 0 2.0 1e-06 
0.0 -1.2863 0 2.0 1e-06 
0.0 -1.2862 0 2.0 1e-06 
0.0 -1.2861 0 2.0 1e-06 
0.0 -1.286 0 2.0 1e-06 
0.0 -1.2859 0 2.0 1e-06 
0.0 -1.2858 0 2.0 1e-06 
0.0 -1.2857 0 2.0 1e-06 
0.0 -1.2856 0 2.0 1e-06 
0.0 -1.2855 0 2.0 1e-06 
0.0 -1.2854 0 2.0 1e-06 
0.0 -1.2853 0 2.0 1e-06 
0.0 -1.2852 0 2.0 1e-06 
0.0 -1.2851 0 2.0 1e-06 
0.0 -1.285 0 2.0 1e-06 
0.0 -1.2849 0 2.0 1e-06 
0.0 -1.2848 0 2.0 1e-06 
0.0 -1.2847 0 2.0 1e-06 
0.0 -1.2846 0 2.0 1e-06 
0.0 -1.2845 0 2.0 1e-06 
0.0 -1.2844 0 2.0 1e-06 
0.0 -1.2843 0 2.0 1e-06 
0.0 -1.2842 0 2.0 1e-06 
0.0 -1.2841 0 2.0 1e-06 
0.0 -1.284 0 2.0 1e-06 
0.0 -1.2839 0 2.0 1e-06 
0.0 -1.2838 0 2.0 1e-06 
0.0 -1.2837 0 2.0 1e-06 
0.0 -1.2836 0 2.0 1e-06 
0.0 -1.2835 0 2.0 1e-06 
0.0 -1.2834 0 2.0 1e-06 
0.0 -1.2833 0 2.0 1e-06 
0.0 -1.2832 0 2.0 1e-06 
0.0 -1.2831 0 2.0 1e-06 
0.0 -1.283 0 2.0 1e-06 
0.0 -1.2829 0 2.0 1e-06 
0.0 -1.2828 0 2.0 1e-06 
0.0 -1.2827 0 2.0 1e-06 
0.0 -1.2826 0 2.0 1e-06 
0.0 -1.2825 0 2.0 1e-06 
0.0 -1.2824 0 2.0 1e-06 
0.0 -1.2823 0 2.0 1e-06 
0.0 -1.2822 0 2.0 1e-06 
0.0 -1.2821 0 2.0 1e-06 
0.0 -1.282 0 2.0 1e-06 
0.0 -1.2819 0 2.0 1e-06 
0.0 -1.2818 0 2.0 1e-06 
0.0 -1.2817 0 2.0 1e-06 
0.0 -1.2816 0 2.0 1e-06 
0.0 -1.2815 0 2.0 1e-06 
0.0 -1.2814 0 2.0 1e-06 
0.0 -1.2813 0 2.0 1e-06 
0.0 -1.2812 0 2.0 1e-06 
0.0 -1.2811 0 2.0 1e-06 
0.0 -1.281 0 2.0 1e-06 
0.0 -1.2809 0 2.0 1e-06 
0.0 -1.2808 0 2.0 1e-06 
0.0 -1.2807 0 2.0 1e-06 
0.0 -1.2806 0 2.0 1e-06 
0.0 -1.2805 0 2.0 1e-06 
0.0 -1.2804 0 2.0 1e-06 
0.0 -1.2803 0 2.0 1e-06 
0.0 -1.2802 0 2.0 1e-06 
0.0 -1.2801 0 2.0 1e-06 
0.0 -1.28 0 2.0 1e-06 
0.0 -1.2799 0 2.0 1e-06 
0.0 -1.2798 0 2.0 1e-06 
0.0 -1.2797 0 2.0 1e-06 
0.0 -1.2796 0 2.0 1e-06 
0.0 -1.2795 0 2.0 1e-06 
0.0 -1.2794 0 2.0 1e-06 
0.0 -1.2793 0 2.0 1e-06 
0.0 -1.2792 0 2.0 1e-06 
0.0 -1.2791 0 2.0 1e-06 
0.0 -1.279 0 2.0 1e-06 
0.0 -1.2789 0 2.0 1e-06 
0.0 -1.2788 0 2.0 1e-06 
0.0 -1.2787 0 2.0 1e-06 
0.0 -1.2786 0 2.0 1e-06 
0.0 -1.2785 0 2.0 1e-06 
0.0 -1.2784 0 2.0 1e-06 
0.0 -1.2783 0 2.0 1e-06 
0.0 -1.2782 0 2.0 1e-06 
0.0 -1.2781 0 2.0 1e-06 
0.0 -1.278 0 2.0 1e-06 
0.0 -1.2779 0 2.0 1e-06 
0.0 -1.2778 0 2.0 1e-06 
0.0 -1.2777 0 2.0 1e-06 
0.0 -1.2776 0 2.0 1e-06 
0.0 -1.2775 0 2.0 1e-06 
0.0 -1.2774 0 2.0 1e-06 
0.0 -1.2773 0 2.0 1e-06 
0.0 -1.2772 0 2.0 1e-06 
0.0 -1.2771 0 2.0 1e-06 
0.0 -1.277 0 2.0 1e-06 
0.0 -1.2769 0 2.0 1e-06 
0.0 -1.2768 0 2.0 1e-06 
0.0 -1.2767 0 2.0 1e-06 
0.0 -1.2766 0 2.0 1e-06 
0.0 -1.2765 0 2.0 1e-06 
0.0 -1.2764 0 2.0 1e-06 
0.0 -1.2763 0 2.0 1e-06 
0.0 -1.2762 0 2.0 1e-06 
0.0 -1.2761 0 2.0 1e-06 
0.0 -1.276 0 2.0 1e-06 
0.0 -1.2759 0 2.0 1e-06 
0.0 -1.2758 0 2.0 1e-06 
0.0 -1.2757 0 2.0 1e-06 
0.0 -1.2756 0 2.0 1e-06 
0.0 -1.2755 0 2.0 1e-06 
0.0 -1.2754 0 2.0 1e-06 
0.0 -1.2753 0 2.0 1e-06 
0.0 -1.2752 0 2.0 1e-06 
0.0 -1.2751 0 2.0 1e-06 
0.0 -1.275 0 2.0 1e-06 
0.0 -1.2749 0 2.0 1e-06 
0.0 -1.2748 0 2.0 1e-06 
0.0 -1.2747 0 2.0 1e-06 
0.0 -1.2746 0 2.0 1e-06 
0.0 -1.2745 0 2.0 1e-06 
0.0 -1.2744 0 2.0 1e-06 
0.0 -1.2743 0 2.0 1e-06 
0.0 -1.2742 0 2.0 1e-06 
0.0 -1.2741 0 2.0 1e-06 
0.0 -1.274 0 2.0 1e-06 
0.0 -1.2739 0 2.0 1e-06 
0.0 -1.2738 0 2.0 1e-06 
0.0 -1.2737 0 2.0 1e-06 
0.0 -1.2736 0 2.0 1e-06 
0.0 -1.2735 0 2.0 1e-06 
0.0 -1.2734 0 2.0 1e-06 
0.0 -1.2733 0 2.0 1e-06 
0.0 -1.2732 0 2.0 1e-06 
0.0 -1.2731 0 2.0 1e-06 
0.0 -1.273 0 2.0 1e-06 
0.0 -1.2729 0 2.0 1e-06 
0.0 -1.2728 0 2.0 1e-06 
0.0 -1.2727 0 2.0 1e-06 
0.0 -1.2726 0 2.0 1e-06 
0.0 -1.2725 0 2.0 1e-06 
0.0 -1.2724 0 2.0 1e-06 
0.0 -1.2723 0 2.0 1e-06 
0.0 -1.2722 0 2.0 1e-06 
0.0 -1.2721 0 2.0 1e-06 
0.0 -1.272 0 2.0 1e-06 
0.0 -1.2719 0 2.0 1e-06 
0.0 -1.2718 0 2.0 1e-06 
0.0 -1.2717 0 2.0 1e-06 
0.0 -1.2716 0 2.0 1e-06 
0.0 -1.2715 0 2.0 1e-06 
0.0 -1.2714 0 2.0 1e-06 
0.0 -1.2713 0 2.0 1e-06 
0.0 -1.2712 0 2.0 1e-06 
0.0 -1.2711 0 2.0 1e-06 
0.0 -1.271 0 2.0 1e-06 
0.0 -1.2709 0 2.0 1e-06 
0.0 -1.2708 0 2.0 1e-06 
0.0 -1.2707 0 2.0 1e-06 
0.0 -1.2706 0 2.0 1e-06 
0.0 -1.2705 0 2.0 1e-06 
0.0 -1.2704 0 2.0 1e-06 
0.0 -1.2703 0 2.0 1e-06 
0.0 -1.2702 0 2.0 1e-06 
0.0 -1.2701 0 2.0 1e-06 
0.0 -1.27 0 2.0 1e-06 
0.0 -1.2699 0 2.0 1e-06 
0.0 -1.2698 0 2.0 1e-06 
0.0 -1.2697 0 2.0 1e-06 
0.0 -1.2696 0 2.0 1e-06 
0.0 -1.2695 0 2.0 1e-06 
0.0 -1.2694 0 2.0 1e-06 
0.0 -1.2693 0 2.0 1e-06 
0.0 -1.2692 0 2.0 1e-06 
0.0 -1.2691 0 2.0 1e-06 
0.0 -1.269 0 2.0 1e-06 
0.0 -1.2689 0 2.0 1e-06 
0.0 -1.2688 0 2.0 1e-06 
0.0 -1.2687 0 2.0 1e-06 
0.0 -1.2686 0 2.0 1e-06 
0.0 -1.2685 0 2.0 1e-06 
0.0 -1.2684 0 2.0 1e-06 
0.0 -1.2683 0 2.0 1e-06 
0.0 -1.2682 0 2.0 1e-06 
0.0 -1.2681 0 2.0 1e-06 
0.0 -1.268 0 2.0 1e-06 
0.0 -1.2679 0 2.0 1e-06 
0.0 -1.2678 0 2.0 1e-06 
0.0 -1.2677 0 2.0 1e-06 
0.0 -1.2676 0 2.0 1e-06 
0.0 -1.2675 0 2.0 1e-06 
0.0 -1.2674 0 2.0 1e-06 
0.0 -1.2673 0 2.0 1e-06 
0.0 -1.2672 0 2.0 1e-06 
0.0 -1.2671 0 2.0 1e-06 
0.0 -1.267 0 2.0 1e-06 
0.0 -1.2669 0 2.0 1e-06 
0.0 -1.2668 0 2.0 1e-06 
0.0 -1.2667 0 2.0 1e-06 
0.0 -1.2666 0 2.0 1e-06 
0.0 -1.2665 0 2.0 1e-06 
0.0 -1.2664 0 2.0 1e-06 
0.0 -1.2663 0 2.0 1e-06 
0.0 -1.2662 0 2.0 1e-06 
0.0 -1.2661 0 2.0 1e-06 
0.0 -1.266 0 2.0 1e-06 
0.0 -1.2659 0 2.0 1e-06 
0.0 -1.2658 0 2.0 1e-06 
0.0 -1.2657 0 2.0 1e-06 
0.0 -1.2656 0 2.0 1e-06 
0.0 -1.2655 0 2.0 1e-06 
0.0 -1.2654 0 2.0 1e-06 
0.0 -1.2653 0 2.0 1e-06 
0.0 -1.2652 0 2.0 1e-06 
0.0 -1.2651 0 2.0 1e-06 
0.0 -1.265 0 2.0 1e-06 
0.0 -1.2649 0 2.0 1e-06 
0.0 -1.2648 0 2.0 1e-06 
0.0 -1.2647 0 2.0 1e-06 
0.0 -1.2646 0 2.0 1e-06 
0.0 -1.2645 0 2.0 1e-06 
0.0 -1.2644 0 2.0 1e-06 
0.0 -1.2643 0 2.0 1e-06 
0.0 -1.2642 0 2.0 1e-06 
0.0 -1.2641 0 2.0 1e-06 
0.0 -1.264 0 2.0 1e-06 
0.0 -1.2639 0 2.0 1e-06 
0.0 -1.2638 0 2.0 1e-06 
0.0 -1.2637 0 2.0 1e-06 
0.0 -1.2636 0 2.0 1e-06 
0.0 -1.2635 0 2.0 1e-06 
0.0 -1.2634 0 2.0 1e-06 
0.0 -1.2633 0 2.0 1e-06 
0.0 -1.2632 0 2.0 1e-06 
0.0 -1.2631 0 2.0 1e-06 
0.0 -1.263 0 2.0 1e-06 
0.0 -1.2629 0 2.0 1e-06 
0.0 -1.2628 0 2.0 1e-06 
0.0 -1.2627 0 2.0 1e-06 
0.0 -1.2626 0 2.0 1e-06 
0.0 -1.2625 0 2.0 1e-06 
0.0 -1.2624 0 2.0 1e-06 
0.0 -1.2623 0 2.0 1e-06 
0.0 -1.2622 0 2.0 1e-06 
0.0 -1.2621 0 2.0 1e-06 
0.0 -1.262 0 2.0 1e-06 
0.0 -1.2619 0 2.0 1e-06 
0.0 -1.2618 0 2.0 1e-06 
0.0 -1.2617 0 2.0 1e-06 
0.0 -1.2616 0 2.0 1e-06 
0.0 -1.2615 0 2.0 1e-06 
0.0 -1.2614 0 2.0 1e-06 
0.0 -1.2613 0 2.0 1e-06 
0.0 -1.2612 0 2.0 1e-06 
0.0 -1.2611 0 2.0 1e-06 
0.0 -1.261 0 2.0 1e-06 
0.0 -1.2609 0 2.0 1e-06 
0.0 -1.2608 0 2.0 1e-06 
0.0 -1.2607 0 2.0 1e-06 
0.0 -1.2606 0 2.0 1e-06 
0.0 -1.2605 0 2.0 1e-06 
0.0 -1.2604 0 2.0 1e-06 
0.0 -1.2603 0 2.0 1e-06 
0.0 -1.2602 0 2.0 1e-06 
0.0 -1.2601 0 2.0 1e-06 
0.0 -1.26 0 2.0 1e-06 
0.0 -1.2599 0 2.0 1e-06 
0.0 -1.2598 0 2.0 1e-06 
0.0 -1.2597 0 2.0 1e-06 
0.0 -1.2596 0 2.0 1e-06 
0.0 -1.2595 0 2.0 1e-06 
0.0 -1.2594 0 2.0 1e-06 
0.0 -1.2593 0 2.0 1e-06 
0.0 -1.2592 0 2.0 1e-06 
0.0 -1.2591 0 2.0 1e-06 
0.0 -1.259 0 2.0 1e-06 
0.0 -1.2589 0 2.0 1e-06 
0.0 -1.2588 0 2.0 1e-06 
0.0 -1.2587 0 2.0 1e-06 
0.0 -1.2586 0 2.0 1e-06 
0.0 -1.2585 0 2.0 1e-06 
0.0 -1.2584 0 2.0 1e-06 
0.0 -1.2583 0 2.0 1e-06 
0.0 -1.2582 0 2.0 1e-06 
0.0 -1.2581 0 2.0 1e-06 
0.0 -1.258 0 2.0 1e-06 
0.0 -1.2579 0 2.0 1e-06 
0.0 -1.2578 0 2.0 1e-06 
0.0 -1.2577 0 2.0 1e-06 
0.0 -1.2576 0 2.0 1e-06 
0.0 -1.2575 0 2.0 1e-06 
0.0 -1.2574 0 2.0 1e-06 
0.0 -1.2573 0 2.0 1e-06 
0.0 -1.2572 0 2.0 1e-06 
0.0 -1.2571 0 2.0 1e-06 
0.0 -1.257 0 2.0 1e-06 
0.0 -1.2569 0 2.0 1e-06 
0.0 -1.2568 0 2.0 1e-06 
0.0 -1.2567 0 2.0 1e-06 
0.0 -1.2566 0 2.0 1e-06 
0.0 -1.2565 0 2.0 1e-06 
0.0 -1.2564 0 2.0 1e-06 
0.0 -1.2563 0 2.0 1e-06 
0.0 -1.2562 0 2.0 1e-06 
0.0 -1.2561 0 2.0 1e-06 
0.0 -1.256 0 2.0 1e-06 
0.0 -1.2559 0 2.0 1e-06 
0.0 -1.2558 0 2.0 1e-06 
0.0 -1.2557 0 2.0 1e-06 
0.0 -1.2556 0 2.0 1e-06 
0.0 -1.2555 0 2.0 1e-06 
0.0 -1.2554 0 2.0 1e-06 
0.0 -1.2553 0 2.0 1e-06 
0.0 -1.2552 0 2.0 1e-06 
0.0 -1.2551 0 2.0 1e-06 
0.0 -1.255 0 2.0 1e-06 
0.0 -1.2549 0 2.0 1e-06 
0.0 -1.2548 0 2.0 1e-06 
0.0 -1.2547 0 2.0 1e-06 
0.0 -1.2546 0 2.0 1e-06 
0.0 -1.2545 0 2.0 1e-06 
0.0 -1.2544 0 2.0 1e-06 
0.0 -1.2543 0 2.0 1e-06 
0.0 -1.2542 0 2.0 1e-06 
0.0 -1.2541 0 2.0 1e-06 
0.0 -1.254 0 2.0 1e-06 
0.0 -1.2539 0 2.0 1e-06 
0.0 -1.2538 0 2.0 1e-06 
0.0 -1.2537 0 2.0 1e-06 
0.0 -1.2536 0 2.0 1e-06 
0.0 -1.2535 0 2.0 1e-06 
0.0 -1.2534 0 2.0 1e-06 
0.0 -1.2533 0 2.0 1e-06 
0.0 -1.2532 0 2.0 1e-06 
0.0 -1.2531 0 2.0 1e-06 
0.0 -1.253 0 2.0 1e-06 
0.0 -1.2529 0 2.0 1e-06 
0.0 -1.2528 0 2.0 1e-06 
0.0 -1.2527 0 2.0 1e-06 
0.0 -1.2526 0 2.0 1e-06 
0.0 -1.2525 0 2.0 1e-06 
0.0 -1.2524 0 2.0 1e-06 
0.0 -1.2523 0 2.0 1e-06 
0.0 -1.2522 0 2.0 1e-06 
0.0 -1.2521 0 2.0 1e-06 
0.0 -1.252 0 2.0 1e-06 
0.0 -1.2519 0 2.0 1e-06 
0.0 -1.2518 0 2.0 1e-06 
0.0 -1.2517 0 2.0 1e-06 
0.0 -1.2516 0 2.0 1e-06 
0.0 -1.2515 0 2.0 1e-06 
0.0 -1.2514 0 2.0 1e-06 
0.0 -1.2513 0 2.0 1e-06 
0.0 -1.2512 0 2.0 1e-06 
0.0 -1.2511 0 2.0 1e-06 
0.0 -1.251 0 2.0 1e-06 
0.0 -1.2509 0 2.0 1e-06 
0.0 -1.2508 0 2.0 1e-06 
0.0 -1.2507 0 2.0 1e-06 
0.0 -1.2506 0 2.0 1e-06 
0.0 -1.2505 0 2.0 1e-06 
0.0 -1.2504 0 2.0 1e-06 
0.0 -1.2503 0 2.0 1e-06 
0.0 -1.2502 0 2.0 1e-06 
0.0 -1.2501 0 2.0 1e-06 
0.0 -1.25 0 2.0 1e-06 
0.0 -1.2499 0 2.0 1e-06 
0.0 -1.2498 0 2.0 1e-06 
0.0 -1.2497 0 2.0 1e-06 
0.0 -1.2496 0 2.0 1e-06 
0.0 -1.2495 0 2.0 1e-06 
0.0 -1.2494 0 2.0 1e-06 
0.0 -1.2493 0 2.0 1e-06 
0.0 -1.2492 0 2.0 1e-06 
0.0 -1.2491 0 2.0 1e-06 
0.0 -1.249 0 2.0 1e-06 
0.0 -1.2489 0 2.0 1e-06 
0.0 -1.2488 0 2.0 1e-06 
0.0 -1.2487 0 2.0 1e-06 
0.0 -1.2486 0 2.0 1e-06 
0.0 -1.2485 0 2.0 1e-06 
0.0 -1.2484 0 2.0 1e-06 
0.0 -1.2483 0 2.0 1e-06 
0.0 -1.2482 0 2.0 1e-06 
0.0 -1.2481 0 2.0 1e-06 
0.0 -1.248 0 2.0 1e-06 
0.0 -1.2479 0 2.0 1e-06 
0.0 -1.2478 0 2.0 1e-06 
0.0 -1.2477 0 2.0 1e-06 
0.0 -1.2476 0 2.0 1e-06 
0.0 -1.2475 0 2.0 1e-06 
0.0 -1.2474 0 2.0 1e-06 
0.0 -1.2473 0 2.0 1e-06 
0.0 -1.2472 0 2.0 1e-06 
0.0 -1.2471 0 2.0 1e-06 
0.0 -1.247 0 2.0 1e-06 
0.0 -1.2469 0 2.0 1e-06 
0.0 -1.2468 0 2.0 1e-06 
0.0 -1.2467 0 2.0 1e-06 
0.0 -1.2466 0 2.0 1e-06 
0.0 -1.2465 0 2.0 1e-06 
0.0 -1.2464 0 2.0 1e-06 
0.0 -1.2463 0 2.0 1e-06 
0.0 -1.2462 0 2.0 1e-06 
0.0 -1.2461 0 2.0 1e-06 
0.0 -1.246 0 2.0 1e-06 
0.0 -1.2459 0 2.0 1e-06 
0.0 -1.2458 0 2.0 1e-06 
0.0 -1.2457 0 2.0 1e-06 
0.0 -1.2456 0 2.0 1e-06 
0.0 -1.2455 0 2.0 1e-06 
0.0 -1.2454 0 2.0 1e-06 
0.0 -1.2453 0 2.0 1e-06 
0.0 -1.2452 0 2.0 1e-06 
0.0 -1.2451 0 2.0 1e-06 
0.0 -1.245 0 2.0 1e-06 
0.0 -1.2449 0 2.0 1e-06 
0.0 -1.2448 0 2.0 1e-06 
0.0 -1.2447 0 2.0 1e-06 
0.0 -1.2446 0 2.0 1e-06 
0.0 -1.2445 0 2.0 1e-06 
0.0 -1.2444 0 2.0 1e-06 
0.0 -1.2443 0 2.0 1e-06 
0.0 -1.2442 0 2.0 1e-06 
0.0 -1.2441 0 2.0 1e-06 
0.0 -1.244 0 2.0 1e-06 
0.0 -1.2439 0 2.0 1e-06 
0.0 -1.2438 0 2.0 1e-06 
0.0 -1.2437 0 2.0 1e-06 
0.0 -1.2436 0 2.0 1e-06 
0.0 -1.2435 0 2.0 1e-06 
0.0 -1.2434 0 2.0 1e-06 
0.0 -1.2433 0 2.0 1e-06 
0.0 -1.2432 0 2.0 1e-06 
0.0 -1.2431 0 2.0 1e-06 
0.0 -1.243 0 2.0 1e-06 
0.0 -1.2429 0 2.0 1e-06 
0.0 -1.2428 0 2.0 1e-06 
0.0 -1.2427 0 2.0 1e-06 
0.0 -1.2426 0 2.0 1e-06 
0.0 -1.2425 0 2.0 1e-06 
0.0 -1.2424 0 2.0 1e-06 
0.0 -1.2423 0 2.0 1e-06 
0.0 -1.2422 0 2.0 1e-06 
0.0 -1.2421 0 2.0 1e-06 
0.0 -1.242 0 2.0 1e-06 
0.0 -1.2419 0 2.0 1e-06 
0.0 -1.2418 0 2.0 1e-06 
0.0 -1.2417 0 2.0 1e-06 
0.0 -1.2416 0 2.0 1e-06 
0.0 -1.2415 0 2.0 1e-06 
0.0 -1.2414 0 2.0 1e-06 
0.0 -1.2413 0 2.0 1e-06 
0.0 -1.2412 0 2.0 1e-06 
0.0 -1.2411 0 2.0 1e-06 
0.0 -1.241 0 2.0 1e-06 
0.0 -1.2409 0 2.0 1e-06 
0.0 -1.2408 0 2.0 1e-06 
0.0 -1.2407 0 2.0 1e-06 
0.0 -1.2406 0 2.0 1e-06 
0.0 -1.2405 0 2.0 1e-06 
0.0 -1.2404 0 2.0 1e-06 
0.0 -1.2403 0 2.0 1e-06 
0.0 -1.2402 0 2.0 1e-06 
0.0 -1.2401 0 2.0 1e-06 
0.0 -1.24 0 2.0 1e-06 
0.0 -1.2399 0 2.0 1e-06 
0.0 -1.2398 0 2.0 1e-06 
0.0 -1.2397 0 2.0 1e-06 
0.0 -1.2396 0 2.0 1e-06 
0.0 -1.2395 0 2.0 1e-06 
0.0 -1.2394 0 2.0 1e-06 
0.0 -1.2393 0 2.0 1e-06 
0.0 -1.2392 0 2.0 1e-06 
0.0 -1.2391 0 2.0 1e-06 
0.0 -1.239 0 2.0 1e-06 
0.0 -1.2389 0 2.0 1e-06 
0.0 -1.2388 0 2.0 1e-06 
0.0 -1.2387 0 2.0 1e-06 
0.0 -1.2386 0 2.0 1e-06 
0.0 -1.2385 0 2.0 1e-06 
0.0 -1.2384 0 2.0 1e-06 
0.0 -1.2383 0 2.0 1e-06 
0.0 -1.2382 0 2.0 1e-06 
0.0 -1.2381 0 2.0 1e-06 
0.0 -1.238 0 2.0 1e-06 
0.0 -1.2379 0 2.0 1e-06 
0.0 -1.2378 0 2.0 1e-06 
0.0 -1.2377 0 2.0 1e-06 
0.0 -1.2376 0 2.0 1e-06 
0.0 -1.2375 0 2.0 1e-06 
0.0 -1.2374 0 2.0 1e-06 
0.0 -1.2373 0 2.0 1e-06 
0.0 -1.2372 0 2.0 1e-06 
0.0 -1.2371 0 2.0 1e-06 
0.0 -1.237 0 2.0 1e-06 
0.0 -1.2369 0 2.0 1e-06 
0.0 -1.2368 0 2.0 1e-06 
0.0 -1.2367 0 2.0 1e-06 
0.0 -1.2366 0 2.0 1e-06 
0.0 -1.2365 0 2.0 1e-06 
0.0 -1.2364 0 2.0 1e-06 
0.0 -1.2363 0 2.0 1e-06 
0.0 -1.2362 0 2.0 1e-06 
0.0 -1.2361 0 2.0 1e-06 
0.0 -1.236 0 2.0 1e-06 
0.0 -1.2359 0 2.0 1e-06 
0.0 -1.2358 0 2.0 1e-06 
0.0 -1.2357 0 2.0 1e-06 
0.0 -1.2356 0 2.0 1e-06 
0.0 -1.2355 0 2.0 1e-06 
0.0 -1.2354 0 2.0 1e-06 
0.0 -1.2353 0 2.0 1e-06 
0.0 -1.2352 0 2.0 1e-06 
0.0 -1.2351 0 2.0 1e-06 
0.0 -1.235 0 2.0 1e-06 
0.0 -1.2349 0 2.0 1e-06 
0.0 -1.2348 0 2.0 1e-06 
0.0 -1.2347 0 2.0 1e-06 
0.0 -1.2346 0 2.0 1e-06 
0.0 -1.2345 0 2.0 1e-06 
0.0 -1.2344 0 2.0 1e-06 
0.0 -1.2343 0 2.0 1e-06 
0.0 -1.2342 0 2.0 1e-06 
0.0 -1.2341 0 2.0 1e-06 
0.0 -1.234 0 2.0 1e-06 
0.0 -1.2339 0 2.0 1e-06 
0.0 -1.2338 0 2.0 1e-06 
0.0 -1.2337 0 2.0 1e-06 
0.0 -1.2336 0 2.0 1e-06 
0.0 -1.2335 0 2.0 1e-06 
0.0 -1.2334 0 2.0 1e-06 
0.0 -1.2333 0 2.0 1e-06 
0.0 -1.2332 0 2.0 1e-06 
0.0 -1.2331 0 2.0 1e-06 
0.0 -1.233 0 2.0 1e-06 
0.0 -1.2329 0 2.0 1e-06 
0.0 -1.2328 0 2.0 1e-06 
0.0 -1.2327 0 2.0 1e-06 
0.0 -1.2326 0 2.0 1e-06 
0.0 -1.2325 0 2.0 1e-06 
0.0 -1.2324 0 2.0 1e-06 
0.0 -1.2323 0 2.0 1e-06 
0.0 -1.2322 0 2.0 1e-06 
0.0 -1.2321 0 2.0 1e-06 
0.0 -1.232 0 2.0 1e-06 
0.0 -1.2319 0 2.0 1e-06 
0.0 -1.2318 0 2.0 1e-06 
0.0 -1.2317 0 2.0 1e-06 
0.0 -1.2316 0 2.0 1e-06 
0.0 -1.2315 0 2.0 1e-06 
0.0 -1.2314 0 2.0 1e-06 
0.0 -1.2313 0 2.0 1e-06 
0.0 -1.2312 0 2.0 1e-06 
0.0 -1.2311 0 2.0 1e-06 
0.0 -1.231 0 2.0 1e-06 
0.0 -1.2309 0 2.0 1e-06 
0.0 -1.2308 0 2.0 1e-06 
0.0 -1.2307 0 2.0 1e-06 
0.0 -1.2306 0 2.0 1e-06 
0.0 -1.2305 0 2.0 1e-06 
0.0 -1.2304 0 2.0 1e-06 
0.0 -1.2303 0 2.0 1e-06 
0.0 -1.2302 0 2.0 1e-06 
0.0 -1.2301 0 2.0 1e-06 
0.0 -1.23 0 2.0 1e-06 
0.0 -1.2299 0 2.0 1e-06 
0.0 -1.2298 0 2.0 1e-06 
0.0 -1.2297 0 2.0 1e-06 
0.0 -1.2296 0 2.0 1e-06 
0.0 -1.2295 0 2.0 1e-06 
0.0 -1.2294 0 2.0 1e-06 
0.0 -1.2293 0 2.0 1e-06 
0.0 -1.2292 0 2.0 1e-06 
0.0 -1.2291 0 2.0 1e-06 
0.0 -1.229 0 2.0 1e-06 
0.0 -1.2289 0 2.0 1e-06 
0.0 -1.2288 0 2.0 1e-06 
0.0 -1.2287 0 2.0 1e-06 
0.0 -1.2286 0 2.0 1e-06 
0.0 -1.2285 0 2.0 1e-06 
0.0 -1.2284 0 2.0 1e-06 
0.0 -1.2283 0 2.0 1e-06 
0.0 -1.2282 0 2.0 1e-06 
0.0 -1.2281 0 2.0 1e-06 
0.0 -1.228 0 2.0 1e-06 
0.0 -1.2279 0 2.0 1e-06 
0.0 -1.2278 0 2.0 1e-06 
0.0 -1.2277 0 2.0 1e-06 
0.0 -1.2276 0 2.0 1e-06 
0.0 -1.2275 0 2.0 1e-06 
0.0 -1.2274 0 2.0 1e-06 
0.0 -1.2273 0 2.0 1e-06 
0.0 -1.2272 0 2.0 1e-06 
0.0 -1.2271 0 2.0 1e-06 
0.0 -1.227 0 2.0 1e-06 
0.0 -1.2269 0 2.0 1e-06 
0.0 -1.2268 0 2.0 1e-06 
0.0 -1.2267 0 2.0 1e-06 
0.0 -1.2266 0 2.0 1e-06 
0.0 -1.2265 0 2.0 1e-06 
0.0 -1.2264 0 2.0 1e-06 
0.0 -1.2263 0 2.0 1e-06 
0.0 -1.2262 0 2.0 1e-06 
0.0 -1.2261 0 2.0 1e-06 
0.0 -1.226 0 2.0 1e-06 
0.0 -1.2259 0 2.0 1e-06 
0.0 -1.2258 0 2.0 1e-06 
0.0 -1.2257 0 2.0 1e-06 
0.0 -1.2256 0 2.0 1e-06 
0.0 -1.2255 0 2.0 1e-06 
0.0 -1.2254 0 2.0 1e-06 
0.0 -1.2253 0 2.0 1e-06 
0.0 -1.2252 0 2.0 1e-06 
0.0 -1.2251 0 2.0 1e-06 
0.0 -1.225 0 2.0 1e-06 
0.0 -1.2249 0 2.0 1e-06 
0.0 -1.2248 0 2.0 1e-06 
0.0 -1.2247 0 2.0 1e-06 
0.0 -1.2246 0 2.0 1e-06 
0.0 -1.2245 0 2.0 1e-06 
0.0 -1.2244 0 2.0 1e-06 
0.0 -1.2243 0 2.0 1e-06 
0.0 -1.2242 0 2.0 1e-06 
0.0 -1.2241 0 2.0 1e-06 
0.0 -1.224 0 2.0 1e-06 
0.0 -1.2239 0 2.0 1e-06 
0.0 -1.2238 0 2.0 1e-06 
0.0 -1.2237 0 2.0 1e-06 
0.0 -1.2236 0 2.0 1e-06 
0.0 -1.2235 0 2.0 1e-06 
0.0 -1.2234 0 2.0 1e-06 
0.0 -1.2233 0 2.0 1e-06 
0.0 -1.2232 0 2.0 1e-06 
0.0 -1.2231 0 2.0 1e-06 
0.0 -1.223 0 2.0 1e-06 
0.0 -1.2229 0 2.0 1e-06 
0.0 -1.2228 0 2.0 1e-06 
0.0 -1.2227 0 2.0 1e-06 
0.0 -1.2226 0 2.0 1e-06 
0.0 -1.2225 0 2.0 1e-06 
0.0 -1.2224 0 2.0 1e-06 
0.0 -1.2223 0 2.0 1e-06 
0.0 -1.2222 0 2.0 1e-06 
0.0 -1.2221 0 2.0 1e-06 
0.0 -1.222 0 2.0 1e-06 
0.0 -1.2219 0 2.0 1e-06 
0.0 -1.2218 0 2.0 1e-06 
0.0 -1.2217 0 2.0 1e-06 
0.0 -1.2216 0 2.0 1e-06 
0.0 -1.2215 0 2.0 1e-06 
0.0 -1.2214 0 2.0 1e-06 
0.0 -1.2213 0 2.0 1e-06 
0.0 -1.2212 0 2.0 1e-06 
0.0 -1.2211 0 2.0 1e-06 
0.0 -1.221 0 2.0 1e-06 
0.0 -1.2209 0 2.0 1e-06 
0.0 -1.2208 0 2.0 1e-06 
0.0 -1.2207 0 2.0 1e-06 
0.0 -1.2206 0 2.0 1e-06 
0.0 -1.2205 0 2.0 1e-06 
0.0 -1.2204 0 2.0 1e-06 
0.0 -1.2203 0 2.0 1e-06 
0.0 -1.2202 0 2.0 1e-06 
0.0 -1.2201 0 2.0 1e-06 
0.0 -1.22 0 2.0 1e-06 
0.0 -1.2199 0 2.0 1e-06 
0.0 -1.2198 0 2.0 1e-06 
0.0 -1.2197 0 2.0 1e-06 
0.0 -1.2196 0 2.0 1e-06 
0.0 -1.2195 0 2.0 1e-06 
0.0 -1.2194 0 2.0 1e-06 
0.0 -1.2193 0 2.0 1e-06 
0.0 -1.2192 0 2.0 1e-06 
0.0 -1.2191 0 2.0 1e-06 
0.0 -1.219 0 2.0 1e-06 
0.0 -1.2189 0 2.0 1e-06 
0.0 -1.2188 0 2.0 1e-06 
0.0 -1.2187 0 2.0 1e-06 
0.0 -1.2186 0 2.0 1e-06 
0.0 -1.2185 0 2.0 1e-06 
0.0 -1.2184 0 2.0 1e-06 
0.0 -1.2183 0 2.0 1e-06 
0.0 -1.2182 0 2.0 1e-06 
0.0 -1.2181 0 2.0 1e-06 
0.0 -1.218 0 2.0 1e-06 
0.0 -1.2179 0 2.0 1e-06 
0.0 -1.2178 0 2.0 1e-06 
0.0 -1.2177 0 2.0 1e-06 
0.0 -1.2176 0 2.0 1e-06 
0.0 -1.2175 0 2.0 1e-06 
0.0 -1.2174 0 2.0 1e-06 
0.0 -1.2173 0 2.0 1e-06 
0.0 -1.2172 0 2.0 1e-06 
0.0 -1.2171 0 2.0 1e-06 
0.0 -1.217 0 2.0 1e-06 
0.0 -1.2169 0 2.0 1e-06 
0.0 -1.2168 0 2.0 1e-06 
0.0 -1.2167 0 2.0 1e-06 
0.0 -1.2166 0 2.0 1e-06 
0.0 -1.2165 0 2.0 1e-06 
0.0 -1.2164 0 2.0 1e-06 
0.0 -1.2163 0 2.0 1e-06 
0.0 -1.2162 0 2.0 1e-06 
0.0 -1.2161 0 2.0 1e-06 
0.0 -1.216 0 2.0 1e-06 
0.0 -1.2159 0 2.0 1e-06 
0.0 -1.2158 0 2.0 1e-06 
0.0 -1.2157 0 2.0 1e-06 
0.0 -1.2156 0 2.0 1e-06 
0.0 -1.2155 0 2.0 1e-06 
0.0 -1.2154 0 2.0 1e-06 
0.0 -1.2153 0 2.0 1e-06 
0.0 -1.2152 0 2.0 1e-06 
0.0 -1.2151 0 2.0 1e-06 
0.0 -1.215 0 2.0 1e-06 
0.0 -1.2149 0 2.0 1e-06 
0.0 -1.2148 0 2.0 1e-06 
0.0 -1.2147 0 2.0 1e-06 
0.0 -1.2146 0 2.0 1e-06 
0.0 -1.2145 0 2.0 1e-06 
0.0 -1.2144 0 2.0 1e-06 
0.0 -1.2143 0 2.0 1e-06 
0.0 -1.2142 0 2.0 1e-06 
0.0 -1.2141 0 2.0 1e-06 
0.0 -1.214 0 2.0 1e-06 
0.0 -1.2139 0 2.0 1e-06 
0.0 -1.2138 0 2.0 1e-06 
0.0 -1.2137 0 2.0 1e-06 
0.0 -1.2136 0 2.0 1e-06 
0.0 -1.2135 0 2.0 1e-06 
0.0 -1.2134 0 2.0 1e-06 
0.0 -1.2133 0 2.0 1e-06 
0.0 -1.2132 0 2.0 1e-06 
0.0 -1.2131 0 2.0 1e-06 
0.0 -1.213 0 2.0 1e-06 
0.0 -1.2129 0 2.0 1e-06 
0.0 -1.2128 0 2.0 1e-06 
0.0 -1.2127 0 2.0 1e-06 
0.0 -1.2126 0 2.0 1e-06 
0.0 -1.2125 0 2.0 1e-06 
0.0 -1.2124 0 2.0 1e-06 
0.0 -1.2123 0 2.0 1e-06 
0.0 -1.2122 0 2.0 1e-06 
0.0 -1.2121 0 2.0 1e-06 
0.0 -1.212 0 2.0 1e-06 
0.0 -1.2119 0 2.0 1e-06 
0.0 -1.2118 0 2.0 1e-06 
0.0 -1.2117 0 2.0 1e-06 
0.0 -1.2116 0 2.0 1e-06 
0.0 -1.2115 0 2.0 1e-06 
0.0 -1.2114 0 2.0 1e-06 
0.0 -1.2113 0 2.0 1e-06 
0.0 -1.2112 0 2.0 1e-06 
0.0 -1.2111 0 2.0 1e-06 
0.0 -1.211 0 2.0 1e-06 
0.0 -1.2109 0 2.0 1e-06 
0.0 -1.2108 0 2.0 1e-06 
0.0 -1.2107 0 2.0 1e-06 
0.0 -1.2106 0 2.0 1e-06 
0.0 -1.2105 0 2.0 1e-06 
0.0 -1.2104 0 2.0 1e-06 
0.0 -1.2103 0 2.0 1e-06 
0.0 -1.2102 0 2.0 1e-06 
0.0 -1.2101 0 2.0 1e-06 
0.0 -1.21 0 2.0 1e-06 
0.0 -1.2099 0 2.0 1e-06 
0.0 -1.2098 0 2.0 1e-06 
0.0 -1.2097 0 2.0 1e-06 
0.0 -1.2096 0 2.0 1e-06 
0.0 -1.2095 0 2.0 1e-06 
0.0 -1.2094 0 2.0 1e-06 
0.0 -1.2093 0 2.0 1e-06 
0.0 -1.2092 0 2.0 1e-06 
0.0 -1.2091 0 2.0 1e-06 
0.0 -1.209 0 2.0 1e-06 
0.0 -1.2089 0 2.0 1e-06 
0.0 -1.2088 0 2.0 1e-06 
0.0 -1.2087 0 2.0 1e-06 
0.0 -1.2086 0 2.0 1e-06 
0.0 -1.2085 0 2.0 1e-06 
0.0 -1.2084 0 2.0 1e-06 
0.0 -1.2083 0 2.0 1e-06 
0.0 -1.2082 0 2.0 1e-06 
0.0 -1.2081 0 2.0 1e-06 
0.0 -1.208 0 2.0 1e-06 
0.0 -1.2079 0 2.0 1e-06 
0.0 -1.2078 0 2.0 1e-06 
0.0 -1.2077 0 2.0 1e-06 
0.0 -1.2076 0 2.0 1e-06 
0.0 -1.2075 0 2.0 1e-06 
0.0 -1.2074 0 2.0 1e-06 
0.0 -1.2073 0 2.0 1e-06 
0.0 -1.2072 0 2.0 1e-06 
0.0 -1.2071 0 2.0 1e-06 
0.0 -1.207 0 2.0 1e-06 
0.0 -1.2069 0 2.0 1e-06 
0.0 -1.2068 0 2.0 1e-06 
0.0 -1.2067 0 2.0 1e-06 
0.0 -1.2066 0 2.0 1e-06 
0.0 -1.2065 0 2.0 1e-06 
0.0 -1.2064 0 2.0 1e-06 
0.0 -1.2063 0 2.0 1e-06 
0.0 -1.2062 0 2.0 1e-06 
0.0 -1.2061 0 2.0 1e-06 
0.0 -1.206 0 2.0 1e-06 
0.0 -1.2059 0 2.0 1e-06 
0.0 -1.2058 0 2.0 1e-06 
0.0 -1.2057 0 2.0 1e-06 
0.0 -1.2056 0 2.0 1e-06 
0.0 -1.2055 0 2.0 1e-06 
0.0 -1.2054 0 2.0 1e-06 
0.0 -1.2053 0 2.0 1e-06 
0.0 -1.2052 0 2.0 1e-06 
0.0 -1.2051 0 2.0 1e-06 
0.0 -1.205 0 2.0 1e-06 
0.0 -1.2049 0 2.0 1e-06 
0.0 -1.2048 0 2.0 1e-06 
0.0 -1.2047 0 2.0 1e-06 
0.0 -1.2046 0 2.0 1e-06 
0.0 -1.2045 0 2.0 1e-06 
0.0 -1.2044 0 2.0 1e-06 
0.0 -1.2043 0 2.0 1e-06 
0.0 -1.2042 0 2.0 1e-06 
0.0 -1.2041 0 2.0 1e-06 
0.0 -1.204 0 2.0 1e-06 
0.0 -1.2039 0 2.0 1e-06 
0.0 -1.2038 0 2.0 1e-06 
0.0 -1.2037 0 2.0 1e-06 
0.0 -1.2036 0 2.0 1e-06 
0.0 -1.2035 0 2.0 1e-06 
0.0 -1.2034 0 2.0 1e-06 
0.0 -1.2033 0 2.0 1e-06 
0.0 -1.2032 0 2.0 1e-06 
0.0 -1.2031 0 2.0 1e-06 
0.0 -1.203 0 2.0 1e-06 
0.0 -1.2029 0 2.0 1e-06 
0.0 -1.2028 0 2.0 1e-06 
0.0 -1.2027 0 2.0 1e-06 
0.0 -1.2026 0 2.0 1e-06 
0.0 -1.2025 0 2.0 1e-06 
0.0 -1.2024 0 2.0 1e-06 
0.0 -1.2023 0 2.0 1e-06 
0.0 -1.2022 0 2.0 1e-06 
0.0 -1.2021 0 2.0 1e-06 
0.0 -1.202 0 2.0 1e-06 
0.0 -1.2019 0 2.0 1e-06 
0.0 -1.2018 0 2.0 1e-06 
0.0 -1.2017 0 2.0 1e-06 
0.0 -1.2016 0 2.0 1e-06 
0.0 -1.2015 0 2.0 1e-06 
0.0 -1.2014 0 2.0 1e-06 
0.0 -1.2013 0 2.0 1e-06 
0.0 -1.2012 0 2.0 1e-06 
0.0 -1.2011 0 2.0 1e-06 
0.0 -1.201 0 2.0 1e-06 
0.0 -1.2009 0 2.0 1e-06 
0.0 -1.2008 0 2.0 1e-06 
0.0 -1.2007 0 2.0 1e-06 
0.0 -1.2006 0 2.0 1e-06 
0.0 -1.2005 0 2.0 1e-06 
0.0 -1.2004 0 2.0 1e-06 
0.0 -1.2003 0 2.0 1e-06 
0.0 -1.2002 0 2.0 1e-06 
0.0 -1.2001 0 2.0 1e-06 
0.0 -1.2 0 2.0 1e-06 
0.0 -1.1999 0 2.0 1e-06 
0.0 -1.1998 0 2.0 1e-06 
0.0 -1.1997 0 2.0 1e-06 
0.0 -1.1996 0 2.0 1e-06 
0.0 -1.1995 0 2.0 1e-06 
0.0 -1.1994 0 2.0 1e-06 
0.0 -1.1993 0 2.0 1e-06 
0.0 -1.1992 0 2.0 1e-06 
0.0 -1.1991 0 2.0 1e-06 
0.0 -1.199 0 2.0 1e-06 
0.0 -1.1989 0 2.0 1e-06 
0.0 -1.1988 0 2.0 1e-06 
0.0 -1.1987 0 2.0 1e-06 
0.0 -1.1986 0 2.0 1e-06 
0.0 -1.1985 0 2.0 1e-06 
0.0 -1.1984 0 2.0 1e-06 
0.0 -1.1983 0 2.0 1e-06 
0.0 -1.1982 0 2.0 1e-06 
0.0 -1.1981 0 2.0 1e-06 
0.0 -1.198 0 2.0 1e-06 
0.0 -1.1979 0 2.0 1e-06 
0.0 -1.1978 0 2.0 1e-06 
0.0 -1.1977 0 2.0 1e-06 
0.0 -1.1976 0 2.0 1e-06 
0.0 -1.1975 0 2.0 1e-06 
0.0 -1.1974 0 2.0 1e-06 
0.0 -1.1973 0 2.0 1e-06 
0.0 -1.1972 0 2.0 1e-06 
0.0 -1.1971 0 2.0 1e-06 
0.0 -1.197 0 2.0 1e-06 
0.0 -1.1969 0 2.0 1e-06 
0.0 -1.1968 0 2.0 1e-06 
0.0 -1.1967 0 2.0 1e-06 
0.0 -1.1966 0 2.0 1e-06 
0.0 -1.1965 0 2.0 1e-06 
0.0 -1.1964 0 2.0 1e-06 
0.0 -1.1963 0 2.0 1e-06 
0.0 -1.1962 0 2.0 1e-06 
0.0 -1.1961 0 2.0 1e-06 
0.0 -1.196 0 2.0 1e-06 
0.0 -1.1959 0 2.0 1e-06 
0.0 -1.1958 0 2.0 1e-06 
0.0 -1.1957 0 2.0 1e-06 
0.0 -1.1956 0 2.0 1e-06 
0.0 -1.1955 0 2.0 1e-06 
0.0 -1.1954 0 2.0 1e-06 
0.0 -1.1953 0 2.0 1e-06 
0.0 -1.1952 0 2.0 1e-06 
0.0 -1.1951 0 2.0 1e-06 
0.0 -1.195 0 2.0 1e-06 
0.0 -1.1949 0 2.0 1e-06 
0.0 -1.1948 0 2.0 1e-06 
0.0 -1.1947 0 2.0 1e-06 
0.0 -1.1946 0 2.0 1e-06 
0.0 -1.1945 0 2.0 1e-06 
0.0 -1.1944 0 2.0 1e-06 
0.0 -1.1943 0 2.0 1e-06 
0.0 -1.1942 0 2.0 1e-06 
0.0 -1.1941 0 2.0 1e-06 
0.0 -1.194 0 2.0 1e-06 
0.0 -1.1939 0 2.0 1e-06 
0.0 -1.1938 0 2.0 1e-06 
0.0 -1.1937 0 2.0 1e-06 
0.0 -1.1936 0 2.0 1e-06 
0.0 -1.1935 0 2.0 1e-06 
0.0 -1.1934 0 2.0 1e-06 
0.0 -1.1933 0 2.0 1e-06 
0.0 -1.1932 0 2.0 1e-06 
0.0 -1.1931 0 2.0 1e-06 
0.0 -1.193 0 2.0 1e-06 
0.0 -1.1929 0 2.0 1e-06 
0.0 -1.1928 0 2.0 1e-06 
0.0 -1.1927 0 2.0 1e-06 
0.0 -1.1926 0 2.0 1e-06 
0.0 -1.1925 0 2.0 1e-06 
0.0 -1.1924 0 2.0 1e-06 
0.0 -1.1923 0 2.0 1e-06 
0.0 -1.1922 0 2.0 1e-06 
0.0 -1.1921 0 2.0 1e-06 
0.0 -1.192 0 2.0 1e-06 
0.0 -1.1919 0 2.0 1e-06 
0.0 -1.1918 0 2.0 1e-06 
0.0 -1.1917 0 2.0 1e-06 
0.0 -1.1916 0 2.0 1e-06 
0.0 -1.1915 0 2.0 1e-06 
0.0 -1.1914 0 2.0 1e-06 
0.0 -1.1913 0 2.0 1e-06 
0.0 -1.1912 0 2.0 1e-06 
0.0 -1.1911 0 2.0 1e-06 
0.0 -1.191 0 2.0 1e-06 
0.0 -1.1909 0 2.0 1e-06 
0.0 -1.1908 0 2.0 1e-06 
0.0 -1.1907 0 2.0 1e-06 
0.0 -1.1906 0 2.0 1e-06 
0.0 -1.1905 0 2.0 1e-06 
0.0 -1.1904 0 2.0 1e-06 
0.0 -1.1903 0 2.0 1e-06 
0.0 -1.1902 0 2.0 1e-06 
0.0 -1.1901 0 2.0 1e-06 
0.0 -1.19 0 2.0 1e-06 
0.0 -1.1899 0 2.0 1e-06 
0.0 -1.1898 0 2.0 1e-06 
0.0 -1.1897 0 2.0 1e-06 
0.0 -1.1896 0 2.0 1e-06 
0.0 -1.1895 0 2.0 1e-06 
0.0 -1.1894 0 2.0 1e-06 
0.0 -1.1893 0 2.0 1e-06 
0.0 -1.1892 0 2.0 1e-06 
0.0 -1.1891 0 2.0 1e-06 
0.0 -1.189 0 2.0 1e-06 
0.0 -1.1889 0 2.0 1e-06 
0.0 -1.1888 0 2.0 1e-06 
0.0 -1.1887 0 2.0 1e-06 
0.0 -1.1886 0 2.0 1e-06 
0.0 -1.1885 0 2.0 1e-06 
0.0 -1.1884 0 2.0 1e-06 
0.0 -1.1883 0 2.0 1e-06 
0.0 -1.1882 0 2.0 1e-06 
0.0 -1.1881 0 2.0 1e-06 
0.0 -1.188 0 2.0 1e-06 
0.0 -1.1879 0 2.0 1e-06 
0.0 -1.1878 0 2.0 1e-06 
0.0 -1.1877 0 2.0 1e-06 
0.0 -1.1876 0 2.0 1e-06 
0.0 -1.1875 0 2.0 1e-06 
0.0 -1.1874 0 2.0 1e-06 
0.0 -1.1873 0 2.0 1e-06 
0.0 -1.1872 0 2.0 1e-06 
0.0 -1.1871 0 2.0 1e-06 
0.0 -1.187 0 2.0 1e-06 
0.0 -1.1869 0 2.0 1e-06 
0.0 -1.1868 0 2.0 1e-06 
0.0 -1.1867 0 2.0 1e-06 
0.0 -1.1866 0 2.0 1e-06 
0.0 -1.1865 0 2.0 1e-06 
0.0 -1.1864 0 2.0 1e-06 
0.0 -1.1863 0 2.0 1e-06 
0.0 -1.1862 0 2.0 1e-06 
0.0 -1.1861 0 2.0 1e-06 
0.0 -1.186 0 2.0 1e-06 
0.0 -1.1859 0 2.0 1e-06 
0.0 -1.1858 0 2.0 1e-06 
0.0 -1.1857 0 2.0 1e-06 
0.0 -1.1856 0 2.0 1e-06 
0.0 -1.1855 0 2.0 1e-06 
0.0 -1.1854 0 2.0 1e-06 
0.0 -1.1853 0 2.0 1e-06 
0.0 -1.1852 0 2.0 1e-06 
0.0 -1.1851 0 2.0 1e-06 
0.0 -1.185 0 2.0 1e-06 
0.0 -1.1849 0 2.0 1e-06 
0.0 -1.1848 0 2.0 1e-06 
0.0 -1.1847 0 2.0 1e-06 
0.0 -1.1846 0 2.0 1e-06 
0.0 -1.1845 0 2.0 1e-06 
0.0 -1.1844 0 2.0 1e-06 
0.0 -1.1843 0 2.0 1e-06 
0.0 -1.1842 0 2.0 1e-06 
0.0 -1.1841 0 2.0 1e-06 
0.0 -1.184 0 2.0 1e-06 
0.0 -1.1839 0 2.0 1e-06 
0.0 -1.1838 0 2.0 1e-06 
0.0 -1.1837 0 2.0 1e-06 
0.0 -1.1836 0 2.0 1e-06 
0.0 -1.1835 0 2.0 1e-06 
0.0 -1.1834 0 2.0 1e-06 
0.0 -1.1833 0 2.0 1e-06 
0.0 -1.1832 0 2.0 1e-06 
0.0 -1.1831 0 2.0 1e-06 
0.0 -1.183 0 2.0 1e-06 
0.0 -1.1829 0 2.0 1e-06 
0.0 -1.1828 0 2.0 1e-06 
0.0 -1.1827 0 2.0 1e-06 
0.0 -1.1826 0 2.0 1e-06 
0.0 -1.1825 0 2.0 1e-06 
0.0 -1.1824 0 2.0 1e-06 
0.0 -1.1823 0 2.0 1e-06 
0.0 -1.1822 0 2.0 1e-06 
0.0 -1.1821 0 2.0 1e-06 
0.0 -1.182 0 2.0 1e-06 
0.0 -1.1819 0 2.0 1e-06 
0.0 -1.1818 0 2.0 1e-06 
0.0 -1.1817 0 2.0 1e-06 
0.0 -1.1816 0 2.0 1e-06 
0.0 -1.1815 0 2.0 1e-06 
0.0 -1.1814 0 2.0 1e-06 
0.0 -1.1813 0 2.0 1e-06 
0.0 -1.1812 0 2.0 1e-06 
0.0 -1.1811 0 2.0 1e-06 
0.0 -1.181 0 2.0 1e-06 
0.0 -1.1809 0 2.0 1e-06 
0.0 -1.1808 0 2.0 1e-06 
0.0 -1.1807 0 2.0 1e-06 
0.0 -1.1806 0 2.0 1e-06 
0.0 -1.1805 0 2.0 1e-06 
0.0 -1.1804 0 2.0 1e-06 
0.0 -1.1803 0 2.0 1e-06 
0.0 -1.1802 0 2.0 1e-06 
0.0 -1.1801 0 2.0 1e-06 
0.0 -1.18 0 2.0 1e-06 
0.0 -1.1799 0 2.0 1e-06 
0.0 -1.1798 0 2.0 1e-06 
0.0 -1.1797 0 2.0 1e-06 
0.0 -1.1796 0 2.0 1e-06 
0.0 -1.1795 0 2.0 1e-06 
0.0 -1.1794 0 2.0 1e-06 
0.0 -1.1793 0 2.0 1e-06 
0.0 -1.1792 0 2.0 1e-06 
0.0 -1.1791 0 2.0 1e-06 
0.0 -1.179 0 2.0 1e-06 
0.0 -1.1789 0 2.0 1e-06 
0.0 -1.1788 0 2.0 1e-06 
0.0 -1.1787 0 2.0 1e-06 
0.0 -1.1786 0 2.0 1e-06 
0.0 -1.1785 0 2.0 1e-06 
0.0 -1.1784 0 2.0 1e-06 
0.0 -1.1783 0 2.0 1e-06 
0.0 -1.1782 0 2.0 1e-06 
0.0 -1.1781 0 2.0 1e-06 
0.0 -1.178 0 2.0 1e-06 
0.0 -1.1779 0 2.0 1e-06 
0.0 -1.1778 0 2.0 1e-06 
0.0 -1.1777 0 2.0 1e-06 
0.0 -1.1776 0 2.0 1e-06 
0.0 -1.1775 0 2.0 1e-06 
0.0 -1.1774 0 2.0 1e-06 
0.0 -1.1773 0 2.0 1e-06 
0.0 -1.1772 0 2.0 1e-06 
0.0 -1.1771 0 2.0 1e-06 
0.0 -1.177 0 2.0 1e-06 
0.0 -1.1769 0 2.0 1e-06 
0.0 -1.1768 0 2.0 1e-06 
0.0 -1.1767 0 2.0 1e-06 
0.0 -1.1766 0 2.0 1e-06 
0.0 -1.1765 0 2.0 1e-06 
0.0 -1.1764 0 2.0 1e-06 
0.0 -1.1763 0 2.0 1e-06 
0.0 -1.1762 0 2.0 1e-06 
0.0 -1.1761 0 2.0 1e-06 
0.0 -1.176 0 2.0 1e-06 
0.0 -1.1759 0 2.0 1e-06 
0.0 -1.1758 0 2.0 1e-06 
0.0 -1.1757 0 2.0 1e-06 
0.0 -1.1756 0 2.0 1e-06 
0.0 -1.1755 0 2.0 1e-06 
0.0 -1.1754 0 2.0 1e-06 
0.0 -1.1753 0 2.0 1e-06 
0.0 -1.1752 0 2.0 1e-06 
0.0 -1.1751 0 2.0 1e-06 
0.0 -1.175 0 2.0 1e-06 
0.0 -1.1749 0 2.0 1e-06 
0.0 -1.1748 0 2.0 1e-06 
0.0 -1.1747 0 2.0 1e-06 
0.0 -1.1746 0 2.0 1e-06 
0.0 -1.1745 0 2.0 1e-06 
0.0 -1.1744 0 2.0 1e-06 
0.0 -1.1743 0 2.0 1e-06 
0.0 -1.1742 0 2.0 1e-06 
0.0 -1.1741 0 2.0 1e-06 
0.0 -1.174 0 2.0 1e-06 
0.0 -1.1739 0 2.0 1e-06 
0.0 -1.1738 0 2.0 1e-06 
0.0 -1.1737 0 2.0 1e-06 
0.0 -1.1736 0 2.0 1e-06 
0.0 -1.1735 0 2.0 1e-06 
0.0 -1.1734 0 2.0 1e-06 
0.0 -1.1733 0 2.0 1e-06 
0.0 -1.1732 0 2.0 1e-06 
0.0 -1.1731 0 2.0 1e-06 
0.0 -1.173 0 2.0 1e-06 
0.0 -1.1729 0 2.0 1e-06 
0.0 -1.1728 0 2.0 1e-06 
0.0 -1.1727 0 2.0 1e-06 
0.0 -1.1726 0 2.0 1e-06 
0.0 -1.1725 0 2.0 1e-06 
0.0 -1.1724 0 2.0 1e-06 
0.0 -1.1723 0 2.0 1e-06 
0.0 -1.1722 0 2.0 1e-06 
0.0 -1.1721 0 2.0 1e-06 
0.0 -1.172 0 2.0 1e-06 
0.0 -1.1719 0 2.0 1e-06 
0.0 -1.1718 0 2.0 1e-06 
0.0 -1.1717 0 2.0 1e-06 
0.0 -1.1716 0 2.0 1e-06 
0.0 -1.1715 0 2.0 1e-06 
0.0 -1.1714 0 2.0 1e-06 
0.0 -1.1713 0 2.0 1e-06 
0.0 -1.1712 0 2.0 1e-06 
0.0 -1.1711 0 2.0 1e-06 
0.0 -1.171 0 2.0 1e-06 
0.0 -1.1709 0 2.0 1e-06 
0.0 -1.1708 0 2.0 1e-06 
0.0 -1.1707 0 2.0 1e-06 
0.0 -1.1706 0 2.0 1e-06 
0.0 -1.1705 0 2.0 1e-06 
0.0 -1.1704 0 2.0 1e-06 
0.0 -1.1703 0 2.0 1e-06 
0.0 -1.1702 0 2.0 1e-06 
0.0 -1.1701 0 2.0 1e-06 
0.0 -1.17 0 2.0 1e-06 
0.0 -1.1699 0 2.0 1e-06 
0.0 -1.1698 0 2.0 1e-06 
0.0 -1.1697 0 2.0 1e-06 
0.0 -1.1696 0 2.0 1e-06 
0.0 -1.1695 0 2.0 1e-06 
0.0 -1.1694 0 2.0 1e-06 
0.0 -1.1693 0 2.0 1e-06 
0.0 -1.1692 0 2.0 1e-06 
0.0 -1.1691 0 2.0 1e-06 
0.0 -1.169 0 2.0 1e-06 
0.0 -1.1689 0 2.0 1e-06 
0.0 -1.1688 0 2.0 1e-06 
0.0 -1.1687 0 2.0 1e-06 
0.0 -1.1686 0 2.0 1e-06 
0.0 -1.1685 0 2.0 1e-06 
0.0 -1.1684 0 2.0 1e-06 
0.0 -1.1683 0 2.0 1e-06 
0.0 -1.1682 0 2.0 1e-06 
0.0 -1.1681 0 2.0 1e-06 
0.0 -1.168 0 2.0 1e-06 
0.0 -1.1679 0 2.0 1e-06 
0.0 -1.1678 0 2.0 1e-06 
0.0 -1.1677 0 2.0 1e-06 
0.0 -1.1676 0 2.0 1e-06 
0.0 -1.1675 0 2.0 1e-06 
0.0 -1.1674 0 2.0 1e-06 
0.0 -1.1673 0 2.0 1e-06 
0.0 -1.1672 0 2.0 1e-06 
0.0 -1.1671 0 2.0 1e-06 
0.0 -1.167 0 2.0 1e-06 
0.0 -1.1669 0 2.0 1e-06 
0.0 -1.1668 0 2.0 1e-06 
0.0 -1.1667 0 2.0 1e-06 
0.0 -1.1666 0 2.0 1e-06 
0.0 -1.1665 0 2.0 1e-06 
0.0 -1.1664 0 2.0 1e-06 
0.0 -1.1663 0 2.0 1e-06 
0.0 -1.1662 0 2.0 1e-06 
0.0 -1.1661 0 2.0 1e-06 
0.0 -1.166 0 2.0 1e-06 
0.0 -1.1659 0 2.0 1e-06 
0.0 -1.1658 0 2.0 1e-06 
0.0 -1.1657 0 2.0 1e-06 
0.0 -1.1656 0 2.0 1e-06 
0.0 -1.1655 0 2.0 1e-06 
0.0 -1.1654 0 2.0 1e-06 
0.0 -1.1653 0 2.0 1e-06 
0.0 -1.1652 0 2.0 1e-06 
0.0 -1.1651 0 2.0 1e-06 
0.0 -1.165 0 2.0 1e-06 
0.0 -1.1649 0 2.0 1e-06 
0.0 -1.1648 0 2.0 1e-06 
0.0 -1.1647 0 2.0 1e-06 
0.0 -1.1646 0 2.0 1e-06 
0.0 -1.1645 0 2.0 1e-06 
0.0 -1.1644 0 2.0 1e-06 
0.0 -1.1643 0 2.0 1e-06 
0.0 -1.1642 0 2.0 1e-06 
0.0 -1.1641 0 2.0 1e-06 
0.0 -1.164 0 2.0 1e-06 
0.0 -1.1639 0 2.0 1e-06 
0.0 -1.1638 0 2.0 1e-06 
0.0 -1.1637 0 2.0 1e-06 
0.0 -1.1636 0 2.0 1e-06 
0.0 -1.1635 0 2.0 1e-06 
0.0 -1.1634 0 2.0 1e-06 
0.0 -1.1633 0 2.0 1e-06 
0.0 -1.1632 0 2.0 1e-06 
0.0 -1.1631 0 2.0 1e-06 
0.0 -1.163 0 2.0 1e-06 
0.0 -1.1629 0 2.0 1e-06 
0.0 -1.1628 0 2.0 1e-06 
0.0 -1.1627 0 2.0 1e-06 
0.0 -1.1626 0 2.0 1e-06 
0.0 -1.1625 0 2.0 1e-06 
0.0 -1.1624 0 2.0 1e-06 
0.0 -1.1623 0 2.0 1e-06 
0.0 -1.1622 0 2.0 1e-06 
0.0 -1.1621 0 2.0 1e-06 
0.0 -1.162 0 2.0 1e-06 
0.0 -1.1619 0 2.0 1e-06 
0.0 -1.1618 0 2.0 1e-06 
0.0 -1.1617 0 2.0 1e-06 
0.0 -1.1616 0 2.0 1e-06 
0.0 -1.1615 0 2.0 1e-06 
0.0 -1.1614 0 2.0 1e-06 
0.0 -1.1613 0 2.0 1e-06 
0.0 -1.1612 0 2.0 1e-06 
0.0 -1.1611 0 2.0 1e-06 
0.0 -1.161 0 2.0 1e-06 
0.0 -1.1609 0 2.0 1e-06 
0.0 -1.1608 0 2.0 1e-06 
0.0 -1.1607 0 2.0 1e-06 
0.0 -1.1606 0 2.0 1e-06 
0.0 -1.1605 0 2.0 1e-06 
0.0 -1.1604 0 2.0 1e-06 
0.0 -1.1603 0 2.0 1e-06 
0.0 -1.1602 0 2.0 1e-06 
0.0 -1.1601 0 2.0 1e-06 
0.0 -1.16 0 2.0 1e-06 
0.0 -1.1599 0 2.0 1e-06 
0.0 -1.1598 0 2.0 1e-06 
0.0 -1.1597 0 2.0 1e-06 
0.0 -1.1596 0 2.0 1e-06 
0.0 -1.1595 0 2.0 1e-06 
0.0 -1.1594 0 2.0 1e-06 
0.0 -1.1593 0 2.0 1e-06 
0.0 -1.1592 0 2.0 1e-06 
0.0 -1.1591 0 2.0 1e-06 
0.0 -1.159 0 2.0 1e-06 
0.0 -1.1589 0 2.0 1e-06 
0.0 -1.1588 0 2.0 1e-06 
0.0 -1.1587 0 2.0 1e-06 
0.0 -1.1586 0 2.0 1e-06 
0.0 -1.1585 0 2.0 1e-06 
0.0 -1.1584 0 2.0 1e-06 
0.0 -1.1583 0 2.0 1e-06 
0.0 -1.1582 0 2.0 1e-06 
0.0 -1.1581 0 2.0 1e-06 
0.0 -1.158 0 2.0 1e-06 
0.0 -1.1579 0 2.0 1e-06 
0.0 -1.1578 0 2.0 1e-06 
0.0 -1.1577 0 2.0 1e-06 
0.0 -1.1576 0 2.0 1e-06 
0.0 -1.1575 0 2.0 1e-06 
0.0 -1.1574 0 2.0 1e-06 
0.0 -1.1573 0 2.0 1e-06 
0.0 -1.1572 0 2.0 1e-06 
0.0 -1.1571 0 2.0 1e-06 
0.0 -1.157 0 2.0 1e-06 
0.0 -1.1569 0 2.0 1e-06 
0.0 -1.1568 0 2.0 1e-06 
0.0 -1.1567 0 2.0 1e-06 
0.0 -1.1566 0 2.0 1e-06 
0.0 -1.1565 0 2.0 1e-06 
0.0 -1.1564 0 2.0 1e-06 
0.0 -1.1563 0 2.0 1e-06 
0.0 -1.1562 0 2.0 1e-06 
0.0 -1.1561 0 2.0 1e-06 
0.0 -1.156 0 2.0 1e-06 
0.0 -1.1559 0 2.0 1e-06 
0.0 -1.1558 0 2.0 1e-06 
0.0 -1.1557 0 2.0 1e-06 
0.0 -1.1556 0 2.0 1e-06 
0.0 -1.1555 0 2.0 1e-06 
0.0 -1.1554 0 2.0 1e-06 
0.0 -1.1553 0 2.0 1e-06 
0.0 -1.1552 0 2.0 1e-06 
0.0 -1.1551 0 2.0 1e-06 
0.0 -1.155 0 2.0 1e-06 
0.0 -1.1549 0 2.0 1e-06 
0.0 -1.1548 0 2.0 1e-06 
0.0 -1.1547 0 2.0 1e-06 
0.0 -1.1546 0 2.0 1e-06 
0.0 -1.1545 0 2.0 1e-06 
0.0 -1.1544 0 2.0 1e-06 
0.0 -1.1543 0 2.0 1e-06 
0.0 -1.1542 0 2.0 1e-06 
0.0 -1.1541 0 2.0 1e-06 
0.0 -1.154 0 2.0 1e-06 
0.0 -1.1539 0 2.0 1e-06 
0.0 -1.1538 0 2.0 1e-06 
0.0 -1.1537 0 2.0 1e-06 
0.0 -1.1536 0 2.0 1e-06 
0.0 -1.1535 0 2.0 1e-06 
0.0 -1.1534 0 2.0 1e-06 
0.0 -1.1533 0 2.0 1e-06 
0.0 -1.1532 0 2.0 1e-06 
0.0 -1.1531 0 2.0 1e-06 
0.0 -1.153 0 2.0 1e-06 
0.0 -1.1529 0 2.0 1e-06 
0.0 -1.1528 0 2.0 1e-06 
0.0 -1.1527 0 2.0 1e-06 
0.0 -1.1526 0 2.0 1e-06 
0.0 -1.1525 0 2.0 1e-06 
0.0 -1.1524 0 2.0 1e-06 
0.0 -1.1523 0 2.0 1e-06 
0.0 -1.1522 0 2.0 1e-06 
0.0 -1.1521 0 2.0 1e-06 
0.0 -1.152 0 2.0 1e-06 
0.0 -1.1519 0 2.0 1e-06 
0.0 -1.1518 0 2.0 1e-06 
0.0 -1.1517 0 2.0 1e-06 
0.0 -1.1516 0 2.0 1e-06 
0.0 -1.1515 0 2.0 1e-06 
0.0 -1.1514 0 2.0 1e-06 
0.0 -1.1513 0 2.0 1e-06 
0.0 -1.1512 0 2.0 1e-06 
0.0 -1.1511 0 2.0 1e-06 
0.0 -1.151 0 2.0 1e-06 
0.0 -1.1509 0 2.0 1e-06 
0.0 -1.1508 0 2.0 1e-06 
0.0 -1.1507 0 2.0 1e-06 
0.0 -1.1506 0 2.0 1e-06 
0.0 -1.1505 0 2.0 1e-06 
0.0 -1.1504 0 2.0 1e-06 
0.0 -1.1503 0 2.0 1e-06 
0.0 -1.1502 0 2.0 1e-06 
0.0 -1.1501 0 2.0 1e-06 
0.0 -1.15 0 2.0 1e-06 
0.0 -1.1499 0 2.0 1e-06 
0.0 -1.1498 0 2.0 1e-06 
0.0 -1.1497 0 2.0 1e-06 
0.0 -1.1496 0 2.0 1e-06 
0.0 -1.1495 0 2.0 1e-06 
0.0 -1.1494 0 2.0 1e-06 
0.0 -1.1493 0 2.0 1e-06 
0.0 -1.1492 0 2.0 1e-06 
0.0 -1.1491 0 2.0 1e-06 
0.0 -1.149 0 2.0 1e-06 
0.0 -1.1489 0 2.0 1e-06 
0.0 -1.1488 0 2.0 1e-06 
0.0 -1.1487 0 2.0 1e-06 
0.0 -1.1486 0 2.0 1e-06 
0.0 -1.1485 0 2.0 1e-06 
0.0 -1.1484 0 2.0 1e-06 
0.0 -1.1483 0 2.0 1e-06 
0.0 -1.1482 0 2.0 1e-06 
0.0 -1.1481 0 2.0 1e-06 
0.0 -1.148 0 2.0 1e-06 
0.0 -1.1479 0 2.0 1e-06 
0.0 -1.1478 0 2.0 1e-06 
0.0 -1.1477 0 2.0 1e-06 
0.0 -1.1476 0 2.0 1e-06 
0.0 -1.1475 0 2.0 1e-06 
0.0 -1.1474 0 2.0 1e-06 
0.0 -1.1473 0 2.0 1e-06 
0.0 -1.1472 0 2.0 1e-06 
0.0 -1.1471 0 2.0 1e-06 
0.0 -1.147 0 2.0 1e-06 
0.0 -1.1469 0 2.0 1e-06 
0.0 -1.1468 0 2.0 1e-06 
0.0 -1.1467 0 2.0 1e-06 
0.0 -1.1466 0 2.0 1e-06 
0.0 -1.1465 0 2.0 1e-06 
0.0 -1.1464 0 2.0 1e-06 
0.0 -1.1463 0 2.0 1e-06 
0.0 -1.1462 0 2.0 1e-06 
0.0 -1.1461 0 2.0 1e-06 
0.0 -1.146 0 2.0 1e-06 
0.0 -1.1459 0 2.0 1e-06 
0.0 -1.1458 0 2.0 1e-06 
0.0 -1.1457 0 2.0 1e-06 
0.0 -1.1456 0 2.0 1e-06 
0.0 -1.1455 0 2.0 1e-06 
0.0 -1.1454 0 2.0 1e-06 
0.0 -1.1453 0 2.0 1e-06 
0.0 -1.1452 0 2.0 1e-06 
0.0 -1.1451 0 2.0 1e-06 
0.0 -1.145 0 2.0 1e-06 
0.0 -1.1449 0 2.0 1e-06 
0.0 -1.1448 0 2.0 1e-06 
0.0 -1.1447 0 2.0 1e-06 
0.0 -1.1446 0 2.0 1e-06 
0.0 -1.1445 0 2.0 1e-06 
0.0 -1.1444 0 2.0 1e-06 
0.0 -1.1443 0 2.0 1e-06 
0.0 -1.1442 0 2.0 1e-06 
0.0 -1.1441 0 2.0 1e-06 
0.0 -1.144 0 2.0 1e-06 
0.0 -1.1439 0 2.0 1e-06 
0.0 -1.1438 0 2.0 1e-06 
0.0 -1.1437 0 2.0 1e-06 
0.0 -1.1436 0 2.0 1e-06 
0.0 -1.1435 0 2.0 1e-06 
0.0 -1.1434 0 2.0 1e-06 
0.0 -1.1433 0 2.0 1e-06 
0.0 -1.1432 0 2.0 1e-06 
0.0 -1.1431 0 2.0 1e-06 
0.0 -1.143 0 2.0 1e-06 
0.0 -1.1429 0 2.0 1e-06 
0.0 -1.1428 0 2.0 1e-06 
0.0 -1.1427 0 2.0 1e-06 
0.0 -1.1426 0 2.0 1e-06 
0.0 -1.1425 0 2.0 1e-06 
0.0 -1.1424 0 2.0 1e-06 
0.0 -1.1423 0 2.0 1e-06 
0.0 -1.1422 0 2.0 1e-06 
0.0 -1.1421 0 2.0 1e-06 
0.0 -1.142 0 2.0 1e-06 
0.0 -1.1419 0 2.0 1e-06 
0.0 -1.1418 0 2.0 1e-06 
0.0 -1.1417 0 2.0 1e-06 
0.0 -1.1416 0 2.0 1e-06 
0.0 -1.1415 0 2.0 1e-06 
0.0 -1.1414 0 2.0 1e-06 
0.0 -1.1413 0 2.0 1e-06 
0.0 -1.1412 0 2.0 1e-06 
0.0 -1.1411 0 2.0 1e-06 
0.0 -1.141 0 2.0 1e-06 
0.0 -1.1409 0 2.0 1e-06 
0.0 -1.1408 0 2.0 1e-06 
0.0 -1.1407 0 2.0 1e-06 
0.0 -1.1406 0 2.0 1e-06 
0.0 -1.1405 0 2.0 1e-06 
0.0 -1.1404 0 2.0 1e-06 
0.0 -1.1403 0 2.0 1e-06 
0.0 -1.1402 0 2.0 1e-06 
0.0 -1.1401 0 2.0 1e-06 
0.0 -1.14 0 2.0 1e-06 
0.0 -1.1399 0 2.0 1e-06 
0.0 -1.1398 0 2.0 1e-06 
0.0 -1.1397 0 2.0 1e-06 
0.0 -1.1396 0 2.0 1e-06 
0.0 -1.1395 0 2.0 1e-06 
0.0 -1.1394 0 2.0 1e-06 
0.0 -1.1393 0 2.0 1e-06 
0.0 -1.1392 0 2.0 1e-06 
0.0 -1.1391 0 2.0 1e-06 
0.0 -1.139 0 2.0 1e-06 
0.0 -1.1389 0 2.0 1e-06 
0.0 -1.1388 0 2.0 1e-06 
0.0 -1.1387 0 2.0 1e-06 
0.0 -1.1386 0 2.0 1e-06 
0.0 -1.1385 0 2.0 1e-06 
0.0 -1.1384 0 2.0 1e-06 
0.0 -1.1383 0 2.0 1e-06 
0.0 -1.1382 0 2.0 1e-06 
0.0 -1.1381 0 2.0 1e-06 
0.0 -1.138 0 2.0 1e-06 
0.0 -1.1379 0 2.0 1e-06 
0.0 -1.1378 0 2.0 1e-06 
0.0 -1.1377 0 2.0 1e-06 
0.0 -1.1376 0 2.0 1e-06 
0.0 -1.1375 0 2.0 1e-06 
0.0 -1.1374 0 2.0 1e-06 
0.0 -1.1373 0 2.0 1e-06 
0.0 -1.1372 0 2.0 1e-06 
0.0 -1.1371 0 2.0 1e-06 
0.0 -1.137 0 2.0 1e-06 
0.0 -1.1369 0 2.0 1e-06 
0.0 -1.1368 0 2.0 1e-06 
0.0 -1.1367 0 2.0 1e-06 
0.0 -1.1366 0 2.0 1e-06 
0.0 -1.1365 0 2.0 1e-06 
0.0 -1.1364 0 2.0 1e-06 
0.0 -1.1363 0 2.0 1e-06 
0.0 -1.1362 0 2.0 1e-06 
0.0 -1.1361 0 2.0 1e-06 
0.0 -1.136 0 2.0 1e-06 
0.0 -1.1359 0 2.0 1e-06 
0.0 -1.1358 0 2.0 1e-06 
0.0 -1.1357 0 2.0 1e-06 
0.0 -1.1356 0 2.0 1e-06 
0.0 -1.1355 0 2.0 1e-06 
0.0 -1.1354 0 2.0 1e-06 
0.0 -1.1353 0 2.0 1e-06 
0.0 -1.1352 0 2.0 1e-06 
0.0 -1.1351 0 2.0 1e-06 
0.0 -1.135 0 2.0 1e-06 
0.0 -1.1349 0 2.0 1e-06 
0.0 -1.1348 0 2.0 1e-06 
0.0 -1.1347 0 2.0 1e-06 
0.0 -1.1346 0 2.0 1e-06 
0.0 -1.1345 0 2.0 1e-06 
0.0 -1.1344 0 2.0 1e-06 
0.0 -1.1343 0 2.0 1e-06 
0.0 -1.1342 0 2.0 1e-06 
0.0 -1.1341 0 2.0 1e-06 
0.0 -1.134 0 2.0 1e-06 
0.0 -1.1339 0 2.0 1e-06 
0.0 -1.1338 0 2.0 1e-06 
0.0 -1.1337 0 2.0 1e-06 
0.0 -1.1336 0 2.0 1e-06 
0.0 -1.1335 0 2.0 1e-06 
0.0 -1.1334 0 2.0 1e-06 
0.0 -1.1333 0 2.0 1e-06 
0.0 -1.1332 0 2.0 1e-06 
0.0 -1.1331 0 2.0 1e-06 
0.0 -1.133 0 2.0 1e-06 
0.0 -1.1329 0 2.0 1e-06 
0.0 -1.1328 0 2.0 1e-06 
0.0 -1.1327 0 2.0 1e-06 
0.0 -1.1326 0 2.0 1e-06 
0.0 -1.1325 0 2.0 1e-06 
0.0 -1.1324 0 2.0 1e-06 
0.0 -1.1323 0 2.0 1e-06 
0.0 -1.1322 0 2.0 1e-06 
0.0 -1.1321 0 2.0 1e-06 
0.0 -1.132 0 2.0 1e-06 
0.0 -1.1319 0 2.0 1e-06 
0.0 -1.1318 0 2.0 1e-06 
0.0 -1.1317 0 2.0 1e-06 
0.0 -1.1316 0 2.0 1e-06 
0.0 -1.1315 0 2.0 1e-06 
0.0 -1.1314 0 2.0 1e-06 
0.0 -1.1313 0 2.0 1e-06 
0.0 -1.1312 0 2.0 1e-06 
0.0 -1.1311 0 2.0 1e-06 
0.0 -1.131 0 2.0 1e-06 
0.0 -1.1309 0 2.0 1e-06 
0.0 -1.1308 0 2.0 1e-06 
0.0 -1.1307 0 2.0 1e-06 
0.0 -1.1306 0 2.0 1e-06 
0.0 -1.1305 0 2.0 1e-06 
0.0 -1.1304 0 2.0 1e-06 
0.0 -1.1303 0 2.0 1e-06 
0.0 -1.1302 0 2.0 1e-06 
0.0 -1.1301 0 2.0 1e-06 
0.0 -1.13 0 2.0 1e-06 
0.0 -1.1299 0 2.0 1e-06 
0.0 -1.1298 0 2.0 1e-06 
0.0 -1.1297 0 2.0 1e-06 
0.0 -1.1296 0 2.0 1e-06 
0.0 -1.1295 0 2.0 1e-06 
0.0 -1.1294 0 2.0 1e-06 
0.0 -1.1293 0 2.0 1e-06 
0.0 -1.1292 0 2.0 1e-06 
0.0 -1.1291 0 2.0 1e-06 
0.0 -1.129 0 2.0 1e-06 
0.0 -1.1289 0 2.0 1e-06 
0.0 -1.1288 0 2.0 1e-06 
0.0 -1.1287 0 2.0 1e-06 
0.0 -1.1286 0 2.0 1e-06 
0.0 -1.1285 0 2.0 1e-06 
0.0 -1.1284 0 2.0 1e-06 
0.0 -1.1283 0 2.0 1e-06 
0.0 -1.1282 0 2.0 1e-06 
0.0 -1.1281 0 2.0 1e-06 
0.0 -1.128 0 2.0 1e-06 
0.0 -1.1279 0 2.0 1e-06 
0.0 -1.1278 0 2.0 1e-06 
0.0 -1.1277 0 2.0 1e-06 
0.0 -1.1276 0 2.0 1e-06 
0.0 -1.1275 0 2.0 1e-06 
0.0 -1.1274 0 2.0 1e-06 
0.0 -1.1273 0 2.0 1e-06 
0.0 -1.1272 0 2.0 1e-06 
0.0 -1.1271 0 2.0 1e-06 
0.0 -1.127 0 2.0 1e-06 
0.0 -1.1269 0 2.0 1e-06 
0.0 -1.1268 0 2.0 1e-06 
0.0 -1.1267 0 2.0 1e-06 
0.0 -1.1266 0 2.0 1e-06 
0.0 -1.1265 0 2.0 1e-06 
0.0 -1.1264 0 2.0 1e-06 
0.0 -1.1263 0 2.0 1e-06 
0.0 -1.1262 0 2.0 1e-06 
0.0 -1.1261 0 2.0 1e-06 
0.0 -1.126 0 2.0 1e-06 
0.0 -1.1259 0 2.0 1e-06 
0.0 -1.1258 0 2.0 1e-06 
0.0 -1.1257 0 2.0 1e-06 
0.0 -1.1256 0 2.0 1e-06 
0.0 -1.1255 0 2.0 1e-06 
0.0 -1.1254 0 2.0 1e-06 
0.0 -1.1253 0 2.0 1e-06 
0.0 -1.1252 0 2.0 1e-06 
0.0 -1.1251 0 2.0 1e-06 
0.0 -1.125 0 2.0 1e-06 
0.0 -1.1249 0 2.0 1e-06 
0.0 -1.1248 0 2.0 1e-06 
0.0 -1.1247 0 2.0 1e-06 
0.0 -1.1246 0 2.0 1e-06 
0.0 -1.1245 0 2.0 1e-06 
0.0 -1.1244 0 2.0 1e-06 
0.0 -1.1243 0 2.0 1e-06 
0.0 -1.1242 0 2.0 1e-06 
0.0 -1.1241 0 2.0 1e-06 
0.0 -1.124 0 2.0 1e-06 
0.0 -1.1239 0 2.0 1e-06 
0.0 -1.1238 0 2.0 1e-06 
0.0 -1.1237 0 2.0 1e-06 
0.0 -1.1236 0 2.0 1e-06 
0.0 -1.1235 0 2.0 1e-06 
0.0 -1.1234 0 2.0 1e-06 
0.0 -1.1233 0 2.0 1e-06 
0.0 -1.1232 0 2.0 1e-06 
0.0 -1.1231 0 2.0 1e-06 
0.0 -1.123 0 2.0 1e-06 
0.0 -1.1229 0 2.0 1e-06 
0.0 -1.1228 0 2.0 1e-06 
0.0 -1.1227 0 2.0 1e-06 
0.0 -1.1226 0 2.0 1e-06 
0.0 -1.1225 0 2.0 1e-06 
0.0 -1.1224 0 2.0 1e-06 
0.0 -1.1223 0 2.0 1e-06 
0.0 -1.1222 0 2.0 1e-06 
0.0 -1.1221 0 2.0 1e-06 
0.0 -1.122 0 2.0 1e-06 
0.0 -1.1219 0 2.0 1e-06 
0.0 -1.1218 0 2.0 1e-06 
0.0 -1.1217 0 2.0 1e-06 
0.0 -1.1216 0 2.0 1e-06 
0.0 -1.1215 0 2.0 1e-06 
0.0 -1.1214 0 2.0 1e-06 
0.0 -1.1213 0 2.0 1e-06 
0.0 -1.1212 0 2.0 1e-06 
0.0 -1.1211 0 2.0 1e-06 
0.0 -1.121 0 2.0 1e-06 
0.0 -1.1209 0 2.0 1e-06 
0.0 -1.1208 0 2.0 1e-06 
0.0 -1.1207 0 2.0 1e-06 
0.0 -1.1206 0 2.0 1e-06 
0.0 -1.1205 0 2.0 1e-06 
0.0 -1.1204 0 2.0 1e-06 
0.0 -1.1203 0 2.0 1e-06 
0.0 -1.1202 0 2.0 1e-06 
0.0 -1.1201 0 2.0 1e-06 
0.0 -1.12 0 2.0 1e-06 
0.0 -1.1199 0 2.0 1e-06 
0.0 -1.1198 0 2.0 1e-06 
0.0 -1.1197 0 2.0 1e-06 
0.0 -1.1196 0 2.0 1e-06 
0.0 -1.1195 0 2.0 1e-06 
0.0 -1.1194 0 2.0 1e-06 
0.0 -1.1193 0 2.0 1e-06 
0.0 -1.1192 0 2.0 1e-06 
0.0 -1.1191 0 2.0 1e-06 
0.0 -1.119 0 2.0 1e-06 
0.0 -1.1189 0 2.0 1e-06 
0.0 -1.1188 0 2.0 1e-06 
0.0 -1.1187 0 2.0 1e-06 
0.0 -1.1186 0 2.0 1e-06 
0.0 -1.1185 0 2.0 1e-06 
0.0 -1.1184 0 2.0 1e-06 
0.0 -1.1183 0 2.0 1e-06 
0.0 -1.1182 0 2.0 1e-06 
0.0 -1.1181 0 2.0 1e-06 
0.0 -1.118 0 2.0 1e-06 
0.0 -1.1179 0 2.0 1e-06 
0.0 -1.1178 0 2.0 1e-06 
0.0 -1.1177 0 2.0 1e-06 
0.0 -1.1176 0 2.0 1e-06 
0.0 -1.1175 0 2.0 1e-06 
0.0 -1.1174 0 2.0 1e-06 
0.0 -1.1173 0 2.0 1e-06 
0.0 -1.1172 0 2.0 1e-06 
0.0 -1.1171 0 2.0 1e-06 
0.0 -1.117 0 2.0 1e-06 
0.0 -1.1169 0 2.0 1e-06 
0.0 -1.1168 0 2.0 1e-06 
0.0 -1.1167 0 2.0 1e-06 
0.0 -1.1166 0 2.0 1e-06 
0.0 -1.1165 0 2.0 1e-06 
0.0 -1.1164 0 2.0 1e-06 
0.0 -1.1163 0 2.0 1e-06 
0.0 -1.1162 0 2.0 1e-06 
0.0 -1.1161 0 2.0 1e-06 
0.0 -1.116 0 2.0 1e-06 
0.0 -1.1159 0 2.0 1e-06 
0.0 -1.1158 0 2.0 1e-06 
0.0 -1.1157 0 2.0 1e-06 
0.0 -1.1156 0 2.0 1e-06 
0.0 -1.1155 0 2.0 1e-06 
0.0 -1.1154 0 2.0 1e-06 
0.0 -1.1153 0 2.0 1e-06 
0.0 -1.1152 0 2.0 1e-06 
0.0 -1.1151 0 2.0 1e-06 
0.0 -1.115 0 2.0 1e-06 
0.0 -1.1149 0 2.0 1e-06 
0.0 -1.1148 0 2.0 1e-06 
0.0 -1.1147 0 2.0 1e-06 
0.0 -1.1146 0 2.0 1e-06 
0.0 -1.1145 0 2.0 1e-06 
0.0 -1.1144 0 2.0 1e-06 
0.0 -1.1143 0 2.0 1e-06 
0.0 -1.1142 0 2.0 1e-06 
0.0 -1.1141 0 2.0 1e-06 
0.0 -1.114 0 2.0 1e-06 
0.0 -1.1139 0 2.0 1e-06 
0.0 -1.1138 0 2.0 1e-06 
0.0 -1.1137 0 2.0 1e-06 
0.0 -1.1136 0 2.0 1e-06 
0.0 -1.1135 0 2.0 1e-06 
0.0 -1.1134 0 2.0 1e-06 
0.0 -1.1133 0 2.0 1e-06 
0.0 -1.1132 0 2.0 1e-06 
0.0 -1.1131 0 2.0 1e-06 
0.0 -1.113 0 2.0 1e-06 
0.0 -1.1129 0 2.0 1e-06 
0.0 -1.1128 0 2.0 1e-06 
0.0 -1.1127 0 2.0 1e-06 
0.0 -1.1126 0 2.0 1e-06 
0.0 -1.1125 0 2.0 1e-06 
0.0 -1.1124 0 2.0 1e-06 
0.0 -1.1123 0 2.0 1e-06 
0.0 -1.1122 0 2.0 1e-06 
0.0 -1.1121 0 2.0 1e-06 
0.0 -1.112 0 2.0 1e-06 
0.0 -1.1119 0 2.0 1e-06 
0.0 -1.1118 0 2.0 1e-06 
0.0 -1.1117 0 2.0 1e-06 
0.0 -1.1116 0 2.0 1e-06 
0.0 -1.1115 0 2.0 1e-06 
0.0 -1.1114 0 2.0 1e-06 
0.0 -1.1113 0 2.0 1e-06 
0.0 -1.1112 0 2.0 1e-06 
0.0 -1.1111 0 2.0 1e-06 
0.0 -1.111 0 2.0 1e-06 
0.0 -1.1109 0 2.0 1e-06 
0.0 -1.1108 0 2.0 1e-06 
0.0 -1.1107 0 2.0 1e-06 
0.0 -1.1106 0 2.0 1e-06 
0.0 -1.1105 0 2.0 1e-06 
0.0 -1.1104 0 2.0 1e-06 
0.0 -1.1103 0 2.0 1e-06 
0.0 -1.1102 0 2.0 1e-06 
0.0 -1.1101 0 2.0 1e-06 
0.0 -1.11 0 2.0 1e-06 
0.0 -1.1099 0 2.0 1e-06 
0.0 -1.1098 0 2.0 1e-06 
0.0 -1.1097 0 2.0 1e-06 
0.0 -1.1096 0 2.0 1e-06 
0.0 -1.1095 0 2.0 1e-06 
0.0 -1.1094 0 2.0 1e-06 
0.0 -1.1093 0 2.0 1e-06 
0.0 -1.1092 0 2.0 1e-06 
0.0 -1.1091 0 2.0 1e-06 
0.0 -1.109 0 2.0 1e-06 
0.0 -1.1089 0 2.0 1e-06 
0.0 -1.1088 0 2.0 1e-06 
0.0 -1.1087 0 2.0 1e-06 
0.0 -1.1086 0 2.0 1e-06 
0.0 -1.1085 0 2.0 1e-06 
0.0 -1.1084 0 2.0 1e-06 
0.0 -1.1083 0 2.0 1e-06 
0.0 -1.1082 0 2.0 1e-06 
0.0 -1.1081 0 2.0 1e-06 
0.0 -1.108 0 2.0 1e-06 
0.0 -1.1079 0 2.0 1e-06 
0.0 -1.1078 0 2.0 1e-06 
0.0 -1.1077 0 2.0 1e-06 
0.0 -1.1076 0 2.0 1e-06 
0.0 -1.1075 0 2.0 1e-06 
0.0 -1.1074 0 2.0 1e-06 
0.0 -1.1073 0 2.0 1e-06 
0.0 -1.1072 0 2.0 1e-06 
0.0 -1.1071 0 2.0 1e-06 
0.0 -1.107 0 2.0 1e-06 
0.0 -1.1069 0 2.0 1e-06 
0.0 -1.1068 0 2.0 1e-06 
0.0 -1.1067 0 2.0 1e-06 
0.0 -1.1066 0 2.0 1e-06 
0.0 -1.1065 0 2.0 1e-06 
0.0 -1.1064 0 2.0 1e-06 
0.0 -1.1063 0 2.0 1e-06 
0.0 -1.1062 0 2.0 1e-06 
0.0 -1.1061 0 2.0 1e-06 
0.0 -1.106 0 2.0 1e-06 
0.0 -1.1059 0 2.0 1e-06 
0.0 -1.1058 0 2.0 1e-06 
0.0 -1.1057 0 2.0 1e-06 
0.0 -1.1056 0 2.0 1e-06 
0.0 -1.1055 0 2.0 1e-06 
0.0 -1.1054 0 2.0 1e-06 
0.0 -1.1053 0 2.0 1e-06 
0.0 -1.1052 0 2.0 1e-06 
0.0 -1.1051 0 2.0 1e-06 
0.0 -1.105 0 2.0 1e-06 
0.0 -1.1049 0 2.0 1e-06 
0.0 -1.1048 0 2.0 1e-06 
0.0 -1.1047 0 2.0 1e-06 
0.0 -1.1046 0 2.0 1e-06 
0.0 -1.1045 0 2.0 1e-06 
0.0 -1.1044 0 2.0 1e-06 
0.0 -1.1043 0 2.0 1e-06 
0.0 -1.1042 0 2.0 1e-06 
0.0 -1.1041 0 2.0 1e-06 
0.0 -1.104 0 2.0 1e-06 
0.0 -1.1039 0 2.0 1e-06 
0.0 -1.1038 0 2.0 1e-06 
0.0 -1.1037 0 2.0 1e-06 
0.0 -1.1036 0 2.0 1e-06 
0.0 -1.1035 0 2.0 1e-06 
0.0 -1.1034 0 2.0 1e-06 
0.0 -1.1033 0 2.0 1e-06 
0.0 -1.1032 0 2.0 1e-06 
0.0 -1.1031 0 2.0 1e-06 
0.0 -1.103 0 2.0 1e-06 
0.0 -1.1029 0 2.0 1e-06 
0.0 -1.1028 0 2.0 1e-06 
0.0 -1.1027 0 2.0 1e-06 
0.0 -1.1026 0 2.0 1e-06 
0.0 -1.1025 0 2.0 1e-06 
0.0 -1.1024 0 2.0 1e-06 
0.0 -1.1023 0 2.0 1e-06 
0.0 -1.1022 0 2.0 1e-06 
0.0 -1.1021 0 2.0 1e-06 
0.0 -1.102 0 2.0 1e-06 
0.0 -1.1019 0 2.0 1e-06 
0.0 -1.1018 0 2.0 1e-06 
0.0 -1.1017 0 2.0 1e-06 
0.0 -1.1016 0 2.0 1e-06 
0.0 -1.1015 0 2.0 1e-06 
0.0 -1.1014 0 2.0 1e-06 
0.0 -1.1013 0 2.0 1e-06 
0.0 -1.1012 0 2.0 1e-06 
0.0 -1.1011 0 2.0 1e-06 
0.0 -1.101 0 2.0 1e-06 
0.0 -1.1009 0 2.0 1e-06 
0.0 -1.1008 0 2.0 1e-06 
0.0 -1.1007 0 2.0 1e-06 
0.0 -1.1006 0 2.0 1e-06 
0.0 -1.1005 0 2.0 1e-06 
0.0 -1.1004 0 2.0 1e-06 
0.0 -1.1003 0 2.0 1e-06 
0.0 -1.1002 0 2.0 1e-06 
0.0 -1.1001 0 2.0 1e-06 
0.0 -1.1 0 2.0 1e-06 
0.0 -1.0999 0 2.0 1e-06 
0.0 -1.0998 0 2.0 1e-06 
0.0 -1.0997 0 2.0 1e-06 
0.0 -1.0996 0 2.0 1e-06 
0.0 -1.0995 0 2.0 1e-06 
0.0 -1.0994 0 2.0 1e-06 
0.0 -1.0993 0 2.0 1e-06 
0.0 -1.0992 0 2.0 1e-06 
0.0 -1.0991 0 2.0 1e-06 
0.0 -1.099 0 2.0 1e-06 
0.0 -1.0989 0 2.0 1e-06 
0.0 -1.0988 0 2.0 1e-06 
0.0 -1.0987 0 2.0 1e-06 
0.0 -1.0986 0 2.0 1e-06 
0.0 -1.0985 0 2.0 1e-06 
0.0 -1.0984 0 2.0 1e-06 
0.0 -1.0983 0 2.0 1e-06 
0.0 -1.0982 0 2.0 1e-06 
0.0 -1.0981 0 2.0 1e-06 
0.0 -1.098 0 2.0 1e-06 
0.0 -1.0979 0 2.0 1e-06 
0.0 -1.0978 0 2.0 1e-06 
0.0 -1.0977 0 2.0 1e-06 
0.0 -1.0976 0 2.0 1e-06 
0.0 -1.0975 0 2.0 1e-06 
0.0 -1.0974 0 2.0 1e-06 
0.0 -1.0973 0 2.0 1e-06 
0.0 -1.0972 0 2.0 1e-06 
0.0 -1.0971 0 2.0 1e-06 
0.0 -1.097 0 2.0 1e-06 
0.0 -1.0969 0 2.0 1e-06 
0.0 -1.0968 0 2.0 1e-06 
0.0 -1.0967 0 2.0 1e-06 
0.0 -1.0966 0 2.0 1e-06 
0.0 -1.0965 0 2.0 1e-06 
0.0 -1.0964 0 2.0 1e-06 
0.0 -1.0963 0 2.0 1e-06 
0.0 -1.0962 0 2.0 1e-06 
0.0 -1.0961 0 2.0 1e-06 
0.0 -1.096 0 2.0 1e-06 
0.0 -1.0959 0 2.0 1e-06 
0.0 -1.0958 0 2.0 1e-06 
0.0 -1.0957 0 2.0 1e-06 
0.0 -1.0956 0 2.0 1e-06 
0.0 -1.0955 0 2.0 1e-06 
0.0 -1.0954 0 2.0 1e-06 
0.0 -1.0953 0 2.0 1e-06 
0.0 -1.0952 0 2.0 1e-06 
0.0 -1.0951 0 2.0 1e-06 
0.0 -1.095 0 2.0 1e-06 
0.0 -1.0949 0 2.0 1e-06 
0.0 -1.0948 0 2.0 1e-06 
0.0 -1.0947 0 2.0 1e-06 
0.0 -1.0946 0 2.0 1e-06 
0.0 -1.0945 0 2.0 1e-06 
0.0 -1.0944 0 2.0 1e-06 
0.0 -1.0943 0 2.0 1e-06 
0.0 -1.0942 0 2.0 1e-06 
0.0 -1.0941 0 2.0 1e-06 
0.0 -1.094 0 2.0 1e-06 
0.0 -1.0939 0 2.0 1e-06 
0.0 -1.0938 0 2.0 1e-06 
0.0 -1.0937 0 2.0 1e-06 
0.0 -1.0936 0 2.0 1e-06 
0.0 -1.0935 0 2.0 1e-06 
0.0 -1.0934 0 2.0 1e-06 
0.0 -1.0933 0 2.0 1e-06 
0.0 -1.0932 0 2.0 1e-06 
0.0 -1.0931 0 2.0 1e-06 
0.0 -1.093 0 2.0 1e-06 
0.0 -1.0929 0 2.0 1e-06 
0.0 -1.0928 0 2.0 1e-06 
0.0 -1.0927 0 2.0 1e-06 
0.0 -1.0926 0 2.0 1e-06 
0.0 -1.0925 0 2.0 1e-06 
0.0 -1.0924 0 2.0 1e-06 
0.0 -1.0923 0 2.0 1e-06 
0.0 -1.0922 0 2.0 1e-06 
0.0 -1.0921 0 2.0 1e-06 
0.0 -1.092 0 2.0 1e-06 
0.0 -1.0919 0 2.0 1e-06 
0.0 -1.0918 0 2.0 1e-06 
0.0 -1.0917 0 2.0 1e-06 
0.0 -1.0916 0 2.0 1e-06 
0.0 -1.0915 0 2.0 1e-06 
0.0 -1.0914 0 2.0 1e-06 
0.0 -1.0913 0 2.0 1e-06 
0.0 -1.0912 0 2.0 1e-06 
0.0 -1.0911 0 2.0 1e-06 
0.0 -1.091 0 2.0 1e-06 
0.0 -1.0909 0 2.0 1e-06 
0.0 -1.0908 0 2.0 1e-06 
0.0 -1.0907 0 2.0 1e-06 
0.0 -1.0906 0 2.0 1e-06 
0.0 -1.0905 0 2.0 1e-06 
0.0 -1.0904 0 2.0 1e-06 
0.0 -1.0903 0 2.0 1e-06 
0.0 -1.0902 0 2.0 1e-06 
0.0 -1.0901 0 2.0 1e-06 
0.0 -1.09 0 2.0 1e-06 
0.0 -1.0899 0 2.0 1e-06 
0.0 -1.0898 0 2.0 1e-06 
0.0 -1.0897 0 2.0 1e-06 
0.0 -1.0896 0 2.0 1e-06 
0.0 -1.0895 0 2.0 1e-06 
0.0 -1.0894 0 2.0 1e-06 
0.0 -1.0893 0 2.0 1e-06 
0.0 -1.0892 0 2.0 1e-06 
0.0 -1.0891 0 2.0 1e-06 
0.0 -1.089 0 2.0 1e-06 
0.0 -1.0889 0 2.0 1e-06 
0.0 -1.0888 0 2.0 1e-06 
0.0 -1.0887 0 2.0 1e-06 
0.0 -1.0886 0 2.0 1e-06 
0.0 -1.0885 0 2.0 1e-06 
0.0 -1.0884 0 2.0 1e-06 
0.0 -1.0883 0 2.0 1e-06 
0.0 -1.0882 0 2.0 1e-06 
0.0 -1.0881 0 2.0 1e-06 
0.0 -1.088 0 2.0 1e-06 
0.0 -1.0879 0 2.0 1e-06 
0.0 -1.0878 0 2.0 1e-06 
0.0 -1.0877 0 2.0 1e-06 
0.0 -1.0876 0 2.0 1e-06 
0.0 -1.0875 0 2.0 1e-06 
0.0 -1.0874 0 2.0 1e-06 
0.0 -1.0873 0 2.0 1e-06 
0.0 -1.0872 0 2.0 1e-06 
0.0 -1.0871 0 2.0 1e-06 
0.0 -1.087 0 2.0 1e-06 
0.0 -1.0869 0 2.0 1e-06 
0.0 -1.0868 0 2.0 1e-06 
0.0 -1.0867 0 2.0 1e-06 
0.0 -1.0866 0 2.0 1e-06 
0.0 -1.0865 0 2.0 1e-06 
0.0 -1.0864 0 2.0 1e-06 
0.0 -1.0863 0 2.0 1e-06 
0.0 -1.0862 0 2.0 1e-06 
0.0 -1.0861 0 2.0 1e-06 
0.0 -1.086 0 2.0 1e-06 
0.0 -1.0859 0 2.0 1e-06 
0.0 -1.0858 0 2.0 1e-06 
0.0 -1.0857 0 2.0 1e-06 
0.0 -1.0856 0 2.0 1e-06 
0.0 -1.0855 0 2.0 1e-06 
0.0 -1.0854 0 2.0 1e-06 
0.0 -1.0853 0 2.0 1e-06 
0.0 -1.0852 0 2.0 1e-06 
0.0 -1.0851 0 2.0 1e-06 
0.0 -1.085 0 2.0 1e-06 
0.0 -1.0849 0 2.0 1e-06 
0.0 -1.0848 0 2.0 1e-06 
0.0 -1.0847 0 2.0 1e-06 
0.0 -1.0846 0 2.0 1e-06 
0.0 -1.0845 0 2.0 1e-06 
0.0 -1.0844 0 2.0 1e-06 
0.0 -1.0843 0 2.0 1e-06 
0.0 -1.0842 0 2.0 1e-06 
0.0 -1.0841 0 2.0 1e-06 
0.0 -1.084 0 2.0 1e-06 
0.0 -1.0839 0 2.0 1e-06 
0.0 -1.0838 0 2.0 1e-06 
0.0 -1.0837 0 2.0 1e-06 
0.0 -1.0836 0 2.0 1e-06 
0.0 -1.0835 0 2.0 1e-06 
0.0 -1.0834 0 2.0 1e-06 
0.0 -1.0833 0 2.0 1e-06 
0.0 -1.0832 0 2.0 1e-06 
0.0 -1.0831 0 2.0 1e-06 
0.0 -1.083 0 2.0 1e-06 
0.0 -1.0829 0 2.0 1e-06 
0.0 -1.0828 0 2.0 1e-06 
0.0 -1.0827 0 2.0 1e-06 
0.0 -1.0826 0 2.0 1e-06 
0.0 -1.0825 0 2.0 1e-06 
0.0 -1.0824 0 2.0 1e-06 
0.0 -1.0823 0 2.0 1e-06 
0.0 -1.0822 0 2.0 1e-06 
0.0 -1.0821 0 2.0 1e-06 
0.0 -1.082 0 2.0 1e-06 
0.0 -1.0819 0 2.0 1e-06 
0.0 -1.0818 0 2.0 1e-06 
0.0 -1.0817 0 2.0 1e-06 
0.0 -1.0816 0 2.0 1e-06 
0.0 -1.0815 0 2.0 1e-06 
0.0 -1.0814 0 2.0 1e-06 
0.0 -1.0813 0 2.0 1e-06 
0.0 -1.0812 0 2.0 1e-06 
0.0 -1.0811 0 2.0 1e-06 
0.0 -1.081 0 2.0 1e-06 
0.0 -1.0809 0 2.0 1e-06 
0.0 -1.0808 0 2.0 1e-06 
0.0 -1.0807 0 2.0 1e-06 
0.0 -1.0806 0 2.0 1e-06 
0.0 -1.0805 0 2.0 1e-06 
0.0 -1.0804 0 2.0 1e-06 
0.0 -1.0803 0 2.0 1e-06 
0.0 -1.0802 0 2.0 1e-06 
0.0 -1.0801 0 2.0 1e-06 
0.0 -1.08 0 2.0 1e-06 
0.0 -1.0799 0 2.0 1e-06 
0.0 -1.0798 0 2.0 1e-06 
0.0 -1.0797 0 2.0 1e-06 
0.0 -1.0796 0 2.0 1e-06 
0.0 -1.0795 0 2.0 1e-06 
0.0 -1.0794 0 2.0 1e-06 
0.0 -1.0793 0 2.0 1e-06 
0.0 -1.0792 0 2.0 1e-06 
0.0 -1.0791 0 2.0 1e-06 
0.0 -1.079 0 2.0 1e-06 
0.0 -1.0789 0 2.0 1e-06 
0.0 -1.0788 0 2.0 1e-06 
0.0 -1.0787 0 2.0 1e-06 
0.0 -1.0786 0 2.0 1e-06 
0.0 -1.0785 0 2.0 1e-06 
0.0 -1.0784 0 2.0 1e-06 
0.0 -1.0783 0 2.0 1e-06 
0.0 -1.0782 0 2.0 1e-06 
0.0 -1.0781 0 2.0 1e-06 
0.0 -1.078 0 2.0 1e-06 
0.0 -1.0779 0 2.0 1e-06 
0.0 -1.0778 0 2.0 1e-06 
0.0 -1.0777 0 2.0 1e-06 
0.0 -1.0776 0 2.0 1e-06 
0.0 -1.0775 0 2.0 1e-06 
0.0 -1.0774 0 2.0 1e-06 
0.0 -1.0773 0 2.0 1e-06 
0.0 -1.0772 0 2.0 1e-06 
0.0 -1.0771 0 2.0 1e-06 
0.0 -1.077 0 2.0 1e-06 
0.0 -1.0769 0 2.0 1e-06 
0.0 -1.0768 0 2.0 1e-06 
0.0 -1.0767 0 2.0 1e-06 
0.0 -1.0766 0 2.0 1e-06 
0.0 -1.0765 0 2.0 1e-06 
0.0 -1.0764 0 2.0 1e-06 
0.0 -1.0763 0 2.0 1e-06 
0.0 -1.0762 0 2.0 1e-06 
0.0 -1.0761 0 2.0 1e-06 
0.0 -1.076 0 2.0 1e-06 
0.0 -1.0759 0 2.0 1e-06 
0.0 -1.0758 0 2.0 1e-06 
0.0 -1.0757 0 2.0 1e-06 
0.0 -1.0756 0 2.0 1e-06 
0.0 -1.0755 0 2.0 1e-06 
0.0 -1.0754 0 2.0 1e-06 
0.0 -1.0753 0 2.0 1e-06 
0.0 -1.0752 0 2.0 1e-06 
0.0 -1.0751 0 2.0 1e-06 
0.0 -1.075 0 2.0 1e-06 
0.0 -1.0749 0 2.0 1e-06 
0.0 -1.0748 0 2.0 1e-06 
0.0 -1.0747 0 2.0 1e-06 
0.0 -1.0746 0 2.0 1e-06 
0.0 -1.0745 0 2.0 1e-06 
0.0 -1.0744 0 2.0 1e-06 
0.0 -1.0743 0 2.0 1e-06 
0.0 -1.0742 0 2.0 1e-06 
0.0 -1.0741 0 2.0 1e-06 
0.0 -1.074 0 2.0 1e-06 
0.0 -1.0739 0 2.0 1e-06 
0.0 -1.0738 0 2.0 1e-06 
0.0 -1.0737 0 2.0 1e-06 
0.0 -1.0736 0 2.0 1e-06 
0.0 -1.0735 0 2.0 1e-06 
0.0 -1.0734 0 2.0 1e-06 
0.0 -1.0733 0 2.0 1e-06 
0.0 -1.0732 0 2.0 1e-06 
0.0 -1.0731 0 2.0 1e-06 
0.0 -1.073 0 2.0 1e-06 
0.0 -1.0729 0 2.0 1e-06 
0.0 -1.0728 0 2.0 1e-06 
0.0 -1.0727 0 2.0 1e-06 
0.0 -1.0726 0 2.0 1e-06 
0.0 -1.0725 0 2.0 1e-06 
0.0 -1.0724 0 2.0 1e-06 
0.0 -1.0723 0 2.0 1e-06 
0.0 -1.0722 0 2.0 1e-06 
0.0 -1.0721 0 2.0 1e-06 
0.0 -1.072 0 2.0 1e-06 
0.0 -1.0719 0 2.0 1e-06 
0.0 -1.0718 0 2.0 1e-06 
0.0 -1.0717 0 2.0 1e-06 
0.0 -1.0716 0 2.0 1e-06 
0.0 -1.0715 0 2.0 1e-06 
0.0 -1.0714 0 2.0 1e-06 
0.0 -1.0713 0 2.0 1e-06 
0.0 -1.0712 0 2.0 1e-06 
0.0 -1.0711 0 2.0 1e-06 
0.0 -1.071 0 2.0 1e-06 
0.0 -1.0709 0 2.0 1e-06 
0.0 -1.0708 0 2.0 1e-06 
0.0 -1.0707 0 2.0 1e-06 
0.0 -1.0706 0 2.0 1e-06 
0.0 -1.0705 0 2.0 1e-06 
0.0 -1.0704 0 2.0 1e-06 
0.0 -1.0703 0 2.0 1e-06 
0.0 -1.0702 0 2.0 1e-06 
0.0 -1.0701 0 2.0 1e-06 
0.0 -1.07 0 2.0 1e-06 
0.0 -1.0699 0 2.0 1e-06 
0.0 -1.0698 0 2.0 1e-06 
0.0 -1.0697 0 2.0 1e-06 
0.0 -1.0696 0 2.0 1e-06 
0.0 -1.0695 0 2.0 1e-06 
0.0 -1.0694 0 2.0 1e-06 
0.0 -1.0693 0 2.0 1e-06 
0.0 -1.0692 0 2.0 1e-06 
0.0 -1.0691 0 2.0 1e-06 
0.0 -1.069 0 2.0 1e-06 
0.0 -1.0689 0 2.0 1e-06 
0.0 -1.0688 0 2.0 1e-06 
0.0 -1.0687 0 2.0 1e-06 
0.0 -1.0686 0 2.0 1e-06 
0.0 -1.0685 0 2.0 1e-06 
0.0 -1.0684 0 2.0 1e-06 
0.0 -1.0683 0 2.0 1e-06 
0.0 -1.0682 0 2.0 1e-06 
0.0 -1.0681 0 2.0 1e-06 
0.0 -1.068 0 2.0 1e-06 
0.0 -1.0679 0 2.0 1e-06 
0.0 -1.0678 0 2.0 1e-06 
0.0 -1.0677 0 2.0 1e-06 
0.0 -1.0676 0 2.0 1e-06 
0.0 -1.0675 0 2.0 1e-06 
0.0 -1.0674 0 2.0 1e-06 
0.0 -1.0673 0 2.0 1e-06 
0.0 -1.0672 0 2.0 1e-06 
0.0 -1.0671 0 2.0 1e-06 
0.0 -1.067 0 2.0 1e-06 
0.0 -1.0669 0 2.0 1e-06 
0.0 -1.0668 0 2.0 1e-06 
0.0 -1.0667 0 2.0 1e-06 
0.0 -1.0666 0 2.0 1e-06 
0.0 -1.0665 0 2.0 1e-06 
0.0 -1.0664 0 2.0 1e-06 
0.0 -1.0663 0 2.0 1e-06 
0.0 -1.0662 0 2.0 1e-06 
0.0 -1.0661 0 2.0 1e-06 
0.0 -1.066 0 2.0 1e-06 
0.0 -1.0659 0 2.0 1e-06 
0.0 -1.0658 0 2.0 1e-06 
0.0 -1.0657 0 2.0 1e-06 
0.0 -1.0656 0 2.0 1e-06 
0.0 -1.0655 0 2.0 1e-06 
0.0 -1.0654 0 2.0 1e-06 
0.0 -1.0653 0 2.0 1e-06 
0.0 -1.0652 0 2.0 1e-06 
0.0 -1.0651 0 2.0 1e-06 
0.0 -1.065 0 2.0 1e-06 
0.0 -1.0649 0 2.0 1e-06 
0.0 -1.0648 0 2.0 1e-06 
0.0 -1.0647 0 2.0 1e-06 
0.0 -1.0646 0 2.0 1e-06 
0.0 -1.0645 0 2.0 1e-06 
0.0 -1.0644 0 2.0 1e-06 
0.0 -1.0643 0 2.0 1e-06 
0.0 -1.0642 0 2.0 1e-06 
0.0 -1.0641 0 2.0 1e-06 
0.0 -1.064 0 2.0 1e-06 
0.0 -1.0639 0 2.0 1e-06 
0.0 -1.0638 0 2.0 1e-06 
0.0 -1.0637 0 2.0 1e-06 
0.0 -1.0636 0 2.0 1e-06 
0.0 -1.0635 0 2.0 1e-06 
0.0 -1.0634 0 2.0 1e-06 
0.0 -1.0633 0 2.0 1e-06 
0.0 -1.0632 0 2.0 1e-06 
0.0 -1.0631 0 2.0 1e-06 
0.0 -1.063 0 2.0 1e-06 
0.0 -1.0629 0 2.0 1e-06 
0.0 -1.0628 0 2.0 1e-06 
0.0 -1.0627 0 2.0 1e-06 
0.0 -1.0626 0 2.0 1e-06 
0.0 -1.0625 0 2.0 1e-06 
0.0 -1.0624 0 2.0 1e-06 
0.0 -1.0623 0 2.0 1e-06 
0.0 -1.0622 0 2.0 1e-06 
0.0 -1.0621 0 2.0 1e-06 
0.0 -1.062 0 2.0 1e-06 
0.0 -1.0619 0 2.0 1e-06 
0.0 -1.0618 0 2.0 1e-06 
0.0 -1.0617 0 2.0 1e-06 
0.0 -1.0616 0 2.0 1e-06 
0.0 -1.0615 0 2.0 1e-06 
0.0 -1.0614 0 2.0 1e-06 
0.0 -1.0613 0 2.0 1e-06 
0.0 -1.0612 0 2.0 1e-06 
0.0 -1.0611 0 2.0 1e-06 
0.0 -1.061 0 2.0 1e-06 
0.0 -1.0609 0 2.0 1e-06 
0.0 -1.0608 0 2.0 1e-06 
0.0 -1.0607 0 2.0 1e-06 
0.0 -1.0606 0 2.0 1e-06 
0.0 -1.0605 0 2.0 1e-06 
0.0 -1.0604 0 2.0 1e-06 
0.0 -1.0603 0 2.0 1e-06 
0.0 -1.0602 0 2.0 1e-06 
0.0 -1.0601 0 2.0 1e-06 
0.0 -1.06 0 2.0 1e-06 
0.0 -1.0599 0 2.0 1e-06 
0.0 -1.0598 0 2.0 1e-06 
0.0 -1.0597 0 2.0 1e-06 
0.0 -1.0596 0 2.0 1e-06 
0.0 -1.0595 0 2.0 1e-06 
0.0 -1.0594 0 2.0 1e-06 
0.0 -1.0593 0 2.0 1e-06 
0.0 -1.0592 0 2.0 1e-06 
0.0 -1.0591 0 2.0 1e-06 
0.0 -1.059 0 2.0 1e-06 
0.0 -1.0589 0 2.0 1e-06 
0.0 -1.0588 0 2.0 1e-06 
0.0 -1.0587 0 2.0 1e-06 
0.0 -1.0586 0 2.0 1e-06 
0.0 -1.0585 0 2.0 1e-06 
0.0 -1.0584 0 2.0 1e-06 
0.0 -1.0583 0 2.0 1e-06 
0.0 -1.0582 0 2.0 1e-06 
0.0 -1.0581 0 2.0 1e-06 
0.0 -1.058 0 2.0 1e-06 
0.0 -1.0579 0 2.0 1e-06 
0.0 -1.0578 0 2.0 1e-06 
0.0 -1.0577 0 2.0 1e-06 
0.0 -1.0576 0 2.0 1e-06 
0.0 -1.0575 0 2.0 1e-06 
0.0 -1.0574 0 2.0 1e-06 
0.0 -1.0573 0 2.0 1e-06 
0.0 -1.0572 0 2.0 1e-06 
0.0 -1.0571 0 2.0 1e-06 
0.0 -1.057 0 2.0 1e-06 
0.0 -1.0569 0 2.0 1e-06 
0.0 -1.0568 0 2.0 1e-06 
0.0 -1.0567 0 2.0 1e-06 
0.0 -1.0566 0 2.0 1e-06 
0.0 -1.0565 0 2.0 1e-06 
0.0 -1.0564 0 2.0 1e-06 
0.0 -1.0563 0 2.0 1e-06 
0.0 -1.0562 0 2.0 1e-06 
0.0 -1.0561 0 2.0 1e-06 
0.0 -1.056 0 2.0 1e-06 
0.0 -1.0559 0 2.0 1e-06 
0.0 -1.0558 0 2.0 1e-06 
0.0 -1.0557 0 2.0 1e-06 
0.0 -1.0556 0 2.0 1e-06 
0.0 -1.0555 0 2.0 1e-06 
0.0 -1.0554 0 2.0 1e-06 
0.0 -1.0553 0 2.0 1e-06 
0.0 -1.0552 0 2.0 1e-06 
0.0 -1.0551 0 2.0 1e-06 
0.0 -1.055 0 2.0 1e-06 
0.0 -1.0549 0 2.0 1e-06 
0.0 -1.0548 0 2.0 1e-06 
0.0 -1.0547 0 2.0 1e-06 
0.0 -1.0546 0 2.0 1e-06 
0.0 -1.0545 0 2.0 1e-06 
0.0 -1.0544 0 2.0 1e-06 
0.0 -1.0543 0 2.0 1e-06 
0.0 -1.0542 0 2.0 1e-06 
0.0 -1.0541 0 2.0 1e-06 
0.0 -1.054 0 2.0 1e-06 
0.0 -1.0539 0 2.0 1e-06 
0.0 -1.0538 0 2.0 1e-06 
0.0 -1.0537 0 2.0 1e-06 
0.0 -1.0536 0 2.0 1e-06 
0.0 -1.0535 0 2.0 1e-06 
0.0 -1.0534 0 2.0 1e-06 
0.0 -1.0533 0 2.0 1e-06 
0.0 -1.0532 0 2.0 1e-06 
0.0 -1.0531 0 2.0 1e-06 
0.0 -1.053 0 2.0 1e-06 
0.0 -1.0529 0 2.0 1e-06 
0.0 -1.0528 0 2.0 1e-06 
0.0 -1.0527 0 2.0 1e-06 
0.0 -1.0526 0 2.0 1e-06 
0.0 -1.0525 0 2.0 1e-06 
0.0 -1.0524 0 2.0 1e-06 
0.0 -1.0523 0 2.0 1e-06 
0.0 -1.0522 0 2.0 1e-06 
0.0 -1.0521 0 2.0 1e-06 
0.0 -1.052 0 2.0 1e-06 
0.0 -1.0519 0 2.0 1e-06 
0.0 -1.0518 0 2.0 1e-06 
0.0 -1.0517 0 2.0 1e-06 
0.0 -1.0516 0 2.0 1e-06 
0.0 -1.0515 0 2.0 1e-06 
0.0 -1.0514 0 2.0 1e-06 
0.0 -1.0513 0 2.0 1e-06 
0.0 -1.0512 0 2.0 1e-06 
0.0 -1.0511 0 2.0 1e-06 
0.0 -1.051 0 2.0 1e-06 
0.0 -1.0509 0 2.0 1e-06 
0.0 -1.0508 0 2.0 1e-06 
0.0 -1.0507 0 2.0 1e-06 
0.0 -1.0506 0 2.0 1e-06 
0.0 -1.0505 0 2.0 1e-06 
0.0 -1.0504 0 2.0 1e-06 
0.0 -1.0503 0 2.0 1e-06 
0.0 -1.0502 0 2.0 1e-06 
0.0 -1.0501 0 2.0 1e-06 
0.0 -1.05 0 2.0 1e-06 
0.0 -1.0499 0 2.0 1e-06 
0.0 -1.0498 0 2.0 1e-06 
0.0 -1.0497 0 2.0 1e-06 
0.0 -1.0496 0 2.0 1e-06 
0.0 -1.0495 0 2.0 1e-06 
0.0 -1.0494 0 2.0 1e-06 
0.0 -1.0493 0 2.0 1e-06 
0.0 -1.0492 0 2.0 1e-06 
0.0 -1.0491 0 2.0 1e-06 
0.0 -1.049 0 2.0 1e-06 
0.0 -1.0489 0 2.0 1e-06 
0.0 -1.0488 0 2.0 1e-06 
0.0 -1.0487 0 2.0 1e-06 
0.0 -1.0486 0 2.0 1e-06 
0.0 -1.0485 0 2.0 1e-06 
0.0 -1.0484 0 2.0 1e-06 
0.0 -1.0483 0 2.0 1e-06 
0.0 -1.0482 0 2.0 1e-06 
0.0 -1.0481 0 2.0 1e-06 
0.0 -1.048 0 2.0 1e-06 
0.0 -1.0479 0 2.0 1e-06 
0.0 -1.0478 0 2.0 1e-06 
0.0 -1.0477 0 2.0 1e-06 
0.0 -1.0476 0 2.0 1e-06 
0.0 -1.0475 0 2.0 1e-06 
0.0 -1.0474 0 2.0 1e-06 
0.0 -1.0473 0 2.0 1e-06 
0.0 -1.0472 0 2.0 1e-06 
0.0 -1.0471 0 2.0 1e-06 
0.0 -1.047 0 2.0 1e-06 
0.0 -1.0469 0 2.0 1e-06 
0.0 -1.0468 0 2.0 1e-06 
0.0 -1.0467 0 2.0 1e-06 
0.0 -1.0466 0 2.0 1e-06 
0.0 -1.0465 0 2.0 1e-06 
0.0 -1.0464 0 2.0 1e-06 
0.0 -1.0463 0 2.0 1e-06 
0.0 -1.0462 0 2.0 1e-06 
0.0 -1.0461 0 2.0 1e-06 
0.0 -1.046 0 2.0 1e-06 
0.0 -1.0459 0 2.0 1e-06 
0.0 -1.0458 0 2.0 1e-06 
0.0 -1.0457 0 2.0 1e-06 
0.0 -1.0456 0 2.0 1e-06 
0.0 -1.0455 0 2.0 1e-06 
0.0 -1.0454 0 2.0 1e-06 
0.0 -1.0453 0 2.0 1e-06 
0.0 -1.0452 0 2.0 1e-06 
0.0 -1.0451 0 2.0 1e-06 
0.0 -1.045 0 2.0 1e-06 
0.0 -1.0449 0 2.0 1e-06 
0.0 -1.0448 0 2.0 1e-06 
0.0 -1.0447 0 2.0 1e-06 
0.0 -1.0446 0 2.0 1e-06 
0.0 -1.0445 0 2.0 1e-06 
0.0 -1.0444 0 2.0 1e-06 
0.0 -1.0443 0 2.0 1e-06 
0.0 -1.0442 0 2.0 1e-06 
0.0 -1.0441 0 2.0 1e-06 
0.0 -1.044 0 2.0 1e-06 
0.0 -1.0439 0 2.0 1e-06 
0.0 -1.0438 0 2.0 1e-06 
0.0 -1.0437 0 2.0 1e-06 
0.0 -1.0436 0 2.0 1e-06 
0.0 -1.0435 0 2.0 1e-06 
0.0 -1.0434 0 2.0 1e-06 
0.0 -1.0433 0 2.0 1e-06 
0.0 -1.0432 0 2.0 1e-06 
0.0 -1.0431 0 2.0 1e-06 
0.0 -1.043 0 2.0 1e-06 
0.0 -1.0429 0 2.0 1e-06 
0.0 -1.0428 0 2.0 1e-06 
0.0 -1.0427 0 2.0 1e-06 
0.0 -1.0426 0 2.0 1e-06 
0.0 -1.0425 0 2.0 1e-06 
0.0 -1.0424 0 2.0 1e-06 
0.0 -1.0423 0 2.0 1e-06 
0.0 -1.0422 0 2.0 1e-06 
0.0 -1.0421 0 2.0 1e-06 
0.0 -1.042 0 2.0 1e-06 
0.0 -1.0419 0 2.0 1e-06 
0.0 -1.0418 0 2.0 1e-06 
0.0 -1.0417 0 2.0 1e-06 
0.0 -1.0416 0 2.0 1e-06 
0.0 -1.0415 0 2.0 1e-06 
0.0 -1.0414 0 2.0 1e-06 
0.0 -1.0413 0 2.0 1e-06 
0.0 -1.0412 0 2.0 1e-06 
0.0 -1.0411 0 2.0 1e-06 
0.0 -1.041 0 2.0 1e-06 
0.0 -1.0409 0 2.0 1e-06 
0.0 -1.0408 0 2.0 1e-06 
0.0 -1.0407 0 2.0 1e-06 
0.0 -1.0406 0 2.0 1e-06 
0.0 -1.0405 0 2.0 1e-06 
0.0 -1.0404 0 2.0 1e-06 
0.0 -1.0403 0 2.0 1e-06 
0.0 -1.0402 0 2.0 1e-06 
0.0 -1.0401 0 2.0 1e-06 
0.0 -1.04 0 2.0 1e-06 
0.0 -1.0399 0 2.0 1e-06 
0.0 -1.0398 0 2.0 1e-06 
0.0 -1.0397 0 2.0 1e-06 
0.0 -1.0396 0 2.0 1e-06 
0.0 -1.0395 0 2.0 1e-06 
0.0 -1.0394 0 2.0 1e-06 
0.0 -1.0393 0 2.0 1e-06 
0.0 -1.0392 0 2.0 1e-06 
0.0 -1.0391 0 2.0 1e-06 
0.0 -1.039 0 2.0 1e-06 
0.0 -1.0389 0 2.0 1e-06 
0.0 -1.0388 0 2.0 1e-06 
0.0 -1.0387 0 2.0 1e-06 
0.0 -1.0386 0 2.0 1e-06 
0.0 -1.0385 0 2.0 1e-06 
0.0 -1.0384 0 2.0 1e-06 
0.0 -1.0383 0 2.0 1e-06 
0.0 -1.0382 0 2.0 1e-06 
0.0 -1.0381 0 2.0 1e-06 
0.0 -1.038 0 2.0 1e-06 
0.0 -1.0379 0 2.0 1e-06 
0.0 -1.0378 0 2.0 1e-06 
0.0 -1.0377 0 2.0 1e-06 
0.0 -1.0376 0 2.0 1e-06 
0.0 -1.0375 0 2.0 1e-06 
0.0 -1.0374 0 2.0 1e-06 
0.0 -1.0373 0 2.0 1e-06 
0.0 -1.0372 0 2.0 1e-06 
0.0 -1.0371 0 2.0 1e-06 
0.0 -1.037 0 2.0 1e-06 
0.0 -1.0369 0 2.0 1e-06 
0.0 -1.0368 0 2.0 1e-06 
0.0 -1.0367 0 2.0 1e-06 
0.0 -1.0366 0 2.0 1e-06 
0.0 -1.0365 0 2.0 1e-06 
0.0 -1.0364 0 2.0 1e-06 
0.0 -1.0363 0 2.0 1e-06 
0.0 -1.0362 0 2.0 1e-06 
0.0 -1.0361 0 2.0 1e-06 
0.0 -1.036 0 2.0 1e-06 
0.0 -1.0359 0 2.0 1e-06 
0.0 -1.0358 0 2.0 1e-06 
0.0 -1.0357 0 2.0 1e-06 
0.0 -1.0356 0 2.0 1e-06 
0.0 -1.0355 0 2.0 1e-06 
0.0 -1.0354 0 2.0 1e-06 
0.0 -1.0353 0 2.0 1e-06 
0.0 -1.0352 0 2.0 1e-06 
0.0 -1.0351 0 2.0 1e-06 
0.0 -1.035 0 2.0 1e-06 
0.0 -1.0349 0 2.0 1e-06 
0.0 -1.0348 0 2.0 1e-06 
0.0 -1.0347 0 2.0 1e-06 
0.0 -1.0346 0 2.0 1e-06 
0.0 -1.0345 0 2.0 1e-06 
0.0 -1.0344 0 2.0 1e-06 
0.0 -1.0343 0 2.0 1e-06 
0.0 -1.0342 0 2.0 1e-06 
0.0 -1.0341 0 2.0 1e-06 
0.0 -1.034 0 2.0 1e-06 
0.0 -1.0339 0 2.0 1e-06 
0.0 -1.0338 0 2.0 1e-06 
0.0 -1.0337 0 2.0 1e-06 
0.0 -1.0336 0 2.0 1e-06 
0.0 -1.0335 0 2.0 1e-06 
0.0 -1.0334 0 2.0 1e-06 
0.0 -1.0333 0 2.0 1e-06 
0.0 -1.0332 0 2.0 1e-06 
0.0 -1.0331 0 2.0 1e-06 
0.0 -1.033 0 2.0 1e-06 
0.0 -1.0329 0 2.0 1e-06 
0.0 -1.0328 0 2.0 1e-06 
0.0 -1.0327 0 2.0 1e-06 
0.0 -1.0326 0 2.0 1e-06 
0.0 -1.0325 0 2.0 1e-06 
0.0 -1.0324 0 2.0 1e-06 
0.0 -1.0323 0 2.0 1e-06 
0.0 -1.0322 0 2.0 1e-06 
0.0 -1.0321 0 2.0 1e-06 
0.0 -1.032 0 2.0 1e-06 
0.0 -1.0319 0 2.0 1e-06 
0.0 -1.0318 0 2.0 1e-06 
0.0 -1.0317 0 2.0 1e-06 
0.0 -1.0316 0 2.0 1e-06 
0.0 -1.0315 0 2.0 1e-06 
0.0 -1.0314 0 2.0 1e-06 
0.0 -1.0313 0 2.0 1e-06 
0.0 -1.0312 0 2.0 1e-06 
0.0 -1.0311 0 2.0 1e-06 
0.0 -1.031 0 2.0 1e-06 
0.0 -1.0309 0 2.0 1e-06 
0.0 -1.0308 0 2.0 1e-06 
0.0 -1.0307 0 2.0 1e-06 
0.0 -1.0306 0 2.0 1e-06 
0.0 -1.0305 0 2.0 1e-06 
0.0 -1.0304 0 2.0 1e-06 
0.0 -1.0303 0 2.0 1e-06 
0.0 -1.0302 0 2.0 1e-06 
0.0 -1.0301 0 2.0 1e-06 
0.0 -1.03 0 2.0 1e-06 
0.0 -1.0299 0 2.0 1e-06 
0.0 -1.0298 0 2.0 1e-06 
0.0 -1.0297 0 2.0 1e-06 
0.0 -1.0296 0 2.0 1e-06 
0.0 -1.0295 0 2.0 1e-06 
0.0 -1.0294 0 2.0 1e-06 
0.0 -1.0293 0 2.0 1e-06 
0.0 -1.0292 0 2.0 1e-06 
0.0 -1.0291 0 2.0 1e-06 
0.0 -1.029 0 2.0 1e-06 
0.0 -1.0289 0 2.0 1e-06 
0.0 -1.0288 0 2.0 1e-06 
0.0 -1.0287 0 2.0 1e-06 
0.0 -1.0286 0 2.0 1e-06 
0.0 -1.0285 0 2.0 1e-06 
0.0 -1.0284 0 2.0 1e-06 
0.0 -1.0283 0 2.0 1e-06 
0.0 -1.0282 0 2.0 1e-06 
0.0 -1.0281 0 2.0 1e-06 
0.0 -1.028 0 2.0 1e-06 
0.0 -1.0279 0 2.0 1e-06 
0.0 -1.0278 0 2.0 1e-06 
0.0 -1.0277 0 2.0 1e-06 
0.0 -1.0276 0 2.0 1e-06 
0.0 -1.0275 0 2.0 1e-06 
0.0 -1.0274 0 2.0 1e-06 
0.0 -1.0273 0 2.0 1e-06 
0.0 -1.0272 0 2.0 1e-06 
0.0 -1.0271 0 2.0 1e-06 
0.0 -1.027 0 2.0 1e-06 
0.0 -1.0269 0 2.0 1e-06 
0.0 -1.0268 0 2.0 1e-06 
0.0 -1.0267 0 2.0 1e-06 
0.0 -1.0266 0 2.0 1e-06 
0.0 -1.0265 0 2.0 1e-06 
0.0 -1.0264 0 2.0 1e-06 
0.0 -1.0263 0 2.0 1e-06 
0.0 -1.0262 0 2.0 1e-06 
0.0 -1.0261 0 2.0 1e-06 
0.0 -1.026 0 2.0 1e-06 
0.0 -1.0259 0 2.0 1e-06 
0.0 -1.0258 0 2.0 1e-06 
0.0 -1.0257 0 2.0 1e-06 
0.0 -1.0256 0 2.0 1e-06 
0.0 -1.0255 0 2.0 1e-06 
0.0 -1.0254 0 2.0 1e-06 
0.0 -1.0253 0 2.0 1e-06 
0.0 -1.0252 0 2.0 1e-06 
0.0 -1.0251 0 2.0 1e-06 
0.0 -1.025 0 2.0 1e-06 
0.0 -1.0249 0 2.0 1e-06 
0.0 -1.0248 0 2.0 1e-06 
0.0 -1.0247 0 2.0 1e-06 
0.0 -1.0246 0 2.0 1e-06 
0.0 -1.0245 0 2.0 1e-06 
0.0 -1.0244 0 2.0 1e-06 
0.0 -1.0243 0 2.0 1e-06 
0.0 -1.0242 0 2.0 1e-06 
0.0 -1.0241 0 2.0 1e-06 
0.0 -1.024 0 2.0 1e-06 
0.0 -1.0239 0 2.0 1e-06 
0.0 -1.0238 0 2.0 1e-06 
0.0 -1.0237 0 2.0 1e-06 
0.0 -1.0236 0 2.0 1e-06 
0.0 -1.0235 0 2.0 1e-06 
0.0 -1.0234 0 2.0 1e-06 
0.0 -1.0233 0 2.0 1e-06 
0.0 -1.0232 0 2.0 1e-06 
0.0 -1.0231 0 2.0 1e-06 
0.0 -1.023 0 2.0 1e-06 
0.0 -1.0229 0 2.0 1e-06 
0.0 -1.0228 0 2.0 1e-06 
0.0 -1.0227 0 2.0 1e-06 
0.0 -1.0226 0 2.0 1e-06 
0.0 -1.0225 0 2.0 1e-06 
0.0 -1.0224 0 2.0 1e-06 
0.0 -1.0223 0 2.0 1e-06 
0.0 -1.0222 0 2.0 1e-06 
0.0 -1.0221 0 2.0 1e-06 
0.0 -1.022 0 2.0 1e-06 
0.0 -1.0219 0 2.0 1e-06 
0.0 -1.0218 0 2.0 1e-06 
0.0 -1.0217 0 2.0 1e-06 
0.0 -1.0216 0 2.0 1e-06 
0.0 -1.0215 0 2.0 1e-06 
0.0 -1.0214 0 2.0 1e-06 
0.0 -1.0213 0 2.0 1e-06 
0.0 -1.0212 0 2.0 1e-06 
0.0 -1.0211 0 2.0 1e-06 
0.0 -1.021 0 2.0 1e-06 
0.0 -1.0209 0 2.0 1e-06 
0.0 -1.0208 0 2.0 1e-06 
0.0 -1.0207 0 2.0 1e-06 
0.0 -1.0206 0 2.0 1e-06 
0.0 -1.0205 0 2.0 1e-06 
0.0 -1.0204 0 2.0 1e-06 
0.0 -1.0203 0 2.0 1e-06 
0.0 -1.0202 0 2.0 1e-06 
0.0 -1.0201 0 2.0 1e-06 
0.0 -1.02 0 2.0 1e-06 
0.0 -1.0199 0 2.0 1e-06 
0.0 -1.0198 0 2.0 1e-06 
0.0 -1.0197 0 2.0 1e-06 
0.0 -1.0196 0 2.0 1e-06 
0.0 -1.0195 0 2.0 1e-06 
0.0 -1.0194 0 2.0 1e-06 
0.0 -1.0193 0 2.0 1e-06 
0.0 -1.0192 0 2.0 1e-06 
0.0 -1.0191 0 2.0 1e-06 
0.0 -1.019 0 2.0 1e-06 
0.0 -1.0189 0 2.0 1e-06 
0.0 -1.0188 0 2.0 1e-06 
0.0 -1.0187 0 2.0 1e-06 
0.0 -1.0186 0 2.0 1e-06 
0.0 -1.0185 0 2.0 1e-06 
0.0 -1.0184 0 2.0 1e-06 
0.0 -1.0183 0 2.0 1e-06 
0.0 -1.0182 0 2.0 1e-06 
0.0 -1.0181 0 2.0 1e-06 
0.0 -1.018 0 2.0 1e-06 
0.0 -1.0179 0 2.0 1e-06 
0.0 -1.0178 0 2.0 1e-06 
0.0 -1.0177 0 2.0 1e-06 
0.0 -1.0176 0 2.0 1e-06 
0.0 -1.0175 0 2.0 1e-06 
0.0 -1.0174 0 2.0 1e-06 
0.0 -1.0173 0 2.0 1e-06 
0.0 -1.0172 0 2.0 1e-06 
0.0 -1.0171 0 2.0 1e-06 
0.0 -1.017 0 2.0 1e-06 
0.0 -1.0169 0 2.0 1e-06 
0.0 -1.0168 0 2.0 1e-06 
0.0 -1.0167 0 2.0 1e-06 
0.0 -1.0166 0 2.0 1e-06 
0.0 -1.0165 0 2.0 1e-06 
0.0 -1.0164 0 2.0 1e-06 
0.0 -1.0163 0 2.0 1e-06 
0.0 -1.0162 0 2.0 1e-06 
0.0 -1.0161 0 2.0 1e-06 
0.0 -1.016 0 2.0 1e-06 
0.0 -1.0159 0 2.0 1e-06 
0.0 -1.0158 0 2.0 1e-06 
0.0 -1.0157 0 2.0 1e-06 
0.0 -1.0156 0 2.0 1e-06 
0.0 -1.0155 0 2.0 1e-06 
0.0 -1.0154 0 2.0 1e-06 
0.0 -1.0153 0 2.0 1e-06 
0.0 -1.0152 0 2.0 1e-06 
0.0 -1.0151 0 2.0 1e-06 
0.0 -1.015 0 2.0 1e-06 
0.0 -1.0149 0 2.0 1e-06 
0.0 -1.0148 0 2.0 1e-06 
0.0 -1.0147 0 2.0 1e-06 
0.0 -1.0146 0 2.0 1e-06 
0.0 -1.0145 0 2.0 1e-06 
0.0 -1.0144 0 2.0 1e-06 
0.0 -1.0143 0 2.0 1e-06 
0.0 -1.0142 0 2.0 1e-06 
0.0 -1.0141 0 2.0 1e-06 
0.0 -1.014 0 2.0 1e-06 
0.0 -1.0139 0 2.0 1e-06 
0.0 -1.0138 0 2.0 1e-06 
0.0 -1.0137 0 2.0 1e-06 
0.0 -1.0136 0 2.0 1e-06 
0.0 -1.0135 0 2.0 1e-06 
0.0 -1.0134 0 2.0 1e-06 
0.0 -1.0133 0 2.0 1e-06 
0.0 -1.0132 0 2.0 1e-06 
0.0 -1.0131 0 2.0 1e-06 
0.0 -1.013 0 2.0 1e-06 
0.0 -1.0129 0 2.0 1e-06 
0.0 -1.0128 0 2.0 1e-06 
0.0 -1.0127 0 2.0 1e-06 
0.0 -1.0126 0 2.0 1e-06 
0.0 -1.0125 0 2.0 1e-06 
0.0 -1.0124 0 2.0 1e-06 
0.0 -1.0123 0 2.0 1e-06 
0.0 -1.0122 0 2.0 1e-06 
0.0 -1.0121 0 2.0 1e-06 
0.0 -1.012 0 2.0 1e-06 
0.0 -1.0119 0 2.0 1e-06 
0.0 -1.0118 0 2.0 1e-06 
0.0 -1.0117 0 2.0 1e-06 
0.0 -1.0116 0 2.0 1e-06 
0.0 -1.0115 0 2.0 1e-06 
0.0 -1.0114 0 2.0 1e-06 
0.0 -1.0113 0 2.0 1e-06 
0.0 -1.0112 0 2.0 1e-06 
0.0 -1.0111 0 2.0 1e-06 
0.0 -1.011 0 2.0 1e-06 
0.0 -1.0109 0 2.0 1e-06 
0.0 -1.0108 0 2.0 1e-06 
0.0 -1.0107 0 2.0 1e-06 
0.0 -1.0106 0 2.0 1e-06 
0.0 -1.0105 0 2.0 1e-06 
0.0 -1.0104 0 2.0 1e-06 
0.0 -1.0103 0 2.0 1e-06 
0.0 -1.0102 0 2.0 1e-06 
0.0 -1.0101 0 2.0 1e-06 
0.0 -1.01 0 2.0 1e-06 
0.0 -1.0099 0 2.0 1e-06 
0.0 -1.0098 0 2.0 1e-06 
0.0 -1.0097 0 2.0 1e-06 
0.0 -1.0096 0 2.0 1e-06 
0.0 -1.0095 0 2.0 1e-06 
0.0 -1.0094 0 2.0 1e-06 
0.0 -1.0093 0 2.0 1e-06 
0.0 -1.0092 0 2.0 1e-06 
0.0 -1.0091 0 2.0 1e-06 
0.0 -1.009 0 2.0 1e-06 
0.0 -1.0089 0 2.0 1e-06 
0.0 -1.0088 0 2.0 1e-06 
0.0 -1.0087 0 2.0 1e-06 
0.0 -1.0086 0 2.0 1e-06 
0.0 -1.0085 0 2.0 1e-06 
0.0 -1.0084 0 2.0 1e-06 
0.0 -1.0083 0 2.0 1e-06 
0.0 -1.0082 0 2.0 1e-06 
0.0 -1.0081 0 2.0 1e-06 
0.0 -1.008 0 2.0 1e-06 
0.0 -1.0079 0 2.0 1e-06 
0.0 -1.0078 0 2.0 1e-06 
0.0 -1.0077 0 2.0 1e-06 
0.0 -1.0076 0 2.0 1e-06 
0.0 -1.0075 0 2.0 1e-06 
0.0 -1.0074 0 2.0 1e-06 
0.0 -1.0073 0 2.0 1e-06 
0.0 -1.0072 0 2.0 1e-06 
0.0 -1.0071 0 2.0 1e-06 
0.0 -1.007 0 2.0 1e-06 
0.0 -1.0069 0 2.0 1e-06 
0.0 -1.0068 0 2.0 1e-06 
0.0 -1.0067 0 2.0 1e-06 
0.0 -1.0066 0 2.0 1e-06 
0.0 -1.0065 0 2.0 1e-06 
0.0 -1.0064 0 2.0 1e-06 
0.0 -1.0063 0 2.0 1e-06 
0.0 -1.0062 0 2.0 1e-06 
0.0 -1.0061 0 2.0 1e-06 
0.0 -1.006 0 2.0 1e-06 
0.0 -1.0059 0 2.0 1e-06 
0.0 -1.0058 0 2.0 1e-06 
0.0 -1.0057 0 2.0 1e-06 
0.0 -1.0056 0 2.0 1e-06 
0.0 -1.0055 0 2.0 1e-06 
0.0 -1.0054 0 2.0 1e-06 
0.0 -1.0053 0 2.0 1e-06 
0.0 -1.0052 0 2.0 1e-06 
0.0 -1.0051 0 2.0 1e-06 
0.0 -1.005 0 2.0 1e-06 
0.0 -1.0049 0 2.0 1e-06 
0.0 -1.0048 0 2.0 1e-06 
0.0 -1.0047 0 2.0 1e-06 
0.0 -1.0046 0 2.0 1e-06 
0.0 -1.0045 0 2.0 1e-06 
0.0 -1.0044 0 2.0 1e-06 
0.0 -1.0043 0 2.0 1e-06 
0.0 -1.0042 0 2.0 1e-06 
0.0 -1.0041 0 2.0 1e-06 
0.0 -1.004 0 2.0 1e-06 
0.0 -1.0039 0 2.0 1e-06 
0.0 -1.0038 0 2.0 1e-06 
0.0 -1.0037 0 2.0 1e-06 
0.0 -1.0036 0 2.0 1e-06 
0.0 -1.0035 0 2.0 1e-06 
0.0 -1.0034 0 2.0 1e-06 
0.0 -1.0033 0 2.0 1e-06 
0.0 -1.0032 0 2.0 1e-06 
0.0 -1.0031 0 2.0 1e-06 
0.0 -1.003 0 2.0 1e-06 
0.0 -1.0029 0 2.0 1e-06 
0.0 -1.0028 0 2.0 1e-06 
0.0 -1.0027 0 2.0 1e-06 
0.0 -1.0026 0 2.0 1e-06 
0.0 -1.0025 0 2.0 1e-06 
0.0 -1.0024 0 2.0 1e-06 
0.0 -1.0023 0 2.0 1e-06 
0.0 -1.0022 0 2.0 1e-06 
0.0 -1.0021 0 2.0 1e-06 
0.0 -1.002 0 2.0 1e-06 
0.0 -1.0019 0 2.0 1e-06 
0.0 -1.0018 0 2.0 1e-06 
0.0 -1.0017 0 2.0 1e-06 
0.0 -1.0016 0 2.0 1e-06 
0.0 -1.0015 0 2.0 1e-06 
0.0 -1.0014 0 2.0 1e-06 
0.0 -1.0013 0 2.0 1e-06 
0.0 -1.0012 0 2.0 1e-06 
0.0 -1.0011 0 2.0 1e-06 
0.0 -1.001 0 2.0 1e-06 
0.0 -1.0009 0 2.0 1e-06 
0.0 -1.0008 0 2.0 1e-06 
0.0 -1.0007 0 2.0 1e-06 
0.0 -1.0006 0 2.0 1e-06 
0.0 -1.0005 0 2.0 1e-06 
0.0 -1.0004 0 2.0 1e-06 
0.0 -1.0003 0 2.0 1e-06 
0.0 -1.0002 0 2.0 1e-06 
0.0 -1.0001 0 2.0 1e-06 
0.0 -1.0 0 2.0 1e-06 
0.0 -0.9999 0 2.0 1e-06 
0.0 -0.9998 0 2.0 1e-06 
0.0 -0.9997 0 2.0 1e-06 
0.0 -0.9996 0 2.0 1e-06 
0.0 -0.9995 0 2.0 1e-06 
0.0 -0.9994 0 2.0 1e-06 
0.0 -0.9993 0 2.0 1e-06 
0.0 -0.9992 0 2.0 1e-06 
0.0 -0.9991 0 2.0 1e-06 
0.0 -0.999 0 2.0 1e-06 
0.0 -0.9989 0 2.0 1e-06 
0.0 -0.9988 0 2.0 1e-06 
0.0 -0.9987 0 2.0 1e-06 
0.0 -0.9986 0 2.0 1e-06 
0.0 -0.9985 0 2.0 1e-06 
0.0 -0.9984 0 2.0 1e-06 
0.0 -0.9983 0 2.0 1e-06 
0.0 -0.9982 0 2.0 1e-06 
0.0 -0.9981 0 2.0 1e-06 
0.0 -0.998 0 2.0 1e-06 
0.0 -0.9979 0 2.0 1e-06 
0.0 -0.9978 0 2.0 1e-06 
0.0 -0.9977 0 2.0 1e-06 
0.0 -0.9976 0 2.0 1e-06 
0.0 -0.9975 0 2.0 1e-06 
0.0 -0.9974 0 2.0 1e-06 
0.0 -0.9973 0 2.0 1e-06 
0.0 -0.9972 0 2.0 1e-06 
0.0 -0.9971 0 2.0 1e-06 
0.0 -0.997 0 2.0 1e-06 
0.0 -0.9969 0 2.0 1e-06 
0.0 -0.9968 0 2.0 1e-06 
0.0 -0.9967 0 2.0 1e-06 
0.0 -0.9966 0 2.0 1e-06 
0.0 -0.9965 0 2.0 1e-06 
0.0 -0.9964 0 2.0 1e-06 
0.0 -0.9963 0 2.0 1e-06 
0.0 -0.9962 0 2.0 1e-06 
0.0 -0.9961 0 2.0 1e-06 
0.0 -0.996 0 2.0 1e-06 
0.0 -0.9959 0 2.0 1e-06 
0.0 -0.9958 0 2.0 1e-06 
0.0 -0.9957 0 2.0 1e-06 
0.0 -0.9956 0 2.0 1e-06 
0.0 -0.9955 0 2.0 1e-06 
0.0 -0.9954 0 2.0 1e-06 
0.0 -0.9953 0 2.0 1e-06 
0.0 -0.9952 0 2.0 1e-06 
0.0 -0.9951 0 2.0 1e-06 
0.0 -0.995 0 2.0 1e-06 
0.0 -0.9949 0 2.0 1e-06 
0.0 -0.9948 0 2.0 1e-06 
0.0 -0.9947 0 2.0 1e-06 
0.0 -0.9946 0 2.0 1e-06 
0.0 -0.9945 0 2.0 1e-06 
0.0 -0.9944 0 2.0 1e-06 
0.0 -0.9943 0 2.0 1e-06 
0.0 -0.9942 0 2.0 1e-06 
0.0 -0.9941 0 2.0 1e-06 
0.0 -0.994 0 2.0 1e-06 
0.0 -0.9939 0 2.0 1e-06 
0.0 -0.9938 0 2.0 1e-06 
0.0 -0.9937 0 2.0 1e-06 
0.0 -0.9936 0 2.0 1e-06 
0.0 -0.9935 0 2.0 1e-06 
0.0 -0.9934 0 2.0 1e-06 
0.0 -0.9933 0 2.0 1e-06 
0.0 -0.9932 0 2.0 1e-06 
0.0 -0.9931 0 2.0 1e-06 
0.0 -0.993 0 2.0 1e-06 
0.0 -0.9929 0 2.0 1e-06 
0.0 -0.9928 0 2.0 1e-06 
0.0 -0.9927 0 2.0 1e-06 
0.0 -0.9926 0 2.0 1e-06 
0.0 -0.9925 0 2.0 1e-06 
0.0 -0.9924 0 2.0 1e-06 
0.0 -0.9923 0 2.0 1e-06 
0.0 -0.9922 0 2.0 1e-06 
0.0 -0.9921 0 2.0 1e-06 
0.0 -0.992 0 2.0 1e-06 
0.0 -0.9919 0 2.0 1e-06 
0.0 -0.9918 0 2.0 1e-06 
0.0 -0.9917 0 2.0 1e-06 
0.0 -0.9916 0 2.0 1e-06 
0.0 -0.9915 0 2.0 1e-06 
0.0 -0.9914 0 2.0 1e-06 
0.0 -0.9913 0 2.0 1e-06 
0.0 -0.9912 0 2.0 1e-06 
0.0 -0.9911 0 2.0 1e-06 
0.0 -0.991 0 2.0 1e-06 
0.0 -0.9909 0 2.0 1e-06 
0.0 -0.9908 0 2.0 1e-06 
0.0 -0.9907 0 2.0 1e-06 
0.0 -0.9906 0 2.0 1e-06 
0.0 -0.9905 0 2.0 1e-06 
0.0 -0.9904 0 2.0 1e-06 
0.0 -0.9903 0 2.0 1e-06 
0.0 -0.9902 0 2.0 1e-06 
0.0 -0.9901 0 2.0 1e-06 
0.0 -0.99 0 2.0 1e-06 
0.0 -0.9899 0 2.0 1e-06 
0.0 -0.9898 0 2.0 1e-06 
0.0 -0.9897 0 2.0 1e-06 
0.0 -0.9896 0 2.0 1e-06 
0.0 -0.9895 0 2.0 1e-06 
0.0 -0.9894 0 2.0 1e-06 
0.0 -0.9893 0 2.0 1e-06 
0.0 -0.9892 0 2.0 1e-06 
0.0 -0.9891 0 2.0 1e-06 
0.0 -0.989 0 2.0 1e-06 
0.0 -0.9889 0 2.0 1e-06 
0.0 -0.9888 0 2.0 1e-06 
0.0 -0.9887 0 2.0 1e-06 
0.0 -0.9886 0 2.0 1e-06 
0.0 -0.9885 0 2.0 1e-06 
0.0 -0.9884 0 2.0 1e-06 
0.0 -0.9883 0 2.0 1e-06 
0.0 -0.9882 0 2.0 1e-06 
0.0 -0.9881 0 2.0 1e-06 
0.0 -0.988 0 2.0 1e-06 
0.0 -0.9879 0 2.0 1e-06 
0.0 -0.9878 0 2.0 1e-06 
0.0 -0.9877 0 2.0 1e-06 
0.0 -0.9876 0 2.0 1e-06 
0.0 -0.9875 0 2.0 1e-06 
0.0 -0.9874 0 2.0 1e-06 
0.0 -0.9873 0 2.0 1e-06 
0.0 -0.9872 0 2.0 1e-06 
0.0 -0.9871 0 2.0 1e-06 
0.0 -0.987 0 2.0 1e-06 
0.0 -0.9869 0 2.0 1e-06 
0.0 -0.9868 0 2.0 1e-06 
0.0 -0.9867 0 2.0 1e-06 
0.0 -0.9866 0 2.0 1e-06 
0.0 -0.9865 0 2.0 1e-06 
0.0 -0.9864 0 2.0 1e-06 
0.0 -0.9863 0 2.0 1e-06 
0.0 -0.9862 0 2.0 1e-06 
0.0 -0.9861 0 2.0 1e-06 
0.0 -0.986 0 2.0 1e-06 
0.0 -0.9859 0 2.0 1e-06 
0.0 -0.9858 0 2.0 1e-06 
0.0 -0.9857 0 2.0 1e-06 
0.0 -0.9856 0 2.0 1e-06 
0.0 -0.9855 0 2.0 1e-06 
0.0 -0.9854 0 2.0 1e-06 
0.0 -0.9853 0 2.0 1e-06 
0.0 -0.9852 0 2.0 1e-06 
0.0 -0.9851 0 2.0 1e-06 
0.0 -0.985 0 2.0 1e-06 
0.0 -0.9849 0 2.0 1e-06 
0.0 -0.9848 0 2.0 1e-06 
0.0 -0.9847 0 2.0 1e-06 
0.0 -0.9846 0 2.0 1e-06 
0.0 -0.9845 0 2.0 1e-06 
0.0 -0.9844 0 2.0 1e-06 
0.0 -0.9843 0 2.0 1e-06 
0.0 -0.9842 0 2.0 1e-06 
0.0 -0.9841 0 2.0 1e-06 
0.0 -0.984 0 2.0 1e-06 
0.0 -0.9839 0 2.0 1e-06 
0.0 -0.9838 0 2.0 1e-06 
0.0 -0.9837 0 2.0 1e-06 
0.0 -0.9836 0 2.0 1e-06 
0.0 -0.9835 0 2.0 1e-06 
0.0 -0.9834 0 2.0 1e-06 
0.0 -0.9833 0 2.0 1e-06 
0.0 -0.9832 0 2.0 1e-06 
0.0 -0.9831 0 2.0 1e-06 
0.0 -0.983 0 2.0 1e-06 
0.0 -0.9829 0 2.0 1e-06 
0.0 -0.9828 0 2.0 1e-06 
0.0 -0.9827 0 2.0 1e-06 
0.0 -0.9826 0 2.0 1e-06 
0.0 -0.9825 0 2.0 1e-06 
0.0 -0.9824 0 2.0 1e-06 
0.0 -0.9823 0 2.0 1e-06 
0.0 -0.9822 0 2.0 1e-06 
0.0 -0.9821 0 2.0 1e-06 
0.0 -0.982 0 2.0 1e-06 
0.0 -0.9819 0 2.0 1e-06 
0.0 -0.9818 0 2.0 1e-06 
0.0 -0.9817 0 2.0 1e-06 
0.0 -0.9816 0 2.0 1e-06 
0.0 -0.9815 0 2.0 1e-06 
0.0 -0.9814 0 2.0 1e-06 
0.0 -0.9813 0 2.0 1e-06 
0.0 -0.9812 0 2.0 1e-06 
0.0 -0.9811 0 2.0 1e-06 
0.0 -0.981 0 2.0 1e-06 
0.0 -0.9809 0 2.0 1e-06 
0.0 -0.9808 0 2.0 1e-06 
0.0 -0.9807 0 2.0 1e-06 
0.0 -0.9806 0 2.0 1e-06 
0.0 -0.9805 0 2.0 1e-06 
0.0 -0.9804 0 2.0 1e-06 
0.0 -0.9803 0 2.0 1e-06 
0.0 -0.9802 0 2.0 1e-06 
0.0 -0.9801 0 2.0 1e-06 
0.0 -0.98 0 2.0 1e-06 
0.0 -0.9799 0 2.0 1e-06 
0.0 -0.9798 0 2.0 1e-06 
0.0 -0.9797 0 2.0 1e-06 
0.0 -0.9796 0 2.0 1e-06 
0.0 -0.9795 0 2.0 1e-06 
0.0 -0.9794 0 2.0 1e-06 
0.0 -0.9793 0 2.0 1e-06 
0.0 -0.9792 0 2.0 1e-06 
0.0 -0.9791 0 2.0 1e-06 
0.0 -0.979 0 2.0 1e-06 
0.0 -0.9789 0 2.0 1e-06 
0.0 -0.9788 0 2.0 1e-06 
0.0 -0.9787 0 2.0 1e-06 
0.0 -0.9786 0 2.0 1e-06 
0.0 -0.9785 0 2.0 1e-06 
0.0 -0.9784 0 2.0 1e-06 
0.0 -0.9783 0 2.0 1e-06 
0.0 -0.9782 0 2.0 1e-06 
0.0 -0.9781 0 2.0 1e-06 
0.0 -0.978 0 2.0 1e-06 
0.0 -0.9779 0 2.0 1e-06 
0.0 -0.9778 0 2.0 1e-06 
0.0 -0.9777 0 2.0 1e-06 
0.0 -0.9776 0 2.0 1e-06 
0.0 -0.9775 0 2.0 1e-06 
0.0 -0.9774 0 2.0 1e-06 
0.0 -0.9773 0 2.0 1e-06 
0.0 -0.9772 0 2.0 1e-06 
0.0 -0.9771 0 2.0 1e-06 
0.0 -0.977 0 2.0 1e-06 
0.0 -0.9769 0 2.0 1e-06 
0.0 -0.9768 0 2.0 1e-06 
0.0 -0.9767 0 2.0 1e-06 
0.0 -0.9766 0 2.0 1e-06 
0.0 -0.9765 0 2.0 1e-06 
0.0 -0.9764 0 2.0 1e-06 
0.0 -0.9763 0 2.0 1e-06 
0.0 -0.9762 0 2.0 1e-06 
0.0 -0.9761 0 2.0 1e-06 
0.0 -0.976 0 2.0 1e-06 
0.0 -0.9759 0 2.0 1e-06 
0.0 -0.9758 0 2.0 1e-06 
0.0 -0.9757 0 2.0 1e-06 
0.0 -0.9756 0 2.0 1e-06 
0.0 -0.9755 0 2.0 1e-06 
0.0 -0.9754 0 2.0 1e-06 
0.0 -0.9753 0 2.0 1e-06 
0.0 -0.9752 0 2.0 1e-06 
0.0 -0.9751 0 2.0 1e-06 
0.0 -0.975 0 2.0 1e-06 
0.0 -0.9749 0 2.0 1e-06 
0.0 -0.9748 0 2.0 1e-06 
0.0 -0.9747 0 2.0 1e-06 
0.0 -0.9746 0 2.0 1e-06 
0.0 -0.9745 0 2.0 1e-06 
0.0 -0.9744 0 2.0 1e-06 
0.0 -0.9743 0 2.0 1e-06 
0.0 -0.9742 0 2.0 1e-06 
0.0 -0.9741 0 2.0 1e-06 
0.0 -0.974 0 2.0 1e-06 
0.0 -0.9739 0 2.0 1e-06 
0.0 -0.9738 0 2.0 1e-06 
0.0 -0.9737 0 2.0 1e-06 
0.0 -0.9736 0 2.0 1e-06 
0.0 -0.9735 0 2.0 1e-06 
0.0 -0.9734 0 2.0 1e-06 
0.0 -0.9733 0 2.0 1e-06 
0.0 -0.9732 0 2.0 1e-06 
0.0 -0.9731 0 2.0 1e-06 
0.0 -0.973 0 2.0 1e-06 
0.0 -0.9729 0 2.0 1e-06 
0.0 -0.9728 0 2.0 1e-06 
0.0 -0.9727 0 2.0 1e-06 
0.0 -0.9726 0 2.0 1e-06 
0.0 -0.9725 0 2.0 1e-06 
0.0 -0.9724 0 2.0 1e-06 
0.0 -0.9723 0 2.0 1e-06 
0.0 -0.9722 0 2.0 1e-06 
0.0 -0.9721 0 2.0 1e-06 
0.0 -0.972 0 2.0 1e-06 
0.0 -0.9719 0 2.0 1e-06 
0.0 -0.9718 0 2.0 1e-06 
0.0 -0.9717 0 2.0 1e-06 
0.0 -0.9716 0 2.0 1e-06 
0.0 -0.9715 0 2.0 1e-06 
0.0 -0.9714 0 2.0 1e-06 
0.0 -0.9713 0 2.0 1e-06 
0.0 -0.9712 0 2.0 1e-06 
0.0 -0.9711 0 2.0 1e-06 
0.0 -0.971 0 2.0 1e-06 
0.0 -0.9709 0 2.0 1e-06 
0.0 -0.9708 0 2.0 1e-06 
0.0 -0.9707 0 2.0 1e-06 
0.0 -0.9706 0 2.0 1e-06 
0.0 -0.9705 0 2.0 1e-06 
0.0 -0.9704 0 2.0 1e-06 
0.0 -0.9703 0 2.0 1e-06 
0.0 -0.9702 0 2.0 1e-06 
0.0 -0.9701 0 2.0 1e-06 
0.0 -0.97 0 2.0 1e-06 
0.0 -0.9699 0 2.0 1e-06 
0.0 -0.9698 0 2.0 1e-06 
0.0 -0.9697 0 2.0 1e-06 
0.0 -0.9696 0 2.0 1e-06 
0.0 -0.9695 0 2.0 1e-06 
0.0 -0.9694 0 2.0 1e-06 
0.0 -0.9693 0 2.0 1e-06 
0.0 -0.9692 0 2.0 1e-06 
0.0 -0.9691 0 2.0 1e-06 
0.0 -0.969 0 2.0 1e-06 
0.0 -0.9689 0 2.0 1e-06 
0.0 -0.9688 0 2.0 1e-06 
0.0 -0.9687 0 2.0 1e-06 
0.0 -0.9686 0 2.0 1e-06 
0.0 -0.9685 0 2.0 1e-06 
0.0 -0.9684 0 2.0 1e-06 
0.0 -0.9683 0 2.0 1e-06 
0.0 -0.9682 0 2.0 1e-06 
0.0 -0.9681 0 2.0 1e-06 
0.0 -0.968 0 2.0 1e-06 
0.0 -0.9679 0 2.0 1e-06 
0.0 -0.9678 0 2.0 1e-06 
0.0 -0.9677 0 2.0 1e-06 
0.0 -0.9676 0 2.0 1e-06 
0.0 -0.9675 0 2.0 1e-06 
0.0 -0.9674 0 2.0 1e-06 
0.0 -0.9673 0 2.0 1e-06 
0.0 -0.9672 0 2.0 1e-06 
0.0 -0.9671 0 2.0 1e-06 
0.0 -0.967 0 2.0 1e-06 
0.0 -0.9669 0 2.0 1e-06 
0.0 -0.9668 0 2.0 1e-06 
0.0 -0.9667 0 2.0 1e-06 
0.0 -0.9666 0 2.0 1e-06 
0.0 -0.9665 0 2.0 1e-06 
0.0 -0.9664 0 2.0 1e-06 
0.0 -0.9663 0 2.0 1e-06 
0.0 -0.9662 0 2.0 1e-06 
0.0 -0.9661 0 2.0 1e-06 
0.0 -0.966 0 2.0 1e-06 
0.0 -0.9659 0 2.0 1e-06 
0.0 -0.9658 0 2.0 1e-06 
0.0 -0.9657 0 2.0 1e-06 
0.0 -0.9656 0 2.0 1e-06 
0.0 -0.9655 0 2.0 1e-06 
0.0 -0.9654 0 2.0 1e-06 
0.0 -0.9653 0 2.0 1e-06 
0.0 -0.9652 0 2.0 1e-06 
0.0 -0.9651 0 2.0 1e-06 
0.0 -0.965 0 2.0 1e-06 
0.0 -0.9649 0 2.0 1e-06 
0.0 -0.9648 0 2.0 1e-06 
0.0 -0.9647 0 2.0 1e-06 
0.0 -0.9646 0 2.0 1e-06 
0.0 -0.9645 0 2.0 1e-06 
0.0 -0.9644 0 2.0 1e-06 
0.0 -0.9643 0 2.0 1e-06 
0.0 -0.9642 0 2.0 1e-06 
0.0 -0.9641 0 2.0 1e-06 
0.0 -0.964 0 2.0 1e-06 
0.0 -0.9639 0 2.0 1e-06 
0.0 -0.9638 0 2.0 1e-06 
0.0 -0.9637 0 2.0 1e-06 
0.0 -0.9636 0 2.0 1e-06 
0.0 -0.9635 0 2.0 1e-06 
0.0 -0.9634 0 2.0 1e-06 
0.0 -0.9633 0 2.0 1e-06 
0.0 -0.9632 0 2.0 1e-06 
0.0 -0.9631 0 2.0 1e-06 
0.0 -0.963 0 2.0 1e-06 
0.0 -0.9629 0 2.0 1e-06 
0.0 -0.9628 0 2.0 1e-06 
0.0 -0.9627 0 2.0 1e-06 
0.0 -0.9626 0 2.0 1e-06 
0.0 -0.9625 0 2.0 1e-06 
0.0 -0.9624 0 2.0 1e-06 
0.0 -0.9623 0 2.0 1e-06 
0.0 -0.9622 0 2.0 1e-06 
0.0 -0.9621 0 2.0 1e-06 
0.0 -0.962 0 2.0 1e-06 
0.0 -0.9619 0 2.0 1e-06 
0.0 -0.9618 0 2.0 1e-06 
0.0 -0.9617 0 2.0 1e-06 
0.0 -0.9616 0 2.0 1e-06 
0.0 -0.9615 0 2.0 1e-06 
0.0 -0.9614 0 2.0 1e-06 
0.0 -0.9613 0 2.0 1e-06 
0.0 -0.9612 0 2.0 1e-06 
0.0 -0.9611 0 2.0 1e-06 
0.0 -0.961 0 2.0 1e-06 
0.0 -0.9609 0 2.0 1e-06 
0.0 -0.9608 0 2.0 1e-06 
0.0 -0.9607 0 2.0 1e-06 
0.0 -0.9606 0 2.0 1e-06 
0.0 -0.9605 0 2.0 1e-06 
0.0 -0.9604 0 2.0 1e-06 
0.0 -0.9603 0 2.0 1e-06 
0.0 -0.9602 0 2.0 1e-06 
0.0 -0.9601 0 2.0 1e-06 
0.0 -0.96 0 2.0 1e-06 
0.0 -0.9599 0 2.0 1e-06 
0.0 -0.9598 0 2.0 1e-06 
0.0 -0.9597 0 2.0 1e-06 
0.0 -0.9596 0 2.0 1e-06 
0.0 -0.9595 0 2.0 1e-06 
0.0 -0.9594 0 2.0 1e-06 
0.0 -0.9593 0 2.0 1e-06 
0.0 -0.9592 0 2.0 1e-06 
0.0 -0.9591 0 2.0 1e-06 
0.0 -0.959 0 2.0 1e-06 
0.0 -0.9589 0 2.0 1e-06 
0.0 -0.9588 0 2.0 1e-06 
0.0 -0.9587 0 2.0 1e-06 
0.0 -0.9586 0 2.0 1e-06 
0.0 -0.9585 0 2.0 1e-06 
0.0 -0.9584 0 2.0 1e-06 
0.0 -0.9583 0 2.0 1e-06 
0.0 -0.9582 0 2.0 1e-06 
0.0 -0.9581 0 2.0 1e-06 
0.0 -0.958 0 2.0 1e-06 
0.0 -0.9579 0 2.0 1e-06 
0.0 -0.9578 0 2.0 1e-06 
0.0 -0.9577 0 2.0 1e-06 
0.0 -0.9576 0 2.0 1e-06 
0.0 -0.9575 0 2.0 1e-06 
0.0 -0.9574 0 2.0 1e-06 
0.0 -0.9573 0 2.0 1e-06 
0.0 -0.9572 0 2.0 1e-06 
0.0 -0.9571 0 2.0 1e-06 
0.0 -0.957 0 2.0 1e-06 
0.0 -0.9569 0 2.0 1e-06 
0.0 -0.9568 0 2.0 1e-06 
0.0 -0.9567 0 2.0 1e-06 
0.0 -0.9566 0 2.0 1e-06 
0.0 -0.9565 0 2.0 1e-06 
0.0 -0.9564 0 2.0 1e-06 
0.0 -0.9563 0 2.0 1e-06 
0.0 -0.9562 0 2.0 1e-06 
0.0 -0.9561 0 2.0 1e-06 
0.0 -0.956 0 2.0 1e-06 
0.0 -0.9559 0 2.0 1e-06 
0.0 -0.9558 0 2.0 1e-06 
0.0 -0.9557 0 2.0 1e-06 
0.0 -0.9556 0 2.0 1e-06 
0.0 -0.9555 0 2.0 1e-06 
0.0 -0.9554 0 2.0 1e-06 
0.0 -0.9553 0 2.0 1e-06 
0.0 -0.9552 0 2.0 1e-06 
0.0 -0.9551 0 2.0 1e-06 
0.0 -0.955 0 2.0 1e-06 
0.0 -0.9549 0 2.0 1e-06 
0.0 -0.9548 0 2.0 1e-06 
0.0 -0.9547 0 2.0 1e-06 
0.0 -0.9546 0 2.0 1e-06 
0.0 -0.9545 0 2.0 1e-06 
0.0 -0.9544 0 2.0 1e-06 
0.0 -0.9543 0 2.0 1e-06 
0.0 -0.9542 0 2.0 1e-06 
0.0 -0.9541 0 2.0 1e-06 
0.0 -0.954 0 2.0 1e-06 
0.0 -0.9539 0 2.0 1e-06 
0.0 -0.9538 0 2.0 1e-06 
0.0 -0.9537 0 2.0 1e-06 
0.0 -0.9536 0 2.0 1e-06 
0.0 -0.9535 0 2.0 1e-06 
0.0 -0.9534 0 2.0 1e-06 
0.0 -0.9533 0 2.0 1e-06 
0.0 -0.9532 0 2.0 1e-06 
0.0 -0.9531 0 2.0 1e-06 
0.0 -0.953 0 2.0 1e-06 
0.0 -0.9529 0 2.0 1e-06 
0.0 -0.9528 0 2.0 1e-06 
0.0 -0.9527 0 2.0 1e-06 
0.0 -0.9526 0 2.0 1e-06 
0.0 -0.9525 0 2.0 1e-06 
0.0 -0.9524 0 2.0 1e-06 
0.0 -0.9523 0 2.0 1e-06 
0.0 -0.9522 0 2.0 1e-06 
0.0 -0.9521 0 2.0 1e-06 
0.0 -0.952 0 2.0 1e-06 
0.0 -0.9519 0 2.0 1e-06 
0.0 -0.9518 0 2.0 1e-06 
0.0 -0.9517 0 2.0 1e-06 
0.0 -0.9516 0 2.0 1e-06 
0.0 -0.9515 0 2.0 1e-06 
0.0 -0.9514 0 2.0 1e-06 
0.0 -0.9513 0 2.0 1e-06 
0.0 -0.9512 0 2.0 1e-06 
0.0 -0.9511 0 2.0 1e-06 
0.0 -0.951 0 2.0 1e-06 
0.0 -0.9509 0 2.0 1e-06 
0.0 -0.9508 0 2.0 1e-06 
0.0 -0.9507 0 2.0 1e-06 
0.0 -0.9506 0 2.0 1e-06 
0.0 -0.9505 0 2.0 1e-06 
0.0 -0.9504 0 2.0 1e-06 
0.0 -0.9503 0 2.0 1e-06 
0.0 -0.9502 0 2.0 1e-06 
0.0 -0.9501 0 2.0 1e-06 
0.0 -0.95 0 2.0 1e-06 
0.0 -0.9499 0 2.0 1e-06 
0.0 -0.9498 0 2.0 1e-06 
0.0 -0.9497 0 2.0 1e-06 
0.0 -0.9496 0 2.0 1e-06 
0.0 -0.9495 0 2.0 1e-06 
0.0 -0.9494 0 2.0 1e-06 
0.0 -0.9493 0 2.0 1e-06 
0.0 -0.9492 0 2.0 1e-06 
0.0 -0.9491 0 2.0 1e-06 
0.0 -0.949 0 2.0 1e-06 
0.0 -0.9489 0 2.0 1e-06 
0.0 -0.9488 0 2.0 1e-06 
0.0 -0.9487 0 2.0 1e-06 
0.0 -0.9486 0 2.0 1e-06 
0.0 -0.9485 0 2.0 1e-06 
0.0 -0.9484 0 2.0 1e-06 
0.0 -0.9483 0 2.0 1e-06 
0.0 -0.9482 0 2.0 1e-06 
0.0 -0.9481 0 2.0 1e-06 
0.0 -0.948 0 2.0 1e-06 
0.0 -0.9479 0 2.0 1e-06 
0.0 -0.9478 0 2.0 1e-06 
0.0 -0.9477 0 2.0 1e-06 
0.0 -0.9476 0 2.0 1e-06 
0.0 -0.9475 0 2.0 1e-06 
0.0 -0.9474 0 2.0 1e-06 
0.0 -0.9473 0 2.0 1e-06 
0.0 -0.9472 0 2.0 1e-06 
0.0 -0.9471 0 2.0 1e-06 
0.0 -0.947 0 2.0 1e-06 
0.0 -0.9469 0 2.0 1e-06 
0.0 -0.9468 0 2.0 1e-06 
0.0 -0.9467 0 2.0 1e-06 
0.0 -0.9466 0 2.0 1e-06 
0.0 -0.9465 0 2.0 1e-06 
0.0 -0.9464 0 2.0 1e-06 
0.0 -0.9463 0 2.0 1e-06 
0.0 -0.9462 0 2.0 1e-06 
0.0 -0.9461 0 2.0 1e-06 
0.0 -0.946 0 2.0 1e-06 
0.0 -0.9459 0 2.0 1e-06 
0.0 -0.9458 0 2.0 1e-06 
0.0 -0.9457 0 2.0 1e-06 
0.0 -0.9456 0 2.0 1e-06 
0.0 -0.9455 0 2.0 1e-06 
0.0 -0.9454 0 2.0 1e-06 
0.0 -0.9453 0 2.0 1e-06 
0.0 -0.9452 0 2.0 1e-06 
0.0 -0.9451 0 2.0 1e-06 
0.0 -0.945 0 2.0 1e-06 
0.0 -0.9449 0 2.0 1e-06 
0.0 -0.9448 0 2.0 1e-06 
0.0 -0.9447 0 2.0 1e-06 
0.0 -0.9446 0 2.0 1e-06 
0.0 -0.9445 0 2.0 1e-06 
0.0 -0.9444 0 2.0 1e-06 
0.0 -0.9443 0 2.0 1e-06 
0.0 -0.9442 0 2.0 1e-06 
0.0 -0.9441 0 2.0 1e-06 
0.0 -0.944 0 2.0 1e-06 
0.0 -0.9439 0 2.0 1e-06 
0.0 -0.9438 0 2.0 1e-06 
0.0 -0.9437 0 2.0 1e-06 
0.0 -0.9436 0 2.0 1e-06 
0.0 -0.9435 0 2.0 1e-06 
0.0 -0.9434 0 2.0 1e-06 
0.0 -0.9433 0 2.0 1e-06 
0.0 -0.9432 0 2.0 1e-06 
0.0 -0.9431 0 2.0 1e-06 
0.0 -0.943 0 2.0 1e-06 
0.0 -0.9429 0 2.0 1e-06 
0.0 -0.9428 0 2.0 1e-06 
0.0 -0.9427 0 2.0 1e-06 
0.0 -0.9426 0 2.0 1e-06 
0.0 -0.9425 0 2.0 1e-06 
0.0 -0.9424 0 2.0 1e-06 
0.0 -0.9423 0 2.0 1e-06 
0.0 -0.9422 0 2.0 1e-06 
0.0 -0.9421 0 2.0 1e-06 
0.0 -0.942 0 2.0 1e-06 
0.0 -0.9419 0 2.0 1e-06 
0.0 -0.9418 0 2.0 1e-06 
0.0 -0.9417 0 2.0 1e-06 
0.0 -0.9416 0 2.0 1e-06 
0.0 -0.9415 0 2.0 1e-06 
0.0 -0.9414 0 2.0 1e-06 
0.0 -0.9413 0 2.0 1e-06 
0.0 -0.9412 0 2.0 1e-06 
0.0 -0.9411 0 2.0 1e-06 
0.0 -0.941 0 2.0 1e-06 
0.0 -0.9409 0 2.0 1e-06 
0.0 -0.9408 0 2.0 1e-06 
0.0 -0.9407 0 2.0 1e-06 
0.0 -0.9406 0 2.0 1e-06 
0.0 -0.9405 0 2.0 1e-06 
0.0 -0.9404 0 2.0 1e-06 
0.0 -0.9403 0 2.0 1e-06 
0.0 -0.9402 0 2.0 1e-06 
0.0 -0.9401 0 2.0 1e-06 
0.0 -0.94 0 2.0 1e-06 
0.0 -0.9399 0 2.0 1e-06 
0.0 -0.9398 0 2.0 1e-06 
0.0 -0.9397 0 2.0 1e-06 
0.0 -0.9396 0 2.0 1e-06 
0.0 -0.9395 0 2.0 1e-06 
0.0 -0.9394 0 2.0 1e-06 
0.0 -0.9393 0 2.0 1e-06 
0.0 -0.9392 0 2.0 1e-06 
0.0 -0.9391 0 2.0 1e-06 
0.0 -0.939 0 2.0 1e-06 
0.0 -0.9389 0 2.0 1e-06 
0.0 -0.9388 0 2.0 1e-06 
0.0 -0.9387 0 2.0 1e-06 
0.0 -0.9386 0 2.0 1e-06 
0.0 -0.9385 0 2.0 1e-06 
0.0 -0.9384 0 2.0 1e-06 
0.0 -0.9383 0 2.0 1e-06 
0.0 -0.9382 0 2.0 1e-06 
0.0 -0.9381 0 2.0 1e-06 
0.0 -0.938 0 2.0 1e-06 
0.0 -0.9379 0 2.0 1e-06 
0.0 -0.9378 0 2.0 1e-06 
0.0 -0.9377 0 2.0 1e-06 
0.0 -0.9376 0 2.0 1e-06 
0.0 -0.9375 0 2.0 1e-06 
0.0 -0.9374 0 2.0 1e-06 
0.0 -0.9373 0 2.0 1e-06 
0.0 -0.9372 0 2.0 1e-06 
0.0 -0.9371 0 2.0 1e-06 
0.0 -0.937 0 2.0 1e-06 
0.0 -0.9369 0 2.0 1e-06 
0.0 -0.9368 0 2.0 1e-06 
0.0 -0.9367 0 2.0 1e-06 
0.0 -0.9366 0 2.0 1e-06 
0.0 -0.9365 0 2.0 1e-06 
0.0 -0.9364 0 2.0 1e-06 
0.0 -0.9363 0 2.0 1e-06 
0.0 -0.9362 0 2.0 1e-06 
0.0 -0.9361 0 2.0 1e-06 
0.0 -0.936 0 2.0 1e-06 
0.0 -0.9359 0 2.0 1e-06 
0.0 -0.9358 0 2.0 1e-06 
0.0 -0.9357 0 2.0 1e-06 
0.0 -0.9356 0 2.0 1e-06 
0.0 -0.9355 0 2.0 1e-06 
0.0 -0.9354 0 2.0 1e-06 
0.0 -0.9353 0 2.0 1e-06 
0.0 -0.9352 0 2.0 1e-06 
0.0 -0.9351 0 2.0 1e-06 
0.0 -0.935 0 2.0 1e-06 
0.0 -0.9349 0 2.0 1e-06 
0.0 -0.9348 0 2.0 1e-06 
0.0 -0.9347 0 2.0 1e-06 
0.0 -0.9346 0 2.0 1e-06 
0.0 -0.9345 0 2.0 1e-06 
0.0 -0.9344 0 2.0 1e-06 
0.0 -0.9343 0 2.0 1e-06 
0.0 -0.9342 0 2.0 1e-06 
0.0 -0.9341 0 2.0 1e-06 
0.0 -0.934 0 2.0 1e-06 
0.0 -0.9339 0 2.0 1e-06 
0.0 -0.9338 0 2.0 1e-06 
0.0 -0.9337 0 2.0 1e-06 
0.0 -0.9336 0 2.0 1e-06 
0.0 -0.9335 0 2.0 1e-06 
0.0 -0.9334 0 2.0 1e-06 
0.0 -0.9333 0 2.0 1e-06 
0.0 -0.9332 0 2.0 1e-06 
0.0 -0.9331 0 2.0 1e-06 
0.0 -0.933 0 2.0 1e-06 
0.0 -0.9329 0 2.0 1e-06 
0.0 -0.9328 0 2.0 1e-06 
0.0 -0.9327 0 2.0 1e-06 
0.0 -0.9326 0 2.0 1e-06 
0.0 -0.9325 0 2.0 1e-06 
0.0 -0.9324 0 2.0 1e-06 
0.0 -0.9323 0 2.0 1e-06 
0.0 -0.9322 0 2.0 1e-06 
0.0 -0.9321 0 2.0 1e-06 
0.0 -0.932 0 2.0 1e-06 
0.0 -0.9319 0 2.0 1e-06 
0.0 -0.9318 0 2.0 1e-06 
0.0 -0.9317 0 2.0 1e-06 
0.0 -0.9316 0 2.0 1e-06 
0.0 -0.9315 0 2.0 1e-06 
0.0 -0.9314 0 2.0 1e-06 
0.0 -0.9313 0 2.0 1e-06 
0.0 -0.9312 0 2.0 1e-06 
0.0 -0.9311 0 2.0 1e-06 
0.0 -0.931 0 2.0 1e-06 
0.0 -0.9309 0 2.0 1e-06 
0.0 -0.9308 0 2.0 1e-06 
0.0 -0.9307 0 2.0 1e-06 
0.0 -0.9306 0 2.0 1e-06 
0.0 -0.9305 0 2.0 1e-06 
0.0 -0.9304 0 2.0 1e-06 
0.0 -0.9303 0 2.0 1e-06 
0.0 -0.9302 0 2.0 1e-06 
0.0 -0.9301 0 2.0 1e-06 
0.0 -0.93 0 2.0 1e-06 
0.0 -0.9299 0 2.0 1e-06 
0.0 -0.9298 0 2.0 1e-06 
0.0 -0.9297 0 2.0 1e-06 
0.0 -0.9296 0 2.0 1e-06 
0.0 -0.9295 0 2.0 1e-06 
0.0 -0.9294 0 2.0 1e-06 
0.0 -0.9293 0 2.0 1e-06 
0.0 -0.9292 0 2.0 1e-06 
0.0 -0.9291 0 2.0 1e-06 
0.0 -0.929 0 2.0 1e-06 
0.0 -0.9289 0 2.0 1e-06 
0.0 -0.9288 0 2.0 1e-06 
0.0 -0.9287 0 2.0 1e-06 
0.0 -0.9286 0 2.0 1e-06 
0.0 -0.9285 0 2.0 1e-06 
0.0 -0.9284 0 2.0 1e-06 
0.0 -0.9283 0 2.0 1e-06 
0.0 -0.9282 0 2.0 1e-06 
0.0 -0.9281 0 2.0 1e-06 
0.0 -0.928 0 2.0 1e-06 
0.0 -0.9279 0 2.0 1e-06 
0.0 -0.9278 0 2.0 1e-06 
0.0 -0.9277 0 2.0 1e-06 
0.0 -0.9276 0 2.0 1e-06 
0.0 -0.9275 0 2.0 1e-06 
0.0 -0.9274 0 2.0 1e-06 
0.0 -0.9273 0 2.0 1e-06 
0.0 -0.9272 0 2.0 1e-06 
0.0 -0.9271 0 2.0 1e-06 
0.0 -0.927 0 2.0 1e-06 
0.0 -0.9269 0 2.0 1e-06 
0.0 -0.9268 0 2.0 1e-06 
0.0 -0.9267 0 2.0 1e-06 
0.0 -0.9266 0 2.0 1e-06 
0.0 -0.9265 0 2.0 1e-06 
0.0 -0.9264 0 2.0 1e-06 
0.0 -0.9263 0 2.0 1e-06 
0.0 -0.9262 0 2.0 1e-06 
0.0 -0.9261 0 2.0 1e-06 
0.0 -0.926 0 2.0 1e-06 
0.0 -0.9259 0 2.0 1e-06 
0.0 -0.9258 0 2.0 1e-06 
0.0 -0.9257 0 2.0 1e-06 
0.0 -0.9256 0 2.0 1e-06 
0.0 -0.9255 0 2.0 1e-06 
0.0 -0.9254 0 2.0 1e-06 
0.0 -0.9253 0 2.0 1e-06 
0.0 -0.9252 0 2.0 1e-06 
0.0 -0.9251 0 2.0 1e-06 
0.0 -0.925 0 2.0 1e-06 
0.0 -0.9249 0 2.0 1e-06 
0.0 -0.9248 0 2.0 1e-06 
0.0 -0.9247 0 2.0 1e-06 
0.0 -0.9246 0 2.0 1e-06 
0.0 -0.9245 0 2.0 1e-06 
0.0 -0.9244 0 2.0 1e-06 
0.0 -0.9243 0 2.0 1e-06 
0.0 -0.9242 0 2.0 1e-06 
0.0 -0.9241 0 2.0 1e-06 
0.0 -0.924 0 2.0 1e-06 
0.0 -0.9239 0 2.0 1e-06 
0.0 -0.9238 0 2.0 1e-06 
0.0 -0.9237 0 2.0 1e-06 
0.0 -0.9236 0 2.0 1e-06 
0.0 -0.9235 0 2.0 1e-06 
0.0 -0.9234 0 2.0 1e-06 
0.0 -0.9233 0 2.0 1e-06 
0.0 -0.9232 0 2.0 1e-06 
0.0 -0.9231 0 2.0 1e-06 
0.0 -0.923 0 2.0 1e-06 
0.0 -0.9229 0 2.0 1e-06 
0.0 -0.9228 0 2.0 1e-06 
0.0 -0.9227 0 2.0 1e-06 
0.0 -0.9226 0 2.0 1e-06 
0.0 -0.9225 0 2.0 1e-06 
0.0 -0.9224 0 2.0 1e-06 
0.0 -0.9223 0 2.0 1e-06 
0.0 -0.9222 0 2.0 1e-06 
0.0 -0.9221 0 2.0 1e-06 
0.0 -0.922 0 2.0 1e-06 
0.0 -0.9219 0 2.0 1e-06 
0.0 -0.9218 0 2.0 1e-06 
0.0 -0.9217 0 2.0 1e-06 
0.0 -0.9216 0 2.0 1e-06 
0.0 -0.9215 0 2.0 1e-06 
0.0 -0.9214 0 2.0 1e-06 
0.0 -0.9213 0 2.0 1e-06 
0.0 -0.9212 0 2.0 1e-06 
0.0 -0.9211 0 2.0 1e-06 
0.0 -0.921 0 2.0 1e-06 
0.0 -0.9209 0 2.0 1e-06 
0.0 -0.9208 0 2.0 1e-06 
0.0 -0.9207 0 2.0 1e-06 
0.0 -0.9206 0 2.0 1e-06 
0.0 -0.9205 0 2.0 1e-06 
0.0 -0.9204 0 2.0 1e-06 
0.0 -0.9203 0 2.0 1e-06 
0.0 -0.9202 0 2.0 1e-06 
0.0 -0.9201 0 2.0 1e-06 
0.0 -0.92 0 2.0 1e-06 
0.0 -0.9199 0 2.0 1e-06 
0.0 -0.9198 0 2.0 1e-06 
0.0 -0.9197 0 2.0 1e-06 
0.0 -0.9196 0 2.0 1e-06 
0.0 -0.9195 0 2.0 1e-06 
0.0 -0.9194 0 2.0 1e-06 
0.0 -0.9193 0 2.0 1e-06 
0.0 -0.9192 0 2.0 1e-06 
0.0 -0.9191 0 2.0 1e-06 
0.0 -0.919 0 2.0 1e-06 
0.0 -0.9189 0 2.0 1e-06 
0.0 -0.9188 0 2.0 1e-06 
0.0 -0.9187 0 2.0 1e-06 
0.0 -0.9186 0 2.0 1e-06 
0.0 -0.9185 0 2.0 1e-06 
0.0 -0.9184 0 2.0 1e-06 
0.0 -0.9183 0 2.0 1e-06 
0.0 -0.9182 0 2.0 1e-06 
0.0 -0.9181 0 2.0 1e-06 
0.0 -0.918 0 2.0 1e-06 
0.0 -0.9179 0 2.0 1e-06 
0.0 -0.9178 0 2.0 1e-06 
0.0 -0.9177 0 2.0 1e-06 
0.0 -0.9176 0 2.0 1e-06 
0.0 -0.9175 0 2.0 1e-06 
0.0 -0.9174 0 2.0 1e-06 
0.0 -0.9173 0 2.0 1e-06 
0.0 -0.9172 0 2.0 1e-06 
0.0 -0.9171 0 2.0 1e-06 
0.0 -0.917 0 2.0 1e-06 
0.0 -0.9169 0 2.0 1e-06 
0.0 -0.9168 0 2.0 1e-06 
0.0 -0.9167 0 2.0 1e-06 
0.0 -0.9166 0 2.0 1e-06 
0.0 -0.9165 0 2.0 1e-06 
0.0 -0.9164 0 2.0 1e-06 
0.0 -0.9163 0 2.0 1e-06 
0.0 -0.9162 0 2.0 1e-06 
0.0 -0.9161 0 2.0 1e-06 
0.0 -0.916 0 2.0 1e-06 
0.0 -0.9159 0 2.0 1e-06 
0.0 -0.9158 0 2.0 1e-06 
0.0 -0.9157 0 2.0 1e-06 
0.0 -0.9156 0 2.0 1e-06 
0.0 -0.9155 0 2.0 1e-06 
0.0 -0.9154 0 2.0 1e-06 
0.0 -0.9153 0 2.0 1e-06 
0.0 -0.9152 0 2.0 1e-06 
0.0 -0.9151 0 2.0 1e-06 
0.0 -0.915 0 2.0 1e-06 
0.0 -0.9149 0 2.0 1e-06 
0.0 -0.9148 0 2.0 1e-06 
0.0 -0.9147 0 2.0 1e-06 
0.0 -0.9146 0 2.0 1e-06 
0.0 -0.9145 0 2.0 1e-06 
0.0 -0.9144 0 2.0 1e-06 
0.0 -0.9143 0 2.0 1e-06 
0.0 -0.9142 0 2.0 1e-06 
0.0 -0.9141 0 2.0 1e-06 
0.0 -0.914 0 2.0 1e-06 
0.0 -0.9139 0 2.0 1e-06 
0.0 -0.9138 0 2.0 1e-06 
0.0 -0.9137 0 2.0 1e-06 
0.0 -0.9136 0 2.0 1e-06 
0.0 -0.9135 0 2.0 1e-06 
0.0 -0.9134 0 2.0 1e-06 
0.0 -0.9133 0 2.0 1e-06 
0.0 -0.9132 0 2.0 1e-06 
0.0 -0.9131 0 2.0 1e-06 
0.0 -0.913 0 2.0 1e-06 
0.0 -0.9129 0 2.0 1e-06 
0.0 -0.9128 0 2.0 1e-06 
0.0 -0.9127 0 2.0 1e-06 
0.0 -0.9126 0 2.0 1e-06 
0.0 -0.9125 0 2.0 1e-06 
0.0 -0.9124 0 2.0 1e-06 
0.0 -0.9123 0 2.0 1e-06 
0.0 -0.9122 0 2.0 1e-06 
0.0 -0.9121 0 2.0 1e-06 
0.0 -0.912 0 2.0 1e-06 
0.0 -0.9119 0 2.0 1e-06 
0.0 -0.9118 0 2.0 1e-06 
0.0 -0.9117 0 2.0 1e-06 
0.0 -0.9116 0 2.0 1e-06 
0.0 -0.9115 0 2.0 1e-06 
0.0 -0.9114 0 2.0 1e-06 
0.0 -0.9113 0 2.0 1e-06 
0.0 -0.9112 0 2.0 1e-06 
0.0 -0.9111 0 2.0 1e-06 
0.0 -0.911 0 2.0 1e-06 
0.0 -0.9109 0 2.0 1e-06 
0.0 -0.9108 0 2.0 1e-06 
0.0 -0.9107 0 2.0 1e-06 
0.0 -0.9106 0 2.0 1e-06 
0.0 -0.9105 0 2.0 1e-06 
0.0 -0.9104 0 2.0 1e-06 
0.0 -0.9103 0 2.0 1e-06 
0.0 -0.9102 0 2.0 1e-06 
0.0 -0.9101 0 2.0 1e-06 
0.0 -0.91 0 2.0 1e-06 
0.0 -0.9099 0 2.0 1e-06 
0.0 -0.9098 0 2.0 1e-06 
0.0 -0.9097 0 2.0 1e-06 
0.0 -0.9096 0 2.0 1e-06 
0.0 -0.9095 0 2.0 1e-06 
0.0 -0.9094 0 2.0 1e-06 
0.0 -0.9093 0 2.0 1e-06 
0.0 -0.9092 0 2.0 1e-06 
0.0 -0.9091 0 2.0 1e-06 
0.0 -0.909 0 2.0 1e-06 
0.0 -0.9089 0 2.0 1e-06 
0.0 -0.9088 0 2.0 1e-06 
0.0 -0.9087 0 2.0 1e-06 
0.0 -0.9086 0 2.0 1e-06 
0.0 -0.9085 0 2.0 1e-06 
0.0 -0.9084 0 2.0 1e-06 
0.0 -0.9083 0 2.0 1e-06 
0.0 -0.9082 0 2.0 1e-06 
0.0 -0.9081 0 2.0 1e-06 
0.0 -0.908 0 2.0 1e-06 
0.0 -0.9079 0 2.0 1e-06 
0.0 -0.9078 0 2.0 1e-06 
0.0 -0.9077 0 2.0 1e-06 
0.0 -0.9076 0 2.0 1e-06 
0.0 -0.9075 0 2.0 1e-06 
0.0 -0.9074 0 2.0 1e-06 
0.0 -0.9073 0 2.0 1e-06 
0.0 -0.9072 0 2.0 1e-06 
0.0 -0.9071 0 2.0 1e-06 
0.0 -0.907 0 2.0 1e-06 
0.0 -0.9069 0 2.0 1e-06 
0.0 -0.9068 0 2.0 1e-06 
0.0 -0.9067 0 2.0 1e-06 
0.0 -0.9066 0 2.0 1e-06 
0.0 -0.9065 0 2.0 1e-06 
0.0 -0.9064 0 2.0 1e-06 
0.0 -0.9063 0 2.0 1e-06 
0.0 -0.9062 0 2.0 1e-06 
0.0 -0.9061 0 2.0 1e-06 
0.0 -0.906 0 2.0 1e-06 
0.0 -0.9059 0 2.0 1e-06 
0.0 -0.9058 0 2.0 1e-06 
0.0 -0.9057 0 2.0 1e-06 
0.0 -0.9056 0 2.0 1e-06 
0.0 -0.9055 0 2.0 1e-06 
0.0 -0.9054 0 2.0 1e-06 
0.0 -0.9053 0 2.0 1e-06 
0.0 -0.9052 0 2.0 1e-06 
0.0 -0.9051 0 2.0 1e-06 
0.0 -0.905 0 2.0 1e-06 
0.0 -0.9049 0 2.0 1e-06 
0.0 -0.9048 0 2.0 1e-06 
0.0 -0.9047 0 2.0 1e-06 
0.0 -0.9046 0 2.0 1e-06 
0.0 -0.9045 0 2.0 1e-06 
0.0 -0.9044 0 2.0 1e-06 
0.0 -0.9043 0 2.0 1e-06 
0.0 -0.9042 0 2.0 1e-06 
0.0 -0.9041 0 2.0 1e-06 
0.0 -0.904 0 2.0 1e-06 
0.0 -0.9039 0 2.0 1e-06 
0.0 -0.9038 0 2.0 1e-06 
0.0 -0.9037 0 2.0 1e-06 
0.0 -0.9036 0 2.0 1e-06 
0.0 -0.9035 0 2.0 1e-06 
0.0 -0.9034 0 2.0 1e-06 
0.0 -0.9033 0 2.0 1e-06 
0.0 -0.9032 0 2.0 1e-06 
0.0 -0.9031 0 2.0 1e-06 
0.0 -0.903 0 2.0 1e-06 
0.0 -0.9029 0 2.0 1e-06 
0.0 -0.9028 0 2.0 1e-06 
0.0 -0.9027 0 2.0 1e-06 
0.0 -0.9026 0 2.0 1e-06 
0.0 -0.9025 0 2.0 1e-06 
0.0 -0.9024 0 2.0 1e-06 
0.0 -0.9023 0 2.0 1e-06 
0.0 -0.9022 0 2.0 1e-06 
0.0 -0.9021 0 2.0 1e-06 
0.0 -0.902 0 2.0 1e-06 
0.0 -0.9019 0 2.0 1e-06 
0.0 -0.9018 0 2.0 1e-06 
0.0 -0.9017 0 2.0 1e-06 
0.0 -0.9016 0 2.0 1e-06 
0.0 -0.9015 0 2.0 1e-06 
0.0 -0.9014 0 2.0 1e-06 
0.0 -0.9013 0 2.0 1e-06 
0.0 -0.9012 0 2.0 1e-06 
0.0 -0.9011 0 2.0 1e-06 
0.0 -0.901 0 2.0 1e-06 
0.0 -0.9009 0 2.0 1e-06 
0.0 -0.9008 0 2.0 1e-06 
0.0 -0.9007 0 2.0 1e-06 
0.0 -0.9006 0 2.0 1e-06 
0.0 -0.9005 0 2.0 1e-06 
0.0 -0.9004 0 2.0 1e-06 
0.0 -0.9003 0 2.0 1e-06 
0.0 -0.9002 0 2.0 1e-06 
0.0 -0.9001 0 2.0 1e-06 
0.0 -0.9 0 2.0 1e-06 
0.0 -0.8999 0 2.0 1e-06 
0.0 -0.8998 0 2.0 1e-06 
0.0 -0.8997 0 2.0 1e-06 
0.0 -0.8996 0 2.0 1e-06 
0.0 -0.8995 0 2.0 1e-06 
0.0 -0.8994 0 2.0 1e-06 
0.0 -0.8993 0 2.0 1e-06 
0.0 -0.8992 0 2.0 1e-06 
0.0 -0.8991 0 2.0 1e-06 
0.0 -0.899 0 2.0 1e-06 
0.0 -0.8989 0 2.0 1e-06 
0.0 -0.8988 0 2.0 1e-06 
0.0 -0.8987 0 2.0 1e-06 
0.0 -0.8986 0 2.0 1e-06 
0.0 -0.8985 0 2.0 1e-06 
0.0 -0.8984 0 2.0 1e-06 
0.0 -0.8983 0 2.0 1e-06 
0.0 -0.8982 0 2.0 1e-06 
0.0 -0.8981 0 2.0 1e-06 
0.0 -0.898 0 2.0 1e-06 
0.0 -0.8979 0 2.0 1e-06 
0.0 -0.8978 0 2.0 1e-06 
0.0 -0.8977 0 2.0 1e-06 
0.0 -0.8976 0 2.0 1e-06 
0.0 -0.8975 0 2.0 1e-06 
0.0 -0.8974 0 2.0 1e-06 
0.0 -0.8973 0 2.0 1e-06 
0.0 -0.8972 0 2.0 1e-06 
0.0 -0.8971 0 2.0 1e-06 
0.0 -0.897 0 2.0 1e-06 
0.0 -0.8969 0 2.0 1e-06 
0.0 -0.8968 0 2.0 1e-06 
0.0 -0.8967 0 2.0 1e-06 
0.0 -0.8966 0 2.0 1e-06 
0.0 -0.8965 0 2.0 1e-06 
0.0 -0.8964 0 2.0 1e-06 
0.0 -0.8963 0 2.0 1e-06 
0.0 -0.8962 0 2.0 1e-06 
0.0 -0.8961 0 2.0 1e-06 
0.0 -0.896 0 2.0 1e-06 
0.0 -0.8959 0 2.0 1e-06 
0.0 -0.8958 0 2.0 1e-06 
0.0 -0.8957 0 2.0 1e-06 
0.0 -0.8956 0 2.0 1e-06 
0.0 -0.8955 0 2.0 1e-06 
0.0 -0.8954 0 2.0 1e-06 
0.0 -0.8953 0 2.0 1e-06 
0.0 -0.8952 0 2.0 1e-06 
0.0 -0.8951 0 2.0 1e-06 
0.0 -0.895 0 2.0 1e-06 
0.0 -0.8949 0 2.0 1e-06 
0.0 -0.8948 0 2.0 1e-06 
0.0 -0.8947 0 2.0 1e-06 
0.0 -0.8946 0 2.0 1e-06 
0.0 -0.8945 0 2.0 1e-06 
0.0 -0.8944 0 2.0 1e-06 
0.0 -0.8943 0 2.0 1e-06 
0.0 -0.8942 0 2.0 1e-06 
0.0 -0.8941 0 2.0 1e-06 
0.0 -0.894 0 2.0 1e-06 
0.0 -0.8939 0 2.0 1e-06 
0.0 -0.8938 0 2.0 1e-06 
0.0 -0.8937 0 2.0 1e-06 
0.0 -0.8936 0 2.0 1e-06 
0.0 -0.8935 0 2.0 1e-06 
0.0 -0.8934 0 2.0 1e-06 
0.0 -0.8933 0 2.0 1e-06 
0.0 -0.8932 0 2.0 1e-06 
0.0 -0.8931 0 2.0 1e-06 
0.0 -0.893 0 2.0 1e-06 
0.0 -0.8929 0 2.0 1e-06 
0.0 -0.8928 0 2.0 1e-06 
0.0 -0.8927 0 2.0 1e-06 
0.0 -0.8926 0 2.0 1e-06 
0.0 -0.8925 0 2.0 1e-06 
0.0 -0.8924 0 2.0 1e-06 
0.0 -0.8923 0 2.0 1e-06 
0.0 -0.8922 0 2.0 1e-06 
0.0 -0.8921 0 2.0 1e-06 
0.0 -0.892 0 2.0 1e-06 
0.0 -0.8919 0 2.0 1e-06 
0.0 -0.8918 0 2.0 1e-06 
0.0 -0.8917 0 2.0 1e-06 
0.0 -0.8916 0 2.0 1e-06 
0.0 -0.8915 0 2.0 1e-06 
0.0 -0.8914 0 2.0 1e-06 
0.0 -0.8913 0 2.0 1e-06 
0.0 -0.8912 0 2.0 1e-06 
0.0 -0.8911 0 2.0 1e-06 
0.0 -0.891 0 2.0 1e-06 
0.0 -0.8909 0 2.0 1e-06 
0.0 -0.8908 0 2.0 1e-06 
0.0 -0.8907 0 2.0 1e-06 
0.0 -0.8906 0 2.0 1e-06 
0.0 -0.8905 0 2.0 1e-06 
0.0 -0.8904 0 2.0 1e-06 
0.0 -0.8903 0 2.0 1e-06 
0.0 -0.8902 0 2.0 1e-06 
0.0 -0.8901 0 2.0 1e-06 
0.0 -0.89 0 2.0 1e-06 
0.0 -0.8899 0 2.0 1e-06 
0.0 -0.8898 0 2.0 1e-06 
0.0 -0.8897 0 2.0 1e-06 
0.0 -0.8896 0 2.0 1e-06 
0.0 -0.8895 0 2.0 1e-06 
0.0 -0.8894 0 2.0 1e-06 
0.0 -0.8893 0 2.0 1e-06 
0.0 -0.8892 0 2.0 1e-06 
0.0 -0.8891 0 2.0 1e-06 
0.0 -0.889 0 2.0 1e-06 
0.0 -0.8889 0 2.0 1e-06 
0.0 -0.8888 0 2.0 1e-06 
0.0 -0.8887 0 2.0 1e-06 
0.0 -0.8886 0 2.0 1e-06 
0.0 -0.8885 0 2.0 1e-06 
0.0 -0.8884 0 2.0 1e-06 
0.0 -0.8883 0 2.0 1e-06 
0.0 -0.8882 0 2.0 1e-06 
0.0 -0.8881 0 2.0 1e-06 
0.0 -0.888 0 2.0 1e-06 
0.0 -0.8879 0 2.0 1e-06 
0.0 -0.8878 0 2.0 1e-06 
0.0 -0.8877 0 2.0 1e-06 
0.0 -0.8876 0 2.0 1e-06 
0.0 -0.8875 0 2.0 1e-06 
0.0 -0.8874 0 2.0 1e-06 
0.0 -0.8873 0 2.0 1e-06 
0.0 -0.8872 0 2.0 1e-06 
0.0 -0.8871 0 2.0 1e-06 
0.0 -0.887 0 2.0 1e-06 
0.0 -0.8869 0 2.0 1e-06 
0.0 -0.8868 0 2.0 1e-06 
0.0 -0.8867 0 2.0 1e-06 
0.0 -0.8866 0 2.0 1e-06 
0.0 -0.8865 0 2.0 1e-06 
0.0 -0.8864 0 2.0 1e-06 
0.0 -0.8863 0 2.0 1e-06 
0.0 -0.8862 0 2.0 1e-06 
0.0 -0.8861 0 2.0 1e-06 
0.0 -0.886 0 2.0 1e-06 
0.0 -0.8859 0 2.0 1e-06 
0.0 -0.8858 0 2.0 1e-06 
0.0 -0.8857 0 2.0 1e-06 
0.0 -0.8856 0 2.0 1e-06 
0.0 -0.8855 0 2.0 1e-06 
0.0 -0.8854 0 2.0 1e-06 
0.0 -0.8853 0 2.0 1e-06 
0.0 -0.8852 0 2.0 1e-06 
0.0 -0.8851 0 2.0 1e-06 
0.0 -0.885 0 2.0 1e-06 
0.0 -0.8849 0 2.0 1e-06 
0.0 -0.8848 0 2.0 1e-06 
0.0 -0.8847 0 2.0 1e-06 
0.0 -0.8846 0 2.0 1e-06 
0.0 -0.8845 0 2.0 1e-06 
0.0 -0.8844 0 2.0 1e-06 
0.0 -0.8843 0 2.0 1e-06 
0.0 -0.8842 0 2.0 1e-06 
0.0 -0.8841 0 2.0 1e-06 
0.0 -0.884 0 2.0 1e-06 
0.0 -0.8839 0 2.0 1e-06 
0.0 -0.8838 0 2.0 1e-06 
0.0 -0.8837 0 2.0 1e-06 
0.0 -0.8836 0 2.0 1e-06 
0.0 -0.8835 0 2.0 1e-06 
0.0 -0.8834 0 2.0 1e-06 
0.0 -0.8833 0 2.0 1e-06 
0.0 -0.8832 0 2.0 1e-06 
0.0 -0.8831 0 2.0 1e-06 
0.0 -0.883 0 2.0 1e-06 
0.0 -0.8829 0 2.0 1e-06 
0.0 -0.8828 0 2.0 1e-06 
0.0 -0.8827 0 2.0 1e-06 
0.0 -0.8826 0 2.0 1e-06 
0.0 -0.8825 0 2.0 1e-06 
0.0 -0.8824 0 2.0 1e-06 
0.0 -0.8823 0 2.0 1e-06 
0.0 -0.8822 0 2.0 1e-06 
0.0 -0.8821 0 2.0 1e-06 
0.0 -0.882 0 2.0 1e-06 
0.0 -0.8819 0 2.0 1e-06 
0.0 -0.8818 0 2.0 1e-06 
0.0 -0.8817 0 2.0 1e-06 
0.0 -0.8816 0 2.0 1e-06 
0.0 -0.8815 0 2.0 1e-06 
0.0 -0.8814 0 2.0 1e-06 
0.0 -0.8813 0 2.0 1e-06 
0.0 -0.8812 0 2.0 1e-06 
0.0 -0.8811 0 2.0 1e-06 
0.0 -0.881 0 2.0 1e-06 
0.0 -0.8809 0 2.0 1e-06 
0.0 -0.8808 0 2.0 1e-06 
0.0 -0.8807 0 2.0 1e-06 
0.0 -0.8806 0 2.0 1e-06 
0.0 -0.8805 0 2.0 1e-06 
0.0 -0.8804 0 2.0 1e-06 
0.0 -0.8803 0 2.0 1e-06 
0.0 -0.8802 0 2.0 1e-06 
0.0 -0.8801 0 2.0 1e-06 
0.0 -0.88 0 2.0 1e-06 
0.0 -0.8799 0 2.0 1e-06 
0.0 -0.8798 0 2.0 1e-06 
0.0 -0.8797 0 2.0 1e-06 
0.0 -0.8796 0 2.0 1e-06 
0.0 -0.8795 0 2.0 1e-06 
0.0 -0.8794 0 2.0 1e-06 
0.0 -0.8793 0 2.0 1e-06 
0.0 -0.8792 0 2.0 1e-06 
0.0 -0.8791 0 2.0 1e-06 
0.0 -0.879 0 2.0 1e-06 
0.0 -0.8789 0 2.0 1e-06 
0.0 -0.8788 0 2.0 1e-06 
0.0 -0.8787 0 2.0 1e-06 
0.0 -0.8786 0 2.0 1e-06 
0.0 -0.8785 0 2.0 1e-06 
0.0 -0.8784 0 2.0 1e-06 
0.0 -0.8783 0 2.0 1e-06 
0.0 -0.8782 0 2.0 1e-06 
0.0 -0.8781 0 2.0 1e-06 
0.0 -0.878 0 2.0 1e-06 
0.0 -0.8779 0 2.0 1e-06 
0.0 -0.8778 0 2.0 1e-06 
0.0 -0.8777 0 2.0 1e-06 
0.0 -0.8776 0 2.0 1e-06 
0.0 -0.8775 0 2.0 1e-06 
0.0 -0.8774 0 2.0 1e-06 
0.0 -0.8773 0 2.0 1e-06 
0.0 -0.8772 0 2.0 1e-06 
0.0 -0.8771 0 2.0 1e-06 
0.0 -0.877 0 2.0 1e-06 
0.0 -0.8769 0 2.0 1e-06 
0.0 -0.8768 0 2.0 1e-06 
0.0 -0.8767 0 2.0 1e-06 
0.0 -0.8766 0 2.0 1e-06 
0.0 -0.8765 0 2.0 1e-06 
0.0 -0.8764 0 2.0 1e-06 
0.0 -0.8763 0 2.0 1e-06 
0.0 -0.8762 0 2.0 1e-06 
0.0 -0.8761 0 2.0 1e-06 
0.0 -0.876 0 2.0 1e-06 
0.0 -0.8759 0 2.0 1e-06 
0.0 -0.8758 0 2.0 1e-06 
0.0 -0.8757 0 2.0 1e-06 
0.0 -0.8756 0 2.0 1e-06 
0.0 -0.8755 0 2.0 1e-06 
0.0 -0.8754 0 2.0 1e-06 
0.0 -0.8753 0 2.0 1e-06 
0.0 -0.8752 0 2.0 1e-06 
0.0 -0.8751 0 2.0 1e-06 
0.0 -0.875 0 2.0 1e-06 
0.0 -0.8749 0 2.0 1e-06 
0.0 -0.8748 0 2.0 1e-06 
0.0 -0.8747 0 2.0 1e-06 
0.0 -0.8746 0 2.0 1e-06 
0.0 -0.8745 0 2.0 1e-06 
0.0 -0.8744 0 2.0 1e-06 
0.0 -0.8743 0 2.0 1e-06 
0.0 -0.8742 0 2.0 1e-06 
0.0 -0.8741 0 2.0 1e-06 
0.0 -0.874 0 2.0 1e-06 
0.0 -0.8739 0 2.0 1e-06 
0.0 -0.8738 0 2.0 1e-06 
0.0 -0.8737 0 2.0 1e-06 
0.0 -0.8736 0 2.0 1e-06 
0.0 -0.8735 0 2.0 1e-06 
0.0 -0.8734 0 2.0 1e-06 
0.0 -0.8733 0 2.0 1e-06 
0.0 -0.8732 0 2.0 1e-06 
0.0 -0.8731 0 2.0 1e-06 
0.0 -0.873 0 2.0 1e-06 
0.0 -0.8729 0 2.0 1e-06 
0.0 -0.8728 0 2.0 1e-06 
0.0 -0.8727 0 2.0 1e-06 
0.0 -0.8726 0 2.0 1e-06 
0.0 -0.8725 0 2.0 1e-06 
0.0 -0.8724 0 2.0 1e-06 
0.0 -0.8723 0 2.0 1e-06 
0.0 -0.8722 0 2.0 1e-06 
0.0 -0.8721 0 2.0 1e-06 
0.0 -0.872 0 2.0 1e-06 
0.0 -0.8719 0 2.0 1e-06 
0.0 -0.8718 0 2.0 1e-06 
0.0 -0.8717 0 2.0 1e-06 
0.0 -0.8716 0 2.0 1e-06 
0.0 -0.8715 0 2.0 1e-06 
0.0 -0.8714 0 2.0 1e-06 
0.0 -0.8713 0 2.0 1e-06 
0.0 -0.8712 0 2.0 1e-06 
0.0 -0.8711 0 2.0 1e-06 
0.0 -0.871 0 2.0 1e-06 
0.0 -0.8709 0 2.0 1e-06 
0.0 -0.8708 0 2.0 1e-06 
0.0 -0.8707 0 2.0 1e-06 
0.0 -0.8706 0 2.0 1e-06 
0.0 -0.8705 0 2.0 1e-06 
0.0 -0.8704 0 2.0 1e-06 
0.0 -0.8703 0 2.0 1e-06 
0.0 -0.8702 0 2.0 1e-06 
0.0 -0.8701 0 2.0 1e-06 
0.0 -0.87 0 2.0 1e-06 
0.0 -0.8699 0 2.0 1e-06 
0.0 -0.8698 0 2.0 1e-06 
0.0 -0.8697 0 2.0 1e-06 
0.0 -0.8696 0 2.0 1e-06 
0.0 -0.8695 0 2.0 1e-06 
0.0 -0.8694 0 2.0 1e-06 
0.0 -0.8693 0 2.0 1e-06 
0.0 -0.8692 0 2.0 1e-06 
0.0 -0.8691 0 2.0 1e-06 
0.0 -0.869 0 2.0 1e-06 
0.0 -0.8689 0 2.0 1e-06 
0.0 -0.8688 0 2.0 1e-06 
0.0 -0.8687 0 2.0 1e-06 
0.0 -0.8686 0 2.0 1e-06 
0.0 -0.8685 0 2.0 1e-06 
0.0 -0.8684 0 2.0 1e-06 
0.0 -0.8683 0 2.0 1e-06 
0.0 -0.8682 0 2.0 1e-06 
0.0 -0.8681 0 2.0 1e-06 
0.0 -0.868 0 2.0 1e-06 
0.0 -0.8679 0 2.0 1e-06 
0.0 -0.8678 0 2.0 1e-06 
0.0 -0.8677 0 2.0 1e-06 
0.0 -0.8676 0 2.0 1e-06 
0.0 -0.8675 0 2.0 1e-06 
0.0 -0.8674 0 2.0 1e-06 
0.0 -0.8673 0 2.0 1e-06 
0.0 -0.8672 0 2.0 1e-06 
0.0 -0.8671 0 2.0 1e-06 
0.0 -0.867 0 2.0 1e-06 
0.0 -0.8669 0 2.0 1e-06 
0.0 -0.8668 0 2.0 1e-06 
0.0 -0.8667 0 2.0 1e-06 
0.0 -0.8666 0 2.0 1e-06 
0.0 -0.8665 0 2.0 1e-06 
0.0 -0.8664 0 2.0 1e-06 
0.0 -0.8663 0 2.0 1e-06 
0.0 -0.8662 0 2.0 1e-06 
0.0 -0.8661 0 2.0 1e-06 
0.0 -0.866 0 2.0 1e-06 
0.0 -0.8659 0 2.0 1e-06 
0.0 -0.8658 0 2.0 1e-06 
0.0 -0.8657 0 2.0 1e-06 
0.0 -0.8656 0 2.0 1e-06 
0.0 -0.8655 0 2.0 1e-06 
0.0 -0.8654 0 2.0 1e-06 
0.0 -0.8653 0 2.0 1e-06 
0.0 -0.8652 0 2.0 1e-06 
0.0 -0.8651 0 2.0 1e-06 
0.0 -0.865 0 2.0 1e-06 
0.0 -0.8649 0 2.0 1e-06 
0.0 -0.8648 0 2.0 1e-06 
0.0 -0.8647 0 2.0 1e-06 
0.0 -0.8646 0 2.0 1e-06 
0.0 -0.8645 0 2.0 1e-06 
0.0 -0.8644 0 2.0 1e-06 
0.0 -0.8643 0 2.0 1e-06 
0.0 -0.8642 0 2.0 1e-06 
0.0 -0.8641 0 2.0 1e-06 
0.0 -0.864 0 2.0 1e-06 
0.0 -0.8639 0 2.0 1e-06 
0.0 -0.8638 0 2.0 1e-06 
0.0 -0.8637 0 2.0 1e-06 
0.0 -0.8636 0 2.0 1e-06 
0.0 -0.8635 0 2.0 1e-06 
0.0 -0.8634 0 2.0 1e-06 
0.0 -0.8633 0 2.0 1e-06 
0.0 -0.8632 0 2.0 1e-06 
0.0 -0.8631 0 2.0 1e-06 
0.0 -0.863 0 2.0 1e-06 
0.0 -0.8629 0 2.0 1e-06 
0.0 -0.8628 0 2.0 1e-06 
0.0 -0.8627 0 2.0 1e-06 
0.0 -0.8626 0 2.0 1e-06 
0.0 -0.8625 0 2.0 1e-06 
0.0 -0.8624 0 2.0 1e-06 
0.0 -0.8623 0 2.0 1e-06 
0.0 -0.8622 0 2.0 1e-06 
0.0 -0.8621 0 2.0 1e-06 
0.0 -0.862 0 2.0 1e-06 
0.0 -0.8619 0 2.0 1e-06 
0.0 -0.8618 0 2.0 1e-06 
0.0 -0.8617 0 2.0 1e-06 
0.0 -0.8616 0 2.0 1e-06 
0.0 -0.8615 0 2.0 1e-06 
0.0 -0.8614 0 2.0 1e-06 
0.0 -0.8613 0 2.0 1e-06 
0.0 -0.8612 0 2.0 1e-06 
0.0 -0.8611 0 2.0 1e-06 
0.0 -0.861 0 2.0 1e-06 
0.0 -0.8609 0 2.0 1e-06 
0.0 -0.8608 0 2.0 1e-06 
0.0 -0.8607 0 2.0 1e-06 
0.0 -0.8606 0 2.0 1e-06 
0.0 -0.8605 0 2.0 1e-06 
0.0 -0.8604 0 2.0 1e-06 
0.0 -0.8603 0 2.0 1e-06 
0.0 -0.8602 0 2.0 1e-06 
0.0 -0.8601 0 2.0 1e-06 
0.0 -0.86 0 2.0 1e-06 
0.0 -0.8599 0 2.0 1e-06 
0.0 -0.8598 0 2.0 1e-06 
0.0 -0.8597 0 2.0 1e-06 
0.0 -0.8596 0 2.0 1e-06 
0.0 -0.8595 0 2.0 1e-06 
0.0 -0.8594 0 2.0 1e-06 
0.0 -0.8593 0 2.0 1e-06 
0.0 -0.8592 0 2.0 1e-06 
0.0 -0.8591 0 2.0 1e-06 
0.0 -0.859 0 2.0 1e-06 
0.0 -0.8589 0 2.0 1e-06 
0.0 -0.8588 0 2.0 1e-06 
0.0 -0.8587 0 2.0 1e-06 
0.0 -0.8586 0 2.0 1e-06 
0.0 -0.8585 0 2.0 1e-06 
0.0 -0.8584 0 2.0 1e-06 
0.0 -0.8583 0 2.0 1e-06 
0.0 -0.8582 0 2.0 1e-06 
0.0 -0.8581 0 2.0 1e-06 
0.0 -0.858 0 2.0 1e-06 
0.0 -0.8579 0 2.0 1e-06 
0.0 -0.8578 0 2.0 1e-06 
0.0 -0.8577 0 2.0 1e-06 
0.0 -0.8576 0 2.0 1e-06 
0.0 -0.8575 0 2.0 1e-06 
0.0 -0.8574 0 2.0 1e-06 
0.0 -0.8573 0 2.0 1e-06 
0.0 -0.8572 0 2.0 1e-06 
0.0 -0.8571 0 2.0 1e-06 
0.0 -0.857 0 2.0 1e-06 
0.0 -0.8569 0 2.0 1e-06 
0.0 -0.8568 0 2.0 1e-06 
0.0 -0.8567 0 2.0 1e-06 
0.0 -0.8566 0 2.0 1e-06 
0.0 -0.8565 0 2.0 1e-06 
0.0 -0.8564 0 2.0 1e-06 
0.0 -0.8563 0 2.0 1e-06 
0.0 -0.8562 0 2.0 1e-06 
0.0 -0.8561 0 2.0 1e-06 
0.0 -0.856 0 2.0 1e-06 
0.0 -0.8559 0 2.0 1e-06 
0.0 -0.8558 0 2.0 1e-06 
0.0 -0.8557 0 2.0 1e-06 
0.0 -0.8556 0 2.0 1e-06 
0.0 -0.8555 0 2.0 1e-06 
0.0 -0.8554 0 2.0 1e-06 
0.0 -0.8553 0 2.0 1e-06 
0.0 -0.8552 0 2.0 1e-06 
0.0 -0.8551 0 2.0 1e-06 
0.0 -0.855 0 2.0 1e-06 
0.0 -0.8549 0 2.0 1e-06 
0.0 -0.8548 0 2.0 1e-06 
0.0 -0.8547 0 2.0 1e-06 
0.0 -0.8546 0 2.0 1e-06 
0.0 -0.8545 0 2.0 1e-06 
0.0 -0.8544 0 2.0 1e-06 
0.0 -0.8543 0 2.0 1e-06 
0.0 -0.8542 0 2.0 1e-06 
0.0 -0.8541 0 2.0 1e-06 
0.0 -0.854 0 2.0 1e-06 
0.0 -0.8539 0 2.0 1e-06 
0.0 -0.8538 0 2.0 1e-06 
0.0 -0.8537 0 2.0 1e-06 
0.0 -0.8536 0 2.0 1e-06 
0.0 -0.8535 0 2.0 1e-06 
0.0 -0.8534 0 2.0 1e-06 
0.0 -0.8533 0 2.0 1e-06 
0.0 -0.8532 0 2.0 1e-06 
0.0 -0.8531 0 2.0 1e-06 
0.0 -0.853 0 2.0 1e-06 
0.0 -0.8529 0 2.0 1e-06 
0.0 -0.8528 0 2.0 1e-06 
0.0 -0.8527 0 2.0 1e-06 
0.0 -0.8526 0 2.0 1e-06 
0.0 -0.8525 0 2.0 1e-06 
0.0 -0.8524 0 2.0 1e-06 
0.0 -0.8523 0 2.0 1e-06 
0.0 -0.8522 0 2.0 1e-06 
0.0 -0.8521 0 2.0 1e-06 
0.0 -0.852 0 2.0 1e-06 
0.0 -0.8519 0 2.0 1e-06 
0.0 -0.8518 0 2.0 1e-06 
0.0 -0.8517 0 2.0 1e-06 
0.0 -0.8516 0 2.0 1e-06 
0.0 -0.8515 0 2.0 1e-06 
0.0 -0.8514 0 2.0 1e-06 
0.0 -0.8513 0 2.0 1e-06 
0.0 -0.8512 0 2.0 1e-06 
0.0 -0.8511 0 2.0 1e-06 
0.0 -0.851 0 2.0 1e-06 
0.0 -0.8509 0 2.0 1e-06 
0.0 -0.8508 0 2.0 1e-06 
0.0 -0.8507 0 2.0 1e-06 
0.0 -0.8506 0 2.0 1e-06 
0.0 -0.8505 0 2.0 1e-06 
0.0 -0.8504 0 2.0 1e-06 
0.0 -0.8503 0 2.0 1e-06 
0.0 -0.8502 0 2.0 1e-06 
0.0 -0.8501 0 2.0 1e-06 
0.0 -0.85 0 2.0 1e-06 
0.0 -0.8499 0 2.0 1e-06 
0.0 -0.8498 0 2.0 1e-06 
0.0 -0.8497 0 2.0 1e-06 
0.0 -0.8496 0 2.0 1e-06 
0.0 -0.8495 0 2.0 1e-06 
0.0 -0.8494 0 2.0 1e-06 
0.0 -0.8493 0 2.0 1e-06 
0.0 -0.8492 0 2.0 1e-06 
0.0 -0.8491 0 2.0 1e-06 
0.0 -0.849 0 2.0 1e-06 
0.0 -0.8489 0 2.0 1e-06 
0.0 -0.8488 0 2.0 1e-06 
0.0 -0.8487 0 2.0 1e-06 
0.0 -0.8486 0 2.0 1e-06 
0.0 -0.8485 0 2.0 1e-06 
0.0 -0.8484 0 2.0 1e-06 
0.0 -0.8483 0 2.0 1e-06 
0.0 -0.8482 0 2.0 1e-06 
0.0 -0.8481 0 2.0 1e-06 
0.0 -0.848 0 2.0 1e-06 
0.0 -0.8479 0 2.0 1e-06 
0.0 -0.8478 0 2.0 1e-06 
0.0 -0.8477 0 2.0 1e-06 
0.0 -0.8476 0 2.0 1e-06 
0.0 -0.8475 0 2.0 1e-06 
0.0 -0.8474 0 2.0 1e-06 
0.0 -0.8473 0 2.0 1e-06 
0.0 -0.8472 0 2.0 1e-06 
0.0 -0.8471 0 2.0 1e-06 
0.0 -0.847 0 2.0 1e-06 
0.0 -0.8469 0 2.0 1e-06 
0.0 -0.8468 0 2.0 1e-06 
0.0 -0.8467 0 2.0 1e-06 
0.0 -0.8466 0 2.0 1e-06 
0.0 -0.8465 0 2.0 1e-06 
0.0 -0.8464 0 2.0 1e-06 
0.0 -0.8463 0 2.0 1e-06 
0.0 -0.8462 0 2.0 1e-06 
0.0 -0.8461 0 2.0 1e-06 
0.0 -0.846 0 2.0 1e-06 
0.0 -0.8459 0 2.0 1e-06 
0.0 -0.8458 0 2.0 1e-06 
0.0 -0.8457 0 2.0 1e-06 
0.0 -0.8456 0 2.0 1e-06 
0.0 -0.8455 0 2.0 1e-06 
0.0 -0.8454 0 2.0 1e-06 
0.0 -0.8453 0 2.0 1e-06 
0.0 -0.8452 0 2.0 1e-06 
0.0 -0.8451 0 2.0 1e-06 
0.0 -0.845 0 2.0 1e-06 
0.0 -0.8449 0 2.0 1e-06 
0.0 -0.8448 0 2.0 1e-06 
0.0 -0.8447 0 2.0 1e-06 
0.0 -0.8446 0 2.0 1e-06 
0.0 -0.8445 0 2.0 1e-06 
0.0 -0.8444 0 2.0 1e-06 
0.0 -0.8443 0 2.0 1e-06 
0.0 -0.8442 0 2.0 1e-06 
0.0 -0.8441 0 2.0 1e-06 
0.0 -0.844 0 2.0 1e-06 
0.0 -0.8439 0 2.0 1e-06 
0.0 -0.8438 0 2.0 1e-06 
0.0 -0.8437 0 2.0 1e-06 
0.0 -0.8436 0 2.0 1e-06 
0.0 -0.8435 0 2.0 1e-06 
0.0 -0.8434 0 2.0 1e-06 
0.0 -0.8433 0 2.0 1e-06 
0.0 -0.8432 0 2.0 1e-06 
0.0 -0.8431 0 2.0 1e-06 
0.0 -0.843 0 2.0 1e-06 
0.0 -0.8429 0 2.0 1e-06 
0.0 -0.8428 0 2.0 1e-06 
0.0 -0.8427 0 2.0 1e-06 
0.0 -0.8426 0 2.0 1e-06 
0.0 -0.8425 0 2.0 1e-06 
0.0 -0.8424 0 2.0 1e-06 
0.0 -0.8423 0 2.0 1e-06 
0.0 -0.8422 0 2.0 1e-06 
0.0 -0.8421 0 2.0 1e-06 
0.0 -0.842 0 2.0 1e-06 
0.0 -0.8419 0 2.0 1e-06 
0.0 -0.8418 0 2.0 1e-06 
0.0 -0.8417 0 2.0 1e-06 
0.0 -0.8416 0 2.0 1e-06 
0.0 -0.8415 0 2.0 1e-06 
0.0 -0.8414 0 2.0 1e-06 
0.0 -0.8413 0 2.0 1e-06 
0.0 -0.8412 0 2.0 1e-06 
0.0 -0.8411 0 2.0 1e-06 
0.0 -0.841 0 2.0 1e-06 
0.0 -0.8409 0 2.0 1e-06 
0.0 -0.8408 0 2.0 1e-06 
0.0 -0.8407 0 2.0 1e-06 
0.0 -0.8406 0 2.0 1e-06 
0.0 -0.8405 0 2.0 1e-06 
0.0 -0.8404 0 2.0 1e-06 
0.0 -0.8403 0 2.0 1e-06 
0.0 -0.8402 0 2.0 1e-06 
0.0 -0.8401 0 2.0 1e-06 
0.0 -0.84 0 2.0 1e-06 
0.0 -0.8399 0 2.0 1e-06 
0.0 -0.8398 0 2.0 1e-06 
0.0 -0.8397 0 2.0 1e-06 
0.0 -0.8396 0 2.0 1e-06 
0.0 -0.8395 0 2.0 1e-06 
0.0 -0.8394 0 2.0 1e-06 
0.0 -0.8393 0 2.0 1e-06 
0.0 -0.8392 0 2.0 1e-06 
0.0 -0.8391 0 2.0 1e-06 
0.0 -0.839 0 2.0 1e-06 
0.0 -0.8389 0 2.0 1e-06 
0.0 -0.8388 0 2.0 1e-06 
0.0 -0.8387 0 2.0 1e-06 
0.0 -0.8386 0 2.0 1e-06 
0.0 -0.8385 0 2.0 1e-06 
0.0 -0.8384 0 2.0 1e-06 
0.0 -0.8383 0 2.0 1e-06 
0.0 -0.8382 0 2.0 1e-06 
0.0 -0.8381 0 2.0 1e-06 
0.0 -0.838 0 2.0 1e-06 
0.0 -0.8379 0 2.0 1e-06 
0.0 -0.8378 0 2.0 1e-06 
0.0 -0.8377 0 2.0 1e-06 
0.0 -0.8376 0 2.0 1e-06 
0.0 -0.8375 0 2.0 1e-06 
0.0 -0.8374 0 2.0 1e-06 
0.0 -0.8373 0 2.0 1e-06 
0.0 -0.8372 0 2.0 1e-06 
0.0 -0.8371 0 2.0 1e-06 
0.0 -0.837 0 2.0 1e-06 
0.0 -0.8369 0 2.0 1e-06 
0.0 -0.8368 0 2.0 1e-06 
0.0 -0.8367 0 2.0 1e-06 
0.0 -0.8366 0 2.0 1e-06 
0.0 -0.8365 0 2.0 1e-06 
0.0 -0.8364 0 2.0 1e-06 
0.0 -0.8363 0 2.0 1e-06 
0.0 -0.8362 0 2.0 1e-06 
0.0 -0.8361 0 2.0 1e-06 
0.0 -0.836 0 2.0 1e-06 
0.0 -0.8359 0 2.0 1e-06 
0.0 -0.8358 0 2.0 1e-06 
0.0 -0.8357 0 2.0 1e-06 
0.0 -0.8356 0 2.0 1e-06 
0.0 -0.8355 0 2.0 1e-06 
0.0 -0.8354 0 2.0 1e-06 
0.0 -0.8353 0 2.0 1e-06 
0.0 -0.8352 0 2.0 1e-06 
0.0 -0.8351 0 2.0 1e-06 
0.0 -0.835 0 2.0 1e-06 
0.0 -0.8349 0 2.0 1e-06 
0.0 -0.8348 0 2.0 1e-06 
0.0 -0.8347 0 2.0 1e-06 
0.0 -0.8346 0 2.0 1e-06 
0.0 -0.8345 0 2.0 1e-06 
0.0 -0.8344 0 2.0 1e-06 
0.0 -0.8343 0 2.0 1e-06 
0.0 -0.8342 0 2.0 1e-06 
0.0 -0.8341 0 2.0 1e-06 
0.0 -0.834 0 2.0 1e-06 
0.0 -0.8339 0 2.0 1e-06 
0.0 -0.8338 0 2.0 1e-06 
0.0 -0.8337 0 2.0 1e-06 
0.0 -0.8336 0 2.0 1e-06 
0.0 -0.8335 0 2.0 1e-06 
0.0 -0.8334 0 2.0 1e-06 
0.0 -0.8333 0 2.0 1e-06 
0.0 -0.8332 0 2.0 1e-06 
0.0 -0.8331 0 2.0 1e-06 
0.0 -0.833 0 2.0 1e-06 
0.0 -0.8329 0 2.0 1e-06 
0.0 -0.8328 0 2.0 1e-06 
0.0 -0.8327 0 2.0 1e-06 
0.0 -0.8326 0 2.0 1e-06 
0.0 -0.8325 0 2.0 1e-06 
0.0 -0.8324 0 2.0 1e-06 
0.0 -0.8323 0 2.0 1e-06 
0.0 -0.8322 0 2.0 1e-06 
0.0 -0.8321 0 2.0 1e-06 
0.0 -0.832 0 2.0 1e-06 
0.0 -0.8319 0 2.0 1e-06 
0.0 -0.8318 0 2.0 1e-06 
0.0 -0.8317 0 2.0 1e-06 
0.0 -0.8316 0 2.0 1e-06 
0.0 -0.8315 0 2.0 1e-06 
0.0 -0.8314 0 2.0 1e-06 
0.0 -0.8313 0 2.0 1e-06 
0.0 -0.8312 0 2.0 1e-06 
0.0 -0.8311 0 2.0 1e-06 
0.0 -0.831 0 2.0 1e-06 
0.0 -0.8309 0 2.0 1e-06 
0.0 -0.8308 0 2.0 1e-06 
0.0 -0.8307 0 2.0 1e-06 
0.0 -0.8306 0 2.0 1e-06 
0.0 -0.8305 0 2.0 1e-06 
0.0 -0.8304 0 2.0 1e-06 
0.0 -0.8303 0 2.0 1e-06 
0.0 -0.8302 0 2.0 1e-06 
0.0 -0.8301 0 2.0 1e-06 
0.0 -0.83 0 2.0 1e-06 
0.0 -0.8299 0 2.0 1e-06 
0.0 -0.8298 0 2.0 1e-06 
0.0 -0.8297 0 2.0 1e-06 
0.0 -0.8296 0 2.0 1e-06 
0.0 -0.8295 0 2.0 1e-06 
0.0 -0.8294 0 2.0 1e-06 
0.0 -0.8293 0 2.0 1e-06 
0.0 -0.8292 0 2.0 1e-06 
0.0 -0.8291 0 2.0 1e-06 
0.0 -0.829 0 2.0 1e-06 
0.0 -0.8289 0 2.0 1e-06 
0.0 -0.8288 0 2.0 1e-06 
0.0 -0.8287 0 2.0 1e-06 
0.0 -0.8286 0 2.0 1e-06 
0.0 -0.8285 0 2.0 1e-06 
0.0 -0.8284 0 2.0 1e-06 
0.0 -0.8283 0 2.0 1e-06 
0.0 -0.8282 0 2.0 1e-06 
0.0 -0.8281 0 2.0 1e-06 
0.0 -0.828 0 2.0 1e-06 
0.0 -0.8279 0 2.0 1e-06 
0.0 -0.8278 0 2.0 1e-06 
0.0 -0.8277 0 2.0 1e-06 
0.0 -0.8276 0 2.0 1e-06 
0.0 -0.8275 0 2.0 1e-06 
0.0 -0.8274 0 2.0 1e-06 
0.0 -0.8273 0 2.0 1e-06 
0.0 -0.8272 0 2.0 1e-06 
0.0 -0.8271 0 2.0 1e-06 
0.0 -0.827 0 2.0 1e-06 
0.0 -0.8269 0 2.0 1e-06 
0.0 -0.8268 0 2.0 1e-06 
0.0 -0.8267 0 2.0 1e-06 
0.0 -0.8266 0 2.0 1e-06 
0.0 -0.8265 0 2.0 1e-06 
0.0 -0.8264 0 2.0 1e-06 
0.0 -0.8263 0 2.0 1e-06 
0.0 -0.8262 0 2.0 1e-06 
0.0 -0.8261 0 2.0 1e-06 
0.0 -0.826 0 2.0 1e-06 
0.0 -0.8259 0 2.0 1e-06 
0.0 -0.8258 0 2.0 1e-06 
0.0 -0.8257 0 2.0 1e-06 
0.0 -0.8256 0 2.0 1e-06 
0.0 -0.8255 0 2.0 1e-06 
0.0 -0.8254 0 2.0 1e-06 
0.0 -0.8253 0 2.0 1e-06 
0.0 -0.8252 0 2.0 1e-06 
0.0 -0.8251 0 2.0 1e-06 
0.0 -0.825 0 2.0 1e-06 
0.0 -0.8249 0 2.0 1e-06 
0.0 -0.8248 0 2.0 1e-06 
0.0 -0.8247 0 2.0 1e-06 
0.0 -0.8246 0 2.0 1e-06 
0.0 -0.8245 0 2.0 1e-06 
0.0 -0.8244 0 2.0 1e-06 
0.0 -0.8243 0 2.0 1e-06 
0.0 -0.8242 0 2.0 1e-06 
0.0 -0.8241 0 2.0 1e-06 
0.0 -0.824 0 2.0 1e-06 
0.0 -0.8239 0 2.0 1e-06 
0.0 -0.8238 0 2.0 1e-06 
0.0 -0.8237 0 2.0 1e-06 
0.0 -0.8236 0 2.0 1e-06 
0.0 -0.8235 0 2.0 1e-06 
0.0 -0.8234 0 2.0 1e-06 
0.0 -0.8233 0 2.0 1e-06 
0.0 -0.8232 0 2.0 1e-06 
0.0 -0.8231 0 2.0 1e-06 
0.0 -0.823 0 2.0 1e-06 
0.0 -0.8229 0 2.0 1e-06 
0.0 -0.8228 0 2.0 1e-06 
0.0 -0.8227 0 2.0 1e-06 
0.0 -0.8226 0 2.0 1e-06 
0.0 -0.8225 0 2.0 1e-06 
0.0 -0.8224 0 2.0 1e-06 
0.0 -0.8223 0 2.0 1e-06 
0.0 -0.8222 0 2.0 1e-06 
0.0 -0.8221 0 2.0 1e-06 
0.0 -0.822 0 2.0 1e-06 
0.0 -0.8219 0 2.0 1e-06 
0.0 -0.8218 0 2.0 1e-06 
0.0 -0.8217 0 2.0 1e-06 
0.0 -0.8216 0 2.0 1e-06 
0.0 -0.8215 0 2.0 1e-06 
0.0 -0.8214 0 2.0 1e-06 
0.0 -0.8213 0 2.0 1e-06 
0.0 -0.8212 0 2.0 1e-06 
0.0 -0.8211 0 2.0 1e-06 
0.0 -0.821 0 2.0 1e-06 
0.0 -0.8209 0 2.0 1e-06 
0.0 -0.8208 0 2.0 1e-06 
0.0 -0.8207 0 2.0 1e-06 
0.0 -0.8206 0 2.0 1e-06 
0.0 -0.8205 0 2.0 1e-06 
0.0 -0.8204 0 2.0 1e-06 
0.0 -0.8203 0 2.0 1e-06 
0.0 -0.8202 0 2.0 1e-06 
0.0 -0.8201 0 2.0 1e-06 
0.0 -0.82 0 2.0 1e-06 
0.0 -0.8199 0 2.0 1e-06 
0.0 -0.8198 0 2.0 1e-06 
0.0 -0.8197 0 2.0 1e-06 
0.0 -0.8196 0 2.0 1e-06 
0.0 -0.8195 0 2.0 1e-06 
0.0 -0.8194 0 2.0 1e-06 
0.0 -0.8193 0 2.0 1e-06 
0.0 -0.8192 0 2.0 1e-06 
0.0 -0.8191 0 2.0 1e-06 
0.0 -0.819 0 2.0 1e-06 
0.0 -0.8189 0 2.0 1e-06 
0.0 -0.8188 0 2.0 1e-06 
0.0 -0.8187 0 2.0 1e-06 
0.0 -0.8186 0 2.0 1e-06 
0.0 -0.8185 0 2.0 1e-06 
0.0 -0.8184 0 2.0 1e-06 
0.0 -0.8183 0 2.0 1e-06 
0.0 -0.8182 0 2.0 1e-06 
0.0 -0.8181 0 2.0 1e-06 
0.0 -0.818 0 2.0 1e-06 
0.0 -0.8179 0 2.0 1e-06 
0.0 -0.8178 0 2.0 1e-06 
0.0 -0.8177 0 2.0 1e-06 
0.0 -0.8176 0 2.0 1e-06 
0.0 -0.8175 0 2.0 1e-06 
0.0 -0.8174 0 2.0 1e-06 
0.0 -0.8173 0 2.0 1e-06 
0.0 -0.8172 0 2.0 1e-06 
0.0 -0.8171 0 2.0 1e-06 
0.0 -0.817 0 2.0 1e-06 
0.0 -0.8169 0 2.0 1e-06 
0.0 -0.8168 0 2.0 1e-06 
0.0 -0.8167 0 2.0 1e-06 
0.0 -0.8166 0 2.0 1e-06 
0.0 -0.8165 0 2.0 1e-06 
0.0 -0.8164 0 2.0 1e-06 
0.0 -0.8163 0 2.0 1e-06 
0.0 -0.8162 0 2.0 1e-06 
0.0 -0.8161 0 2.0 1e-06 
0.0 -0.816 0 2.0 1e-06 
0.0 -0.8159 0 2.0 1e-06 
0.0 -0.8158 0 2.0 1e-06 
0.0 -0.8157 0 2.0 1e-06 
0.0 -0.8156 0 2.0 1e-06 
0.0 -0.8155 0 2.0 1e-06 
0.0 -0.8154 0 2.0 1e-06 
0.0 -0.8153 0 2.0 1e-06 
0.0 -0.8152 0 2.0 1e-06 
0.0 -0.8151 0 2.0 1e-06 
0.0 -0.815 0 2.0 1e-06 
0.0 -0.8149 0 2.0 1e-06 
0.0 -0.8148 0 2.0 1e-06 
0.0 -0.8147 0 2.0 1e-06 
0.0 -0.8146 0 2.0 1e-06 
0.0 -0.8145 0 2.0 1e-06 
0.0 -0.8144 0 2.0 1e-06 
0.0 -0.8143 0 2.0 1e-06 
0.0 -0.8142 0 2.0 1e-06 
0.0 -0.8141 0 2.0 1e-06 
0.0 -0.814 0 2.0 1e-06 
0.0 -0.8139 0 2.0 1e-06 
0.0 -0.8138 0 2.0 1e-06 
0.0 -0.8137 0 2.0 1e-06 
0.0 -0.8136 0 2.0 1e-06 
0.0 -0.8135 0 2.0 1e-06 
0.0 -0.8134 0 2.0 1e-06 
0.0 -0.8133 0 2.0 1e-06 
0.0 -0.8132 0 2.0 1e-06 
0.0 -0.8131 0 2.0 1e-06 
0.0 -0.813 0 2.0 1e-06 
0.0 -0.8129 0 2.0 1e-06 
0.0 -0.8128 0 2.0 1e-06 
0.0 -0.8127 0 2.0 1e-06 
0.0 -0.8126 0 2.0 1e-06 
0.0 -0.8125 0 2.0 1e-06 
0.0 -0.8124 0 2.0 1e-06 
0.0 -0.8123 0 2.0 1e-06 
0.0 -0.8122 0 2.0 1e-06 
0.0 -0.8121 0 2.0 1e-06 
0.0 -0.812 0 2.0 1e-06 
0.0 -0.8119 0 2.0 1e-06 
0.0 -0.8118 0 2.0 1e-06 
0.0 -0.8117 0 2.0 1e-06 
0.0 -0.8116 0 2.0 1e-06 
0.0 -0.8115 0 2.0 1e-06 
0.0 -0.8114 0 2.0 1e-06 
0.0 -0.8113 0 2.0 1e-06 
0.0 -0.8112 0 2.0 1e-06 
0.0 -0.8111 0 2.0 1e-06 
0.0 -0.811 0 2.0 1e-06 
0.0 -0.8109 0 2.0 1e-06 
0.0 -0.8108 0 2.0 1e-06 
0.0 -0.8107 0 2.0 1e-06 
0.0 -0.8106 0 2.0 1e-06 
0.0 -0.8105 0 2.0 1e-06 
0.0 -0.8104 0 2.0 1e-06 
0.0 -0.8103 0 2.0 1e-06 
0.0 -0.8102 0 2.0 1e-06 
0.0 -0.8101 0 2.0 1e-06 
0.0 -0.81 0 2.0 1e-06 
0.0 -0.8099 0 2.0 1e-06 
0.0 -0.8098 0 2.0 1e-06 
0.0 -0.8097 0 2.0 1e-06 
0.0 -0.8096 0 2.0 1e-06 
0.0 -0.8095 0 2.0 1e-06 
0.0 -0.8094 0 2.0 1e-06 
0.0 -0.8093 0 2.0 1e-06 
0.0 -0.8092 0 2.0 1e-06 
0.0 -0.8091 0 2.0 1e-06 
0.0 -0.809 0 2.0 1e-06 
0.0 -0.8089 0 2.0 1e-06 
0.0 -0.8088 0 2.0 1e-06 
0.0 -0.8087 0 2.0 1e-06 
0.0 -0.8086 0 2.0 1e-06 
0.0 -0.8085 0 2.0 1e-06 
0.0 -0.8084 0 2.0 1e-06 
0.0 -0.8083 0 2.0 1e-06 
0.0 -0.8082 0 2.0 1e-06 
0.0 -0.8081 0 2.0 1e-06 
0.0 -0.808 0 2.0 1e-06 
0.0 -0.8079 0 2.0 1e-06 
0.0 -0.8078 0 2.0 1e-06 
0.0 -0.8077 0 2.0 1e-06 
0.0 -0.8076 0 2.0 1e-06 
0.0 -0.8075 0 2.0 1e-06 
0.0 -0.8074 0 2.0 1e-06 
0.0 -0.8073 0 2.0 1e-06 
0.0 -0.8072 0 2.0 1e-06 
0.0 -0.8071 0 2.0 1e-06 
0.0 -0.807 0 2.0 1e-06 
0.0 -0.8069 0 2.0 1e-06 
0.0 -0.8068 0 2.0 1e-06 
0.0 -0.8067 0 2.0 1e-06 
0.0 -0.8066 0 2.0 1e-06 
0.0 -0.8065 0 2.0 1e-06 
0.0 -0.8064 0 2.0 1e-06 
0.0 -0.8063 0 2.0 1e-06 
0.0 -0.8062 0 2.0 1e-06 
0.0 -0.8061 0 2.0 1e-06 
0.0 -0.806 0 2.0 1e-06 
0.0 -0.8059 0 2.0 1e-06 
0.0 -0.8058 0 2.0 1e-06 
0.0 -0.8057 0 2.0 1e-06 
0.0 -0.8056 0 2.0 1e-06 
0.0 -0.8055 0 2.0 1e-06 
0.0 -0.8054 0 2.0 1e-06 
0.0 -0.8053 0 2.0 1e-06 
0.0 -0.8052 0 2.0 1e-06 
0.0 -0.8051 0 2.0 1e-06 
0.0 -0.805 0 2.0 1e-06 
0.0 -0.8049 0 2.0 1e-06 
0.0 -0.8048 0 2.0 1e-06 
0.0 -0.8047 0 2.0 1e-06 
0.0 -0.8046 0 2.0 1e-06 
0.0 -0.8045 0 2.0 1e-06 
0.0 -0.8044 0 2.0 1e-06 
0.0 -0.8043 0 2.0 1e-06 
0.0 -0.8042 0 2.0 1e-06 
0.0 -0.8041 0 2.0 1e-06 
0.0 -0.804 0 2.0 1e-06 
0.0 -0.8039 0 2.0 1e-06 
0.0 -0.8038 0 2.0 1e-06 
0.0 -0.8037 0 2.0 1e-06 
0.0 -0.8036 0 2.0 1e-06 
0.0 -0.8035 0 2.0 1e-06 
0.0 -0.8034 0 2.0 1e-06 
0.0 -0.8033 0 2.0 1e-06 
0.0 -0.8032 0 2.0 1e-06 
0.0 -0.8031 0 2.0 1e-06 
0.0 -0.803 0 2.0 1e-06 
0.0 -0.8029 0 2.0 1e-06 
0.0 -0.8028 0 2.0 1e-06 
0.0 -0.8027 0 2.0 1e-06 
0.0 -0.8026 0 2.0 1e-06 
0.0 -0.8025 0 2.0 1e-06 
0.0 -0.8024 0 2.0 1e-06 
0.0 -0.8023 0 2.0 1e-06 
0.0 -0.8022 0 2.0 1e-06 
0.0 -0.8021 0 2.0 1e-06 
0.0 -0.802 0 2.0 1e-06 
0.0 -0.8019 0 2.0 1e-06 
0.0 -0.8018 0 2.0 1e-06 
0.0 -0.8017 0 2.0 1e-06 
0.0 -0.8016 0 2.0 1e-06 
0.0 -0.8015 0 2.0 1e-06 
0.0 -0.8014 0 2.0 1e-06 
0.0 -0.8013 0 2.0 1e-06 
0.0 -0.8012 0 2.0 1e-06 
0.0 -0.8011 0 2.0 1e-06 
0.0 -0.801 0 2.0 1e-06 
0.0 -0.8009 0 2.0 1e-06 
0.0 -0.8008 0 2.0 1e-06 
0.0 -0.8007 0 2.0 1e-06 
0.0 -0.8006 0 2.0 1e-06 
0.0 -0.8005 0 2.0 1e-06 
0.0 -0.8004 0 2.0 1e-06 
0.0 -0.8003 0 2.0 1e-06 
0.0 -0.8002 0 2.0 1e-06 
0.0 -0.8001 0 2.0 1e-06 
0.0 -0.8 0 2.0 1e-06 
0.0 -0.7999 0 2.0 1e-06 
0.0 -0.7998 0 2.0 1e-06 
0.0 -0.7997 0 2.0 1e-06 
0.0 -0.7996 0 2.0 1e-06 
0.0 -0.7995 0 2.0 1e-06 
0.0 -0.7994 0 2.0 1e-06 
0.0 -0.7993 0 2.0 1e-06 
0.0 -0.7992 0 2.0 1e-06 
0.0 -0.7991 0 2.0 1e-06 
0.0 -0.799 0 2.0 1e-06 
0.0 -0.7989 0 2.0 1e-06 
0.0 -0.7988 0 2.0 1e-06 
0.0 -0.7987 0 2.0 1e-06 
0.0 -0.7986 0 2.0 1e-06 
0.0 -0.7985 0 2.0 1e-06 
0.0 -0.7984 0 2.0 1e-06 
0.0 -0.7983 0 2.0 1e-06 
0.0 -0.7982 0 2.0 1e-06 
0.0 -0.7981 0 2.0 1e-06 
0.0 -0.798 0 2.0 1e-06 
0.0 -0.7979 0 2.0 1e-06 
0.0 -0.7978 0 2.0 1e-06 
0.0 -0.7977 0 2.0 1e-06 
0.0 -0.7976 0 2.0 1e-06 
0.0 -0.7975 0 2.0 1e-06 
0.0 -0.7974 0 2.0 1e-06 
0.0 -0.7973 0 2.0 1e-06 
0.0 -0.7972 0 2.0 1e-06 
0.0 -0.7971 0 2.0 1e-06 
0.0 -0.797 0 2.0 1e-06 
0.0 -0.7969 0 2.0 1e-06 
0.0 -0.7968 0 2.0 1e-06 
0.0 -0.7967 0 2.0 1e-06 
0.0 -0.7966 0 2.0 1e-06 
0.0 -0.7965 0 2.0 1e-06 
0.0 -0.7964 0 2.0 1e-06 
0.0 -0.7963 0 2.0 1e-06 
0.0 -0.7962 0 2.0 1e-06 
0.0 -0.7961 0 2.0 1e-06 
0.0 -0.796 0 2.0 1e-06 
0.0 -0.7959 0 2.0 1e-06 
0.0 -0.7958 0 2.0 1e-06 
0.0 -0.7957 0 2.0 1e-06 
0.0 -0.7956 0 2.0 1e-06 
0.0 -0.7955 0 2.0 1e-06 
0.0 -0.7954 0 2.0 1e-06 
0.0 -0.7953 0 2.0 1e-06 
0.0 -0.7952 0 2.0 1e-06 
0.0 -0.7951 0 2.0 1e-06 
0.0 -0.795 0 2.0 1e-06 
0.0 -0.7949 0 2.0 1e-06 
0.0 -0.7948 0 2.0 1e-06 
0.0 -0.7947 0 2.0 1e-06 
0.0 -0.7946 0 2.0 1e-06 
0.0 -0.7945 0 2.0 1e-06 
0.0 -0.7944 0 2.0 1e-06 
0.0 -0.7943 0 2.0 1e-06 
0.0 -0.7942 0 2.0 1e-06 
0.0 -0.7941 0 2.0 1e-06 
0.0 -0.794 0 2.0 1e-06 
0.0 -0.7939 0 2.0 1e-06 
0.0 -0.7938 0 2.0 1e-06 
0.0 -0.7937 0 2.0 1e-06 
0.0 -0.7936 0 2.0 1e-06 
0.0 -0.7935 0 2.0 1e-06 
0.0 -0.7934 0 2.0 1e-06 
0.0 -0.7933 0 2.0 1e-06 
0.0 -0.7932 0 2.0 1e-06 
0.0 -0.7931 0 2.0 1e-06 
0.0 -0.793 0 2.0 1e-06 
0.0 -0.7929 0 2.0 1e-06 
0.0 -0.7928 0 2.0 1e-06 
0.0 -0.7927 0 2.0 1e-06 
0.0 -0.7926 0 2.0 1e-06 
0.0 -0.7925 0 2.0 1e-06 
0.0 -0.7924 0 2.0 1e-06 
0.0 -0.7923 0 2.0 1e-06 
0.0 -0.7922 0 2.0 1e-06 
0.0 -0.7921 0 2.0 1e-06 
0.0 -0.792 0 2.0 1e-06 
0.0 -0.7919 0 2.0 1e-06 
0.0 -0.7918 0 2.0 1e-06 
0.0 -0.7917 0 2.0 1e-06 
0.0 -0.7916 0 2.0 1e-06 
0.0 -0.7915 0 2.0 1e-06 
0.0 -0.7914 0 2.0 1e-06 
0.0 -0.7913 0 2.0 1e-06 
0.0 -0.7912 0 2.0 1e-06 
0.0 -0.7911 0 2.0 1e-06 
0.0 -0.791 0 2.0 1e-06 
0.0 -0.7909 0 2.0 1e-06 
0.0 -0.7908 0 2.0 1e-06 
0.0 -0.7907 0 2.0 1e-06 
0.0 -0.7906 0 2.0 1e-06 
0.0 -0.7905 0 2.0 1e-06 
0.0 -0.7904 0 2.0 1e-06 
0.0 -0.7903 0 2.0 1e-06 
0.0 -0.7902 0 2.0 1e-06 
0.0 -0.7901 0 2.0 1e-06 
0.0 -0.79 0 2.0 1e-06 
0.0 -0.7899 0 2.0 1e-06 
0.0 -0.7898 0 2.0 1e-06 
0.0 -0.7897 0 2.0 1e-06 
0.0 -0.7896 0 2.0 1e-06 
0.0 -0.7895 0 2.0 1e-06 
0.0 -0.7894 0 2.0 1e-06 
0.0 -0.7893 0 2.0 1e-06 
0.0 -0.7892 0 2.0 1e-06 
0.0 -0.7891 0 2.0 1e-06 
0.0 -0.789 0 2.0 1e-06 
0.0 -0.7889 0 2.0 1e-06 
0.0 -0.7888 0 2.0 1e-06 
0.0 -0.7887 0 2.0 1e-06 
0.0 -0.7886 0 2.0 1e-06 
0.0 -0.7885 0 2.0 1e-06 
0.0 -0.7884 0 2.0 1e-06 
0.0 -0.7883 0 2.0 1e-06 
0.0 -0.7882 0 2.0 1e-06 
0.0 -0.7881 0 2.0 1e-06 
0.0 -0.788 0 2.0 1e-06 
0.0 -0.7879 0 2.0 1e-06 
0.0 -0.7878 0 2.0 1e-06 
0.0 -0.7877 0 2.0 1e-06 
0.0 -0.7876 0 2.0 1e-06 
0.0 -0.7875 0 2.0 1e-06 
0.0 -0.7874 0 2.0 1e-06 
0.0 -0.7873 0 2.0 1e-06 
0.0 -0.7872 0 2.0 1e-06 
0.0 -0.7871 0 2.0 1e-06 
0.0 -0.787 0 2.0 1e-06 
0.0 -0.7869 0 2.0 1e-06 
0.0 -0.7868 0 2.0 1e-06 
0.0 -0.7867 0 2.0 1e-06 
0.0 -0.7866 0 2.0 1e-06 
0.0 -0.7865 0 2.0 1e-06 
0.0 -0.7864 0 2.0 1e-06 
0.0 -0.7863 0 2.0 1e-06 
0.0 -0.7862 0 2.0 1e-06 
0.0 -0.7861 0 2.0 1e-06 
0.0 -0.786 0 2.0 1e-06 
0.0 -0.7859 0 2.0 1e-06 
0.0 -0.7858 0 2.0 1e-06 
0.0 -0.7857 0 2.0 1e-06 
0.0 -0.7856 0 2.0 1e-06 
0.0 -0.7855 0 2.0 1e-06 
0.0 -0.7854 0 2.0 1e-06 
0.0 -0.7853 0 2.0 1e-06 
0.0 -0.7852 0 2.0 1e-06 
0.0 -0.7851 0 2.0 1e-06 
0.0 -0.785 0 2.0 1e-06 
0.0 -0.7849 0 2.0 1e-06 
0.0 -0.7848 0 2.0 1e-06 
0.0 -0.7847 0 2.0 1e-06 
0.0 -0.7846 0 2.0 1e-06 
0.0 -0.7845 0 2.0 1e-06 
0.0 -0.7844 0 2.0 1e-06 
0.0 -0.7843 0 2.0 1e-06 
0.0 -0.7842 0 2.0 1e-06 
0.0 -0.7841 0 2.0 1e-06 
0.0 -0.784 0 2.0 1e-06 
0.0 -0.7839 0 2.0 1e-06 
0.0 -0.7838 0 2.0 1e-06 
0.0 -0.7837 0 2.0 1e-06 
0.0 -0.7836 0 2.0 1e-06 
0.0 -0.7835 0 2.0 1e-06 
0.0 -0.7834 0 2.0 1e-06 
0.0 -0.7833 0 2.0 1e-06 
0.0 -0.7832 0 2.0 1e-06 
0.0 -0.7831 0 2.0 1e-06 
0.0 -0.783 0 2.0 1e-06 
0.0 -0.7829 0 2.0 1e-06 
0.0 -0.7828 0 2.0 1e-06 
0.0 -0.7827 0 2.0 1e-06 
0.0 -0.7826 0 2.0 1e-06 
0.0 -0.7825 0 2.0 1e-06 
0.0 -0.7824 0 2.0 1e-06 
0.0 -0.7823 0 2.0 1e-06 
0.0 -0.7822 0 2.0 1e-06 
0.0 -0.7821 0 2.0 1e-06 
0.0 -0.782 0 2.0 1e-06 
0.0 -0.7819 0 2.0 1e-06 
0.0 -0.7818 0 2.0 1e-06 
0.0 -0.7817 0 2.0 1e-06 
0.0 -0.7816 0 2.0 1e-06 
0.0 -0.7815 0 2.0 1e-06 
0.0 -0.7814 0 2.0 1e-06 
0.0 -0.7813 0 2.0 1e-06 
0.0 -0.7812 0 2.0 1e-06 
0.0 -0.7811 0 2.0 1e-06 
0.0 -0.781 0 2.0 1e-06 
0.0 -0.7809 0 2.0 1e-06 
0.0 -0.7808 0 2.0 1e-06 
0.0 -0.7807 0 2.0 1e-06 
0.0 -0.7806 0 2.0 1e-06 
0.0 -0.7805 0 2.0 1e-06 
0.0 -0.7804 0 2.0 1e-06 
0.0 -0.7803 0 2.0 1e-06 
0.0 -0.7802 0 2.0 1e-06 
0.0 -0.7801 0 2.0 1e-06 
0.0 -0.78 0 2.0 1e-06 
0.0 -0.7799 0 2.0 1e-06 
0.0 -0.7798 0 2.0 1e-06 
0.0 -0.7797 0 2.0 1e-06 
0.0 -0.7796 0 2.0 1e-06 
0.0 -0.7795 0 2.0 1e-06 
0.0 -0.7794 0 2.0 1e-06 
0.0 -0.7793 0 2.0 1e-06 
0.0 -0.7792 0 2.0 1e-06 
0.0 -0.7791 0 2.0 1e-06 
0.0 -0.779 0 2.0 1e-06 
0.0 -0.7789 0 2.0 1e-06 
0.0 -0.7788 0 2.0 1e-06 
0.0 -0.7787 0 2.0 1e-06 
0.0 -0.7786 0 2.0 1e-06 
0.0 -0.7785 0 2.0 1e-06 
0.0 -0.7784 0 2.0 1e-06 
0.0 -0.7783 0 2.0 1e-06 
0.0 -0.7782 0 2.0 1e-06 
0.0 -0.7781 0 2.0 1e-06 
0.0 -0.778 0 2.0 1e-06 
0.0 -0.7779 0 2.0 1e-06 
0.0 -0.7778 0 2.0 1e-06 
0.0 -0.7777 0 2.0 1e-06 
0.0 -0.7776 0 2.0 1e-06 
0.0 -0.7775 0 2.0 1e-06 
0.0 -0.7774 0 2.0 1e-06 
0.0 -0.7773 0 2.0 1e-06 
0.0 -0.7772 0 2.0 1e-06 
0.0 -0.7771 0 2.0 1e-06 
0.0 -0.777 0 2.0 1e-06 
0.0 -0.7769 0 2.0 1e-06 
0.0 -0.7768 0 2.0 1e-06 
0.0 -0.7767 0 2.0 1e-06 
0.0 -0.7766 0 2.0 1e-06 
0.0 -0.7765 0 2.0 1e-06 
0.0 -0.7764 0 2.0 1e-06 
0.0 -0.7763 0 2.0 1e-06 
0.0 -0.7762 0 2.0 1e-06 
0.0 -0.7761 0 2.0 1e-06 
0.0 -0.776 0 2.0 1e-06 
0.0 -0.7759 0 2.0 1e-06 
0.0 -0.7758 0 2.0 1e-06 
0.0 -0.7757 0 2.0 1e-06 
0.0 -0.7756 0 2.0 1e-06 
0.0 -0.7755 0 2.0 1e-06 
0.0 -0.7754 0 2.0 1e-06 
0.0 -0.7753 0 2.0 1e-06 
0.0 -0.7752 0 2.0 1e-06 
0.0 -0.7751 0 2.0 1e-06 
0.0 -0.775 0 2.0 1e-06 
0.0 -0.7749 0 2.0 1e-06 
0.0 -0.7748 0 2.0 1e-06 
0.0 -0.7747 0 2.0 1e-06 
0.0 -0.7746 0 2.0 1e-06 
0.0 -0.7745 0 2.0 1e-06 
0.0 -0.7744 0 2.0 1e-06 
0.0 -0.7743 0 2.0 1e-06 
0.0 -0.7742 0 2.0 1e-06 
0.0 -0.7741 0 2.0 1e-06 
0.0 -0.774 0 2.0 1e-06 
0.0 -0.7739 0 2.0 1e-06 
0.0 -0.7738 0 2.0 1e-06 
0.0 -0.7737 0 2.0 1e-06 
0.0 -0.7736 0 2.0 1e-06 
0.0 -0.7735 0 2.0 1e-06 
0.0 -0.7734 0 2.0 1e-06 
0.0 -0.7733 0 2.0 1e-06 
0.0 -0.7732 0 2.0 1e-06 
0.0 -0.7731 0 2.0 1e-06 
0.0 -0.773 0 2.0 1e-06 
0.0 -0.7729 0 2.0 1e-06 
0.0 -0.7728 0 2.0 1e-06 
0.0 -0.7727 0 2.0 1e-06 
0.0 -0.7726 0 2.0 1e-06 
0.0 -0.7725 0 2.0 1e-06 
0.0 -0.7724 0 2.0 1e-06 
0.0 -0.7723 0 2.0 1e-06 
0.0 -0.7722 0 2.0 1e-06 
0.0 -0.7721 0 2.0 1e-06 
0.0 -0.772 0 2.0 1e-06 
0.0 -0.7719 0 2.0 1e-06 
0.0 -0.7718 0 2.0 1e-06 
0.0 -0.7717 0 2.0 1e-06 
0.0 -0.7716 0 2.0 1e-06 
0.0 -0.7715 0 2.0 1e-06 
0.0 -0.7714 0 2.0 1e-06 
0.0 -0.7713 0 2.0 1e-06 
0.0 -0.7712 0 2.0 1e-06 
0.0 -0.7711 0 2.0 1e-06 
0.0 -0.771 0 2.0 1e-06 
0.0 -0.7709 0 2.0 1e-06 
0.0 -0.7708 0 2.0 1e-06 
0.0 -0.7707 0 2.0 1e-06 
0.0 -0.7706 0 2.0 1e-06 
0.0 -0.7705 0 2.0 1e-06 
0.0 -0.7704 0 2.0 1e-06 
0.0 -0.7703 0 2.0 1e-06 
0.0 -0.7702 0 2.0 1e-06 
0.0 -0.7701 0 2.0 1e-06 
0.0 -0.77 0 2.0 1e-06 
0.0 -0.7699 0 2.0 1e-06 
0.0 -0.7698 0 2.0 1e-06 
0.0 -0.7697 0 2.0 1e-06 
0.0 -0.7696 0 2.0 1e-06 
0.0 -0.7695 0 2.0 1e-06 
0.0 -0.7694 0 2.0 1e-06 
0.0 -0.7693 0 2.0 1e-06 
0.0 -0.7692 0 2.0 1e-06 
0.0 -0.7691 0 2.0 1e-06 
0.0 -0.769 0 2.0 1e-06 
0.0 -0.7689 0 2.0 1e-06 
0.0 -0.7688 0 2.0 1e-06 
0.0 -0.7687 0 2.0 1e-06 
0.0 -0.7686 0 2.0 1e-06 
0.0 -0.7685 0 2.0 1e-06 
0.0 -0.7684 0 2.0 1e-06 
0.0 -0.7683 0 2.0 1e-06 
0.0 -0.7682 0 2.0 1e-06 
0.0 -0.7681 0 2.0 1e-06 
0.0 -0.768 0 2.0 1e-06 
0.0 -0.7679 0 2.0 1e-06 
0.0 -0.7678 0 2.0 1e-06 
0.0 -0.7677 0 2.0 1e-06 
0.0 -0.7676 0 2.0 1e-06 
0.0 -0.7675 0 2.0 1e-06 
0.0 -0.7674 0 2.0 1e-06 
0.0 -0.7673 0 2.0 1e-06 
0.0 -0.7672 0 2.0 1e-06 
0.0 -0.7671 0 2.0 1e-06 
0.0 -0.767 0 2.0 1e-06 
0.0 -0.7669 0 2.0 1e-06 
0.0 -0.7668 0 2.0 1e-06 
0.0 -0.7667 0 2.0 1e-06 
0.0 -0.7666 0 2.0 1e-06 
0.0 -0.7665 0 2.0 1e-06 
0.0 -0.7664 0 2.0 1e-06 
0.0 -0.7663 0 2.0 1e-06 
0.0 -0.7662 0 2.0 1e-06 
0.0 -0.7661 0 2.0 1e-06 
0.0 -0.766 0 2.0 1e-06 
0.0 -0.7659 0 2.0 1e-06 
0.0 -0.7658 0 2.0 1e-06 
0.0 -0.7657 0 2.0 1e-06 
0.0 -0.7656 0 2.0 1e-06 
0.0 -0.7655 0 2.0 1e-06 
0.0 -0.7654 0 2.0 1e-06 
0.0 -0.7653 0 2.0 1e-06 
0.0 -0.7652 0 2.0 1e-06 
0.0 -0.7651 0 2.0 1e-06 
0.0 -0.765 0 2.0 1e-06 
0.0 -0.7649 0 2.0 1e-06 
0.0 -0.7648 0 2.0 1e-06 
0.0 -0.7647 0 2.0 1e-06 
0.0 -0.7646 0 2.0 1e-06 
0.0 -0.7645 0 2.0 1e-06 
0.0 -0.7644 0 2.0 1e-06 
0.0 -0.7643 0 2.0 1e-06 
0.0 -0.7642 0 2.0 1e-06 
0.0 -0.7641 0 2.0 1e-06 
0.0 -0.764 0 2.0 1e-06 
0.0 -0.7639 0 2.0 1e-06 
0.0 -0.7638 0 2.0 1e-06 
0.0 -0.7637 0 2.0 1e-06 
0.0 -0.7636 0 2.0 1e-06 
0.0 -0.7635 0 2.0 1e-06 
0.0 -0.7634 0 2.0 1e-06 
0.0 -0.7633 0 2.0 1e-06 
0.0 -0.7632 0 2.0 1e-06 
0.0 -0.7631 0 2.0 1e-06 
0.0 -0.763 0 2.0 1e-06 
0.0 -0.7629 0 2.0 1e-06 
0.0 -0.7628 0 2.0 1e-06 
0.0 -0.7627 0 2.0 1e-06 
0.0 -0.7626 0 2.0 1e-06 
0.0 -0.7625 0 2.0 1e-06 
0.0 -0.7624 0 2.0 1e-06 
0.0 -0.7623 0 2.0 1e-06 
0.0 -0.7622 0 2.0 1e-06 
0.0 -0.7621 0 2.0 1e-06 
0.0 -0.762 0 2.0 1e-06 
0.0 -0.7619 0 2.0 1e-06 
0.0 -0.7618 0 2.0 1e-06 
0.0 -0.7617 0 2.0 1e-06 
0.0 -0.7616 0 2.0 1e-06 
0.0 -0.7615 0 2.0 1e-06 
0.0 -0.7614 0 2.0 1e-06 
0.0 -0.7613 0 2.0 1e-06 
0.0 -0.7612 0 2.0 1e-06 
0.0 -0.7611 0 2.0 1e-06 
0.0 -0.761 0 2.0 1e-06 
0.0 -0.7609 0 2.0 1e-06 
0.0 -0.7608 0 2.0 1e-06 
0.0 -0.7607 0 2.0 1e-06 
0.0 -0.7606 0 2.0 1e-06 
0.0 -0.7605 0 2.0 1e-06 
0.0 -0.7604 0 2.0 1e-06 
0.0 -0.7603 0 2.0 1e-06 
0.0 -0.7602 0 2.0 1e-06 
0.0 -0.7601 0 2.0 1e-06 
0.0 -0.76 0 2.0 1e-06 
0.0 -0.7599 0 2.0 1e-06 
0.0 -0.7598 0 2.0 1e-06 
0.0 -0.7597 0 2.0 1e-06 
0.0 -0.7596 0 2.0 1e-06 
0.0 -0.7595 0 2.0 1e-06 
0.0 -0.7594 0 2.0 1e-06 
0.0 -0.7593 0 2.0 1e-06 
0.0 -0.7592 0 2.0 1e-06 
0.0 -0.7591 0 2.0 1e-06 
0.0 -0.759 0 2.0 1e-06 
0.0 -0.7589 0 2.0 1e-06 
0.0 -0.7588 0 2.0 1e-06 
0.0 -0.7587 0 2.0 1e-06 
0.0 -0.7586 0 2.0 1e-06 
0.0 -0.7585 0 2.0 1e-06 
0.0 -0.7584 0 2.0 1e-06 
0.0 -0.7583 0 2.0 1e-06 
0.0 -0.7582 0 2.0 1e-06 
0.0 -0.7581 0 2.0 1e-06 
0.0 -0.758 0 2.0 1e-06 
0.0 -0.7579 0 2.0 1e-06 
0.0 -0.7578 0 2.0 1e-06 
0.0 -0.7577 0 2.0 1e-06 
0.0 -0.7576 0 2.0 1e-06 
0.0 -0.7575 0 2.0 1e-06 
0.0 -0.7574 0 2.0 1e-06 
0.0 -0.7573 0 2.0 1e-06 
0.0 -0.7572 0 2.0 1e-06 
0.0 -0.7571 0 2.0 1e-06 
0.0 -0.757 0 2.0 1e-06 
0.0 -0.7569 0 2.0 1e-06 
0.0 -0.7568 0 2.0 1e-06 
0.0 -0.7567 0 2.0 1e-06 
0.0 -0.7566 0 2.0 1e-06 
0.0 -0.7565 0 2.0 1e-06 
0.0 -0.7564 0 2.0 1e-06 
0.0 -0.7563 0 2.0 1e-06 
0.0 -0.7562 0 2.0 1e-06 
0.0 -0.7561 0 2.0 1e-06 
0.0 -0.756 0 2.0 1e-06 
0.0 -0.7559 0 2.0 1e-06 
0.0 -0.7558 0 2.0 1e-06 
0.0 -0.7557 0 2.0 1e-06 
0.0 -0.7556 0 2.0 1e-06 
0.0 -0.7555 0 2.0 1e-06 
0.0 -0.7554 0 2.0 1e-06 
0.0 -0.7553 0 2.0 1e-06 
0.0 -0.7552 0 2.0 1e-06 
0.0 -0.7551 0 2.0 1e-06 
0.0 -0.755 0 2.0 1e-06 
0.0 -0.7549 0 2.0 1e-06 
0.0 -0.7548 0 2.0 1e-06 
0.0 -0.7547 0 2.0 1e-06 
0.0 -0.7546 0 2.0 1e-06 
0.0 -0.7545 0 2.0 1e-06 
0.0 -0.7544 0 2.0 1e-06 
0.0 -0.7543 0 2.0 1e-06 
0.0 -0.7542 0 2.0 1e-06 
0.0 -0.7541 0 2.0 1e-06 
0.0 -0.754 0 2.0 1e-06 
0.0 -0.7539 0 2.0 1e-06 
0.0 -0.7538 0 2.0 1e-06 
0.0 -0.7537 0 2.0 1e-06 
0.0 -0.7536 0 2.0 1e-06 
0.0 -0.7535 0 2.0 1e-06 
0.0 -0.7534 0 2.0 1e-06 
0.0 -0.7533 0 2.0 1e-06 
0.0 -0.7532 0 2.0 1e-06 
0.0 -0.7531 0 2.0 1e-06 
0.0 -0.753 0 2.0 1e-06 
0.0 -0.7529 0 2.0 1e-06 
0.0 -0.7528 0 2.0 1e-06 
0.0 -0.7527 0 2.0 1e-06 
0.0 -0.7526 0 2.0 1e-06 
0.0 -0.7525 0 2.0 1e-06 
0.0 -0.7524 0 2.0 1e-06 
0.0 -0.7523 0 2.0 1e-06 
0.0 -0.7522 0 2.0 1e-06 
0.0 -0.7521 0 2.0 1e-06 
0.0 -0.752 0 2.0 1e-06 
0.0 -0.7519 0 2.0 1e-06 
0.0 -0.7518 0 2.0 1e-06 
0.0 -0.7517 0 2.0 1e-06 
0.0 -0.7516 0 2.0 1e-06 
0.0 -0.7515 0 2.0 1e-06 
0.0 -0.7514 0 2.0 1e-06 
0.0 -0.7513 0 2.0 1e-06 
0.0 -0.7512 0 2.0 1e-06 
0.0 -0.7511 0 2.0 1e-06 
0.0 -0.751 0 2.0 1e-06 
0.0 -0.7509 0 2.0 1e-06 
0.0 -0.7508 0 2.0 1e-06 
0.0 -0.7507 0 2.0 1e-06 
0.0 -0.7506 0 2.0 1e-06 
0.0 -0.7505 0 2.0 1e-06 
0.0 -0.7504 0 2.0 1e-06 
0.0 -0.7503 0 2.0 1e-06 
0.0 -0.7502 0 2.0 1e-06 
0.0 -0.7501 0 2.0 1e-06 
0.0 -0.75 0 2.0 1e-06 
0.0 -0.7499 0 2.0 1e-06 
0.0 -0.7498 0 2.0 1e-06 
0.0 -0.7497 0 2.0 1e-06 
0.0 -0.7496 0 2.0 1e-06 
0.0 -0.7495 0 2.0 1e-06 
0.0 -0.7494 0 2.0 1e-06 
0.0 -0.7493 0 2.0 1e-06 
0.0 -0.7492 0 2.0 1e-06 
0.0 -0.7491 0 2.0 1e-06 
0.0 -0.749 0 2.0 1e-06 
0.0 -0.7489 0 2.0 1e-06 
0.0 -0.7488 0 2.0 1e-06 
0.0 -0.7487 0 2.0 1e-06 
0.0 -0.7486 0 2.0 1e-06 
0.0 -0.7485 0 2.0 1e-06 
0.0 -0.7484 0 2.0 1e-06 
0.0 -0.7483 0 2.0 1e-06 
0.0 -0.7482 0 2.0 1e-06 
0.0 -0.7481 0 2.0 1e-06 
0.0 -0.748 0 2.0 1e-06 
0.0 -0.7479 0 2.0 1e-06 
0.0 -0.7478 0 2.0 1e-06 
0.0 -0.7477 0 2.0 1e-06 
0.0 -0.7476 0 2.0 1e-06 
0.0 -0.7475 0 2.0 1e-06 
0.0 -0.7474 0 2.0 1e-06 
0.0 -0.7473 0 2.0 1e-06 
0.0 -0.7472 0 2.0 1e-06 
0.0 -0.7471 0 2.0 1e-06 
0.0 -0.747 0 2.0 1e-06 
0.0 -0.7469 0 2.0 1e-06 
0.0 -0.7468 0 2.0 1e-06 
0.0 -0.7467 0 2.0 1e-06 
0.0 -0.7466 0 2.0 1e-06 
0.0 -0.7465 0 2.0 1e-06 
0.0 -0.7464 0 2.0 1e-06 
0.0 -0.7463 0 2.0 1e-06 
0.0 -0.7462 0 2.0 1e-06 
0.0 -0.7461 0 2.0 1e-06 
0.0 -0.746 0 2.0 1e-06 
0.0 -0.7459 0 2.0 1e-06 
0.0 -0.7458 0 2.0 1e-06 
0.0 -0.7457 0 2.0 1e-06 
0.0 -0.7456 0 2.0 1e-06 
0.0 -0.7455 0 2.0 1e-06 
0.0 -0.7454 0 2.0 1e-06 
0.0 -0.7453 0 2.0 1e-06 
0.0 -0.7452 0 2.0 1e-06 
0.0 -0.7451 0 2.0 1e-06 
0.0 -0.745 0 2.0 1e-06 
0.0 -0.7449 0 2.0 1e-06 
0.0 -0.7448 0 2.0 1e-06 
0.0 -0.7447 0 2.0 1e-06 
0.0 -0.7446 0 2.0 1e-06 
0.0 -0.7445 0 2.0 1e-06 
0.0 -0.7444 0 2.0 1e-06 
0.0 -0.7443 0 2.0 1e-06 
0.0 -0.7442 0 2.0 1e-06 
0.0 -0.7441 0 2.0 1e-06 
0.0 -0.744 0 2.0 1e-06 
0.0 -0.7439 0 2.0 1e-06 
0.0 -0.7438 0 2.0 1e-06 
0.0 -0.7437 0 2.0 1e-06 
0.0 -0.7436 0 2.0 1e-06 
0.0 -0.7435 0 2.0 1e-06 
0.0 -0.7434 0 2.0 1e-06 
0.0 -0.7433 0 2.0 1e-06 
0.0 -0.7432 0 2.0 1e-06 
0.0 -0.7431 0 2.0 1e-06 
0.0 -0.743 0 2.0 1e-06 
0.0 -0.7429 0 2.0 1e-06 
0.0 -0.7428 0 2.0 1e-06 
0.0 -0.7427 0 2.0 1e-06 
0.0 -0.7426 0 2.0 1e-06 
0.0 -0.7425 0 2.0 1e-06 
0.0 -0.7424 0 2.0 1e-06 
0.0 -0.7423 0 2.0 1e-06 
0.0 -0.7422 0 2.0 1e-06 
0.0 -0.7421 0 2.0 1e-06 
0.0 -0.742 0 2.0 1e-06 
0.0 -0.7419 0 2.0 1e-06 
0.0 -0.7418 0 2.0 1e-06 
0.0 -0.7417 0 2.0 1e-06 
0.0 -0.7416 0 2.0 1e-06 
0.0 -0.7415 0 2.0 1e-06 
0.0 -0.7414 0 2.0 1e-06 
0.0 -0.7413 0 2.0 1e-06 
0.0 -0.7412 0 2.0 1e-06 
0.0 -0.7411 0 2.0 1e-06 
0.0 -0.741 0 2.0 1e-06 
0.0 -0.7409 0 2.0 1e-06 
0.0 -0.7408 0 2.0 1e-06 
0.0 -0.7407 0 2.0 1e-06 
0.0 -0.7406 0 2.0 1e-06 
0.0 -0.7405 0 2.0 1e-06 
0.0 -0.7404 0 2.0 1e-06 
0.0 -0.7403 0 2.0 1e-06 
0.0 -0.7402 0 2.0 1e-06 
0.0 -0.7401 0 2.0 1e-06 
0.0 -0.74 0 2.0 1e-06 
0.0 -0.7399 0 2.0 1e-06 
0.0 -0.7398 0 2.0 1e-06 
0.0 -0.7397 0 2.0 1e-06 
0.0 -0.7396 0 2.0 1e-06 
0.0 -0.7395 0 2.0 1e-06 
0.0 -0.7394 0 2.0 1e-06 
0.0 -0.7393 0 2.0 1e-06 
0.0 -0.7392 0 2.0 1e-06 
0.0 -0.7391 0 2.0 1e-06 
0.0 -0.739 0 2.0 1e-06 
0.0 -0.7389 0 2.0 1e-06 
0.0 -0.7388 0 2.0 1e-06 
0.0 -0.7387 0 2.0 1e-06 
0.0 -0.7386 0 2.0 1e-06 
0.0 -0.7385 0 2.0 1e-06 
0.0 -0.7384 0 2.0 1e-06 
0.0 -0.7383 0 2.0 1e-06 
0.0 -0.7382 0 2.0 1e-06 
0.0 -0.7381 0 2.0 1e-06 
0.0 -0.738 0 2.0 1e-06 
0.0 -0.7379 0 2.0 1e-06 
0.0 -0.7378 0 2.0 1e-06 
0.0 -0.7377 0 2.0 1e-06 
0.0 -0.7376 0 2.0 1e-06 
0.0 -0.7375 0 2.0 1e-06 
0.0 -0.7374 0 2.0 1e-06 
0.0 -0.7373 0 2.0 1e-06 
0.0 -0.7372 0 2.0 1e-06 
0.0 -0.7371 0 2.0 1e-06 
0.0 -0.737 0 2.0 1e-06 
0.0 -0.7369 0 2.0 1e-06 
0.0 -0.7368 0 2.0 1e-06 
0.0 -0.7367 0 2.0 1e-06 
0.0 -0.7366 0 2.0 1e-06 
0.0 -0.7365 0 2.0 1e-06 
0.0 -0.7364 0 2.0 1e-06 
0.0 -0.7363 0 2.0 1e-06 
0.0 -0.7362 0 2.0 1e-06 
0.0 -0.7361 0 2.0 1e-06 
0.0 -0.736 0 2.0 1e-06 
0.0 -0.7359 0 2.0 1e-06 
0.0 -0.7358 0 2.0 1e-06 
0.0 -0.7357 0 2.0 1e-06 
0.0 -0.7356 0 2.0 1e-06 
0.0 -0.7355 0 2.0 1e-06 
0.0 -0.7354 0 2.0 1e-06 
0.0 -0.7353 0 2.0 1e-06 
0.0 -0.7352 0 2.0 1e-06 
0.0 -0.7351 0 2.0 1e-06 
0.0 -0.735 0 2.0 1e-06 
0.0 -0.7349 0 2.0 1e-06 
0.0 -0.7348 0 2.0 1e-06 
0.0 -0.7347 0 2.0 1e-06 
0.0 -0.7346 0 2.0 1e-06 
0.0 -0.7345 0 2.0 1e-06 
0.0 -0.7344 0 2.0 1e-06 
0.0 -0.7343 0 2.0 1e-06 
0.0 -0.7342 0 2.0 1e-06 
0.0 -0.7341 0 2.0 1e-06 
0.0 -0.734 0 2.0 1e-06 
0.0 -0.7339 0 2.0 1e-06 
0.0 -0.7338 0 2.0 1e-06 
0.0 -0.7337 0 2.0 1e-06 
0.0 -0.7336 0 2.0 1e-06 
0.0 -0.7335 0 2.0 1e-06 
0.0 -0.7334 0 2.0 1e-06 
0.0 -0.7333 0 2.0 1e-06 
0.0 -0.7332 0 2.0 1e-06 
0.0 -0.7331 0 2.0 1e-06 
0.0 -0.733 0 2.0 1e-06 
0.0 -0.7329 0 2.0 1e-06 
0.0 -0.7328 0 2.0 1e-06 
0.0 -0.7327 0 2.0 1e-06 
0.0 -0.7326 0 2.0 1e-06 
0.0 -0.7325 0 2.0 1e-06 
0.0 -0.7324 0 2.0 1e-06 
0.0 -0.7323 0 2.0 1e-06 
0.0 -0.7322 0 2.0 1e-06 
0.0 -0.7321 0 2.0 1e-06 
0.0 -0.732 0 2.0 1e-06 
0.0 -0.7319 0 2.0 1e-06 
0.0 -0.7318 0 2.0 1e-06 
0.0 -0.7317 0 2.0 1e-06 
0.0 -0.7316 0 2.0 1e-06 
0.0 -0.7315 0 2.0 1e-06 
0.0 -0.7314 0 2.0 1e-06 
0.0 -0.7313 0 2.0 1e-06 
0.0 -0.7312 0 2.0 1e-06 
0.0 -0.7311 0 2.0 1e-06 
0.0 -0.731 0 2.0 1e-06 
0.0 -0.7309 0 2.0 1e-06 
0.0 -0.7308 0 2.0 1e-06 
0.0 -0.7307 0 2.0 1e-06 
0.0 -0.7306 0 2.0 1e-06 
0.0 -0.7305 0 2.0 1e-06 
0.0 -0.7304 0 2.0 1e-06 
0.0 -0.7303 0 2.0 1e-06 
0.0 -0.7302 0 2.0 1e-06 
0.0 -0.7301 0 2.0 1e-06 
0.0 -0.73 0 2.0 1e-06 
0.0 -0.7299 0 2.0 1e-06 
0.0 -0.7298 0 2.0 1e-06 
0.0 -0.7297 0 2.0 1e-06 
0.0 -0.7296 0 2.0 1e-06 
0.0 -0.7295 0 2.0 1e-06 
0.0 -0.7294 0 2.0 1e-06 
0.0 -0.7293 0 2.0 1e-06 
0.0 -0.7292 0 2.0 1e-06 
0.0 -0.7291 0 2.0 1e-06 
0.0 -0.729 0 2.0 1e-06 
0.0 -0.7289 0 2.0 1e-06 
0.0 -0.7288 0 2.0 1e-06 
0.0 -0.7287 0 2.0 1e-06 
0.0 -0.7286 0 2.0 1e-06 
0.0 -0.7285 0 2.0 1e-06 
0.0 -0.7284 0 2.0 1e-06 
0.0 -0.7283 0 2.0 1e-06 
0.0 -0.7282 0 2.0 1e-06 
0.0 -0.7281 0 2.0 1e-06 
0.0 -0.728 0 2.0 1e-06 
0.0 -0.7279 0 2.0 1e-06 
0.0 -0.7278 0 2.0 1e-06 
0.0 -0.7277 0 2.0 1e-06 
0.0 -0.7276 0 2.0 1e-06 
0.0 -0.7275 0 2.0 1e-06 
0.0 -0.7274 0 2.0 1e-06 
0.0 -0.7273 0 2.0 1e-06 
0.0 -0.7272 0 2.0 1e-06 
0.0 -0.7271 0 2.0 1e-06 
0.0 -0.727 0 2.0 1e-06 
0.0 -0.7269 0 2.0 1e-06 
0.0 -0.7268 0 2.0 1e-06 
0.0 -0.7267 0 2.0 1e-06 
0.0 -0.7266 0 2.0 1e-06 
0.0 -0.7265 0 2.0 1e-06 
0.0 -0.7264 0 2.0 1e-06 
0.0 -0.7263 0 2.0 1e-06 
0.0 -0.7262 0 2.0 1e-06 
0.0 -0.7261 0 2.0 1e-06 
0.0 -0.726 0 2.0 1e-06 
0.0 -0.7259 0 2.0 1e-06 
0.0 -0.7258 0 2.0 1e-06 
0.0 -0.7257 0 2.0 1e-06 
0.0 -0.7256 0 2.0 1e-06 
0.0 -0.7255 0 2.0 1e-06 
0.0 -0.7254 0 2.0 1e-06 
0.0 -0.7253 0 2.0 1e-06 
0.0 -0.7252 0 2.0 1e-06 
0.0 -0.7251 0 2.0 1e-06 
0.0 -0.725 0 2.0 1e-06 
0.0 -0.7249 0 2.0 1e-06 
0.0 -0.7248 0 2.0 1e-06 
0.0 -0.7247 0 2.0 1e-06 
0.0 -0.7246 0 2.0 1e-06 
0.0 -0.7245 0 2.0 1e-06 
0.0 -0.7244 0 2.0 1e-06 
0.0 -0.7243 0 2.0 1e-06 
0.0 -0.7242 0 2.0 1e-06 
0.0 -0.7241 0 2.0 1e-06 
0.0 -0.724 0 2.0 1e-06 
0.0 -0.7239 0 2.0 1e-06 
0.0 -0.7238 0 2.0 1e-06 
0.0 -0.7237 0 2.0 1e-06 
0.0 -0.7236 0 2.0 1e-06 
0.0 -0.7235 0 2.0 1e-06 
0.0 -0.7234 0 2.0 1e-06 
0.0 -0.7233 0 2.0 1e-06 
0.0 -0.7232 0 2.0 1e-06 
0.0 -0.7231 0 2.0 1e-06 
0.0 -0.723 0 2.0 1e-06 
0.0 -0.7229 0 2.0 1e-06 
0.0 -0.7228 0 2.0 1e-06 
0.0 -0.7227 0 2.0 1e-06 
0.0 -0.7226 0 2.0 1e-06 
0.0 -0.7225 0 2.0 1e-06 
0.0 -0.7224 0 2.0 1e-06 
0.0 -0.7223 0 2.0 1e-06 
0.0 -0.7222 0 2.0 1e-06 
0.0 -0.7221 0 2.0 1e-06 
0.0 -0.722 0 2.0 1e-06 
0.0 -0.7219 0 2.0 1e-06 
0.0 -0.7218 0 2.0 1e-06 
0.0 -0.7217 0 2.0 1e-06 
0.0 -0.7216 0 2.0 1e-06 
0.0 -0.7215 0 2.0 1e-06 
0.0 -0.7214 0 2.0 1e-06 
0.0 -0.7213 0 2.0 1e-06 
0.0 -0.7212 0 2.0 1e-06 
0.0 -0.7211 0 2.0 1e-06 
0.0 -0.721 0 2.0 1e-06 
0.0 -0.7209 0 2.0 1e-06 
0.0 -0.7208 0 2.0 1e-06 
0.0 -0.7207 0 2.0 1e-06 
0.0 -0.7206 0 2.0 1e-06 
0.0 -0.7205 0 2.0 1e-06 
0.0 -0.7204 0 2.0 1e-06 
0.0 -0.7203 0 2.0 1e-06 
0.0 -0.7202 0 2.0 1e-06 
0.0 -0.7201 0 2.0 1e-06 
0.0 -0.72 0 2.0 1e-06 
0.0 -0.7199 0 2.0 1e-06 
0.0 -0.7198 0 2.0 1e-06 
0.0 -0.7197 0 2.0 1e-06 
0.0 -0.7196 0 2.0 1e-06 
0.0 -0.7195 0 2.0 1e-06 
0.0 -0.7194 0 2.0 1e-06 
0.0 -0.7193 0 2.0 1e-06 
0.0 -0.7192 0 2.0 1e-06 
0.0 -0.7191 0 2.0 1e-06 
0.0 -0.719 0 2.0 1e-06 
0.0 -0.7189 0 2.0 1e-06 
0.0 -0.7188 0 2.0 1e-06 
0.0 -0.7187 0 2.0 1e-06 
0.0 -0.7186 0 2.0 1e-06 
0.0 -0.7185 0 2.0 1e-06 
0.0 -0.7184 0 2.0 1e-06 
0.0 -0.7183 0 2.0 1e-06 
0.0 -0.7182 0 2.0 1e-06 
0.0 -0.7181 0 2.0 1e-06 
0.0 -0.718 0 2.0 1e-06 
0.0 -0.7179 0 2.0 1e-06 
0.0 -0.7178 0 2.0 1e-06 
0.0 -0.7177 0 2.0 1e-06 
0.0 -0.7176 0 2.0 1e-06 
0.0 -0.7175 0 2.0 1e-06 
0.0 -0.7174 0 2.0 1e-06 
0.0 -0.7173 0 2.0 1e-06 
0.0 -0.7172 0 2.0 1e-06 
0.0 -0.7171 0 2.0 1e-06 
0.0 -0.717 0 2.0 1e-06 
0.0 -0.7169 0 2.0 1e-06 
0.0 -0.7168 0 2.0 1e-06 
0.0 -0.7167 0 2.0 1e-06 
0.0 -0.7166 0 2.0 1e-06 
0.0 -0.7165 0 2.0 1e-06 
0.0 -0.7164 0 2.0 1e-06 
0.0 -0.7163 0 2.0 1e-06 
0.0 -0.7162 0 2.0 1e-06 
0.0 -0.7161 0 2.0 1e-06 
0.0 -0.716 0 2.0 1e-06 
0.0 -0.7159 0 2.0 1e-06 
0.0 -0.7158 0 2.0 1e-06 
0.0 -0.7157 0 2.0 1e-06 
0.0 -0.7156 0 2.0 1e-06 
0.0 -0.7155 0 2.0 1e-06 
0.0 -0.7154 0 2.0 1e-06 
0.0 -0.7153 0 2.0 1e-06 
0.0 -0.7152 0 2.0 1e-06 
0.0 -0.7151 0 2.0 1e-06 
0.0 -0.715 0 2.0 1e-06 
0.0 -0.7149 0 2.0 1e-06 
0.0 -0.7148 0 2.0 1e-06 
0.0 -0.7147 0 2.0 1e-06 
0.0 -0.7146 0 2.0 1e-06 
0.0 -0.7145 0 2.0 1e-06 
0.0 -0.7144 0 2.0 1e-06 
0.0 -0.7143 0 2.0 1e-06 
0.0 -0.7142 0 2.0 1e-06 
0.0 -0.7141 0 2.0 1e-06 
0.0 -0.714 0 2.0 1e-06 
0.0 -0.7139 0 2.0 1e-06 
0.0 -0.7138 0 2.0 1e-06 
0.0 -0.7137 0 2.0 1e-06 
0.0 -0.7136 0 2.0 1e-06 
0.0 -0.7135 0 2.0 1e-06 
0.0 -0.7134 0 2.0 1e-06 
0.0 -0.7133 0 2.0 1e-06 
0.0 -0.7132 0 2.0 1e-06 
0.0 -0.7131 0 2.0 1e-06 
0.0 -0.713 0 2.0 1e-06 
0.0 -0.7129 0 2.0 1e-06 
0.0 -0.7128 0 2.0 1e-06 
0.0 -0.7127 0 2.0 1e-06 
0.0 -0.7126 0 2.0 1e-06 
0.0 -0.7125 0 2.0 1e-06 
0.0 -0.7124 0 2.0 1e-06 
0.0 -0.7123 0 2.0 1e-06 
0.0 -0.7122 0 2.0 1e-06 
0.0 -0.7121 0 2.0 1e-06 
0.0 -0.712 0 2.0 1e-06 
0.0 -0.7119 0 2.0 1e-06 
0.0 -0.7118 0 2.0 1e-06 
0.0 -0.7117 0 2.0 1e-06 
0.0 -0.7116 0 2.0 1e-06 
0.0 -0.7115 0 2.0 1e-06 
0.0 -0.7114 0 2.0 1e-06 
0.0 -0.7113 0 2.0 1e-06 
0.0 -0.7112 0 2.0 1e-06 
0.0 -0.7111 0 2.0 1e-06 
0.0 -0.711 0 2.0 1e-06 
0.0 -0.7109 0 2.0 1e-06 
0.0 -0.7108 0 2.0 1e-06 
0.0 -0.7107 0 2.0 1e-06 
0.0 -0.7106 0 2.0 1e-06 
0.0 -0.7105 0 2.0 1e-06 
0.0 -0.7104 0 2.0 1e-06 
0.0 -0.7103 0 2.0 1e-06 
0.0 -0.7102 0 2.0 1e-06 
0.0 -0.7101 0 2.0 1e-06 
0.0 -0.71 0 2.0 1e-06 
0.0 -0.7099 0 2.0 1e-06 
0.0 -0.7098 0 2.0 1e-06 
0.0 -0.7097 0 2.0 1e-06 
0.0 -0.7096 0 2.0 1e-06 
0.0 -0.7095 0 2.0 1e-06 
0.0 -0.7094 0 2.0 1e-06 
0.0 -0.7093 0 2.0 1e-06 
0.0 -0.7092 0 2.0 1e-06 
0.0 -0.7091 0 2.0 1e-06 
0.0 -0.709 0 2.0 1e-06 
0.0 -0.7089 0 2.0 1e-06 
0.0 -0.7088 0 2.0 1e-06 
0.0 -0.7087 0 2.0 1e-06 
0.0 -0.7086 0 2.0 1e-06 
0.0 -0.7085 0 2.0 1e-06 
0.0 -0.7084 0 2.0 1e-06 
0.0 -0.7083 0 2.0 1e-06 
0.0 -0.7082 0 2.0 1e-06 
0.0 -0.7081 0 2.0 1e-06 
0.0 -0.708 0 2.0 1e-06 
0.0 -0.7079 0 2.0 1e-06 
0.0 -0.7078 0 2.0 1e-06 
0.0 -0.7077 0 2.0 1e-06 
0.0 -0.7076 0 2.0 1e-06 
0.0 -0.7075 0 2.0 1e-06 
0.0 -0.7074 0 2.0 1e-06 
0.0 -0.7073 0 2.0 1e-06 
0.0 -0.7072 0 2.0 1e-06 
0.0 -0.7071 0 2.0 1e-06 
0.0 -0.707 0 2.0 1e-06 
0.0 -0.7069 0 2.0 1e-06 
0.0 -0.7068 0 2.0 1e-06 
0.0 -0.7067 0 2.0 1e-06 
0.0 -0.7066 0 2.0 1e-06 
0.0 -0.7065 0 2.0 1e-06 
0.0 -0.7064 0 2.0 1e-06 
0.0 -0.7063 0 2.0 1e-06 
0.0 -0.7062 0 2.0 1e-06 
0.0 -0.7061 0 2.0 1e-06 
0.0 -0.706 0 2.0 1e-06 
0.0 -0.7059 0 2.0 1e-06 
0.0 -0.7058 0 2.0 1e-06 
0.0 -0.7057 0 2.0 1e-06 
0.0 -0.7056 0 2.0 1e-06 
0.0 -0.7055 0 2.0 1e-06 
0.0 -0.7054 0 2.0 1e-06 
0.0 -0.7053 0 2.0 1e-06 
0.0 -0.7052 0 2.0 1e-06 
0.0 -0.7051 0 2.0 1e-06 
0.0 -0.705 0 2.0 1e-06 
0.0 -0.7049 0 2.0 1e-06 
0.0 -0.7048 0 2.0 1e-06 
0.0 -0.7047 0 2.0 1e-06 
0.0 -0.7046 0 2.0 1e-06 
0.0 -0.7045 0 2.0 1e-06 
0.0 -0.7044 0 2.0 1e-06 
0.0 -0.7043 0 2.0 1e-06 
0.0 -0.7042 0 2.0 1e-06 
0.0 -0.7041 0 2.0 1e-06 
0.0 -0.704 0 2.0 1e-06 
0.0 -0.7039 0 2.0 1e-06 
0.0 -0.7038 0 2.0 1e-06 
0.0 -0.7037 0 2.0 1e-06 
0.0 -0.7036 0 2.0 1e-06 
0.0 -0.7035 0 2.0 1e-06 
0.0 -0.7034 0 2.0 1e-06 
0.0 -0.7033 0 2.0 1e-06 
0.0 -0.7032 0 2.0 1e-06 
0.0 -0.7031 0 2.0 1e-06 
0.0 -0.703 0 2.0 1e-06 
0.0 -0.7029 0 2.0 1e-06 
0.0 -0.7028 0 2.0 1e-06 
0.0 -0.7027 0 2.0 1e-06 
0.0 -0.7026 0 2.0 1e-06 
0.0 -0.7025 0 2.0 1e-06 
0.0 -0.7024 0 2.0 1e-06 
0.0 -0.7023 0 2.0 1e-06 
0.0 -0.7022 0 2.0 1e-06 
0.0 -0.7021 0 2.0 1e-06 
0.0 -0.702 0 2.0 1e-06 
0.0 -0.7019 0 2.0 1e-06 
0.0 -0.7018 0 2.0 1e-06 
0.0 -0.7017 0 2.0 1e-06 
0.0 -0.7016 0 2.0 1e-06 
0.0 -0.7015 0 2.0 1e-06 
0.0 -0.7014 0 2.0 1e-06 
0.0 -0.7013 0 2.0 1e-06 
0.0 -0.7012 0 2.0 1e-06 
0.0 -0.7011 0 2.0 1e-06 
0.0 -0.701 0 2.0 1e-06 
0.0 -0.7009 0 2.0 1e-06 
0.0 -0.7008 0 2.0 1e-06 
0.0 -0.7007 0 2.0 1e-06 
0.0 -0.7006 0 2.0 1e-06 
0.0 -0.7005 0 2.0 1e-06 
0.0 -0.7004 0 2.0 1e-06 
0.0 -0.7003 0 2.0 1e-06 
0.0 -0.7002 0 2.0 1e-06 
0.0 -0.7001 0 2.0 1e-06 
0.0 -0.7 0 2.0 1e-06 
0.0 -0.6999 0 2.0 1e-06 
0.0 -0.6998 0 2.0 1e-06 
0.0 -0.6997 0 2.0 1e-06 
0.0 -0.6996 0 2.0 1e-06 
0.0 -0.6995 0 2.0 1e-06 
0.0 -0.6994 0 2.0 1e-06 
0.0 -0.6993 0 2.0 1e-06 
0.0 -0.6992 0 2.0 1e-06 
0.0 -0.6991 0 2.0 1e-06 
0.0 -0.699 0 2.0 1e-06 
0.0 -0.6989 0 2.0 1e-06 
0.0 -0.6988 0 2.0 1e-06 
0.0 -0.6987 0 2.0 1e-06 
0.0 -0.6986 0 2.0 1e-06 
0.0 -0.6985 0 2.0 1e-06 
0.0 -0.6984 0 2.0 1e-06 
0.0 -0.6983 0 2.0 1e-06 
0.0 -0.6982 0 2.0 1e-06 
0.0 -0.6981 0 2.0 1e-06 
0.0 -0.698 0 2.0 1e-06 
0.0 -0.6979 0 2.0 1e-06 
0.0 -0.6978 0 2.0 1e-06 
0.0 -0.6977 0 2.0 1e-06 
0.0 -0.6976 0 2.0 1e-06 
0.0 -0.6975 0 2.0 1e-06 
0.0 -0.6974 0 2.0 1e-06 
0.0 -0.6973 0 2.0 1e-06 
0.0 -0.6972 0 2.0 1e-06 
0.0 -0.6971 0 2.0 1e-06 
0.0 -0.697 0 2.0 1e-06 
0.0 -0.6969 0 2.0 1e-06 
0.0 -0.6968 0 2.0 1e-06 
0.0 -0.6967 0 2.0 1e-06 
0.0 -0.6966 0 2.0 1e-06 
0.0 -0.6965 0 2.0 1e-06 
0.0 -0.6964 0 2.0 1e-06 
0.0 -0.6963 0 2.0 1e-06 
0.0 -0.6962 0 2.0 1e-06 
0.0 -0.6961 0 2.0 1e-06 
0.0 -0.696 0 2.0 1e-06 
0.0 -0.6959 0 2.0 1e-06 
0.0 -0.6958 0 2.0 1e-06 
0.0 -0.6957 0 2.0 1e-06 
0.0 -0.6956 0 2.0 1e-06 
0.0 -0.6955 0 2.0 1e-06 
0.0 -0.6954 0 2.0 1e-06 
0.0 -0.6953 0 2.0 1e-06 
0.0 -0.6952 0 2.0 1e-06 
0.0 -0.6951 0 2.0 1e-06 
0.0 -0.695 0 2.0 1e-06 
0.0 -0.6949 0 2.0 1e-06 
0.0 -0.6948 0 2.0 1e-06 
0.0 -0.6947 0 2.0 1e-06 
0.0 -0.6946 0 2.0 1e-06 
0.0 -0.6945 0 2.0 1e-06 
0.0 -0.6944 0 2.0 1e-06 
0.0 -0.6943 0 2.0 1e-06 
0.0 -0.6942 0 2.0 1e-06 
0.0 -0.6941 0 2.0 1e-06 
0.0 -0.694 0 2.0 1e-06 
0.0 -0.6939 0 2.0 1e-06 
0.0 -0.6938 0 2.0 1e-06 
0.0 -0.6937 0 2.0 1e-06 
0.0 -0.6936 0 2.0 1e-06 
0.0 -0.6935 0 2.0 1e-06 
0.0 -0.6934 0 2.0 1e-06 
0.0 -0.6933 0 2.0 1e-06 
0.0 -0.6932 0 2.0 1e-06 
0.0 -0.6931 0 2.0 1e-06 
0.0 -0.693 0 2.0 1e-06 
0.0 -0.6929 0 2.0 1e-06 
0.0 -0.6928 0 2.0 1e-06 
0.0 -0.6927 0 2.0 1e-06 
0.0 -0.6926 0 2.0 1e-06 
0.0 -0.6925 0 2.0 1e-06 
0.0 -0.6924 0 2.0 1e-06 
0.0 -0.6923 0 2.0 1e-06 
0.0 -0.6922 0 2.0 1e-06 
0.0 -0.6921 0 2.0 1e-06 
0.0 -0.692 0 2.0 1e-06 
0.0 -0.6919 0 2.0 1e-06 
0.0 -0.6918 0 2.0 1e-06 
0.0 -0.6917 0 2.0 1e-06 
0.0 -0.6916 0 2.0 1e-06 
0.0 -0.6915 0 2.0 1e-06 
0.0 -0.6914 0 2.0 1e-06 
0.0 -0.6913 0 2.0 1e-06 
0.0 -0.6912 0 2.0 1e-06 
0.0 -0.6911 0 2.0 1e-06 
0.0 -0.691 0 2.0 1e-06 
0.0 -0.6909 0 2.0 1e-06 
0.0 -0.6908 0 2.0 1e-06 
0.0 -0.6907 0 2.0 1e-06 
0.0 -0.6906 0 2.0 1e-06 
0.0 -0.6905 0 2.0 1e-06 
0.0 -0.6904 0 2.0 1e-06 
0.0 -0.6903 0 2.0 1e-06 
0.0 -0.6902 0 2.0 1e-06 
0.0 -0.6901 0 2.0 1e-06 
0.0 -0.69 0 2.0 1e-06 
0.0 -0.6899 0 2.0 1e-06 
0.0 -0.6898 0 2.0 1e-06 
0.0 -0.6897 0 2.0 1e-06 
0.0 -0.6896 0 2.0 1e-06 
0.0 -0.6895 0 2.0 1e-06 
0.0 -0.6894 0 2.0 1e-06 
0.0 -0.6893 0 2.0 1e-06 
0.0 -0.6892 0 2.0 1e-06 
0.0 -0.6891 0 2.0 1e-06 
0.0 -0.689 0 2.0 1e-06 
0.0 -0.6889 0 2.0 1e-06 
0.0 -0.6888 0 2.0 1e-06 
0.0 -0.6887 0 2.0 1e-06 
0.0 -0.6886 0 2.0 1e-06 
0.0 -0.6885 0 2.0 1e-06 
0.0 -0.6884 0 2.0 1e-06 
0.0 -0.6883 0 2.0 1e-06 
0.0 -0.6882 0 2.0 1e-06 
0.0 -0.6881 0 2.0 1e-06 
0.0 -0.688 0 2.0 1e-06 
0.0 -0.6879 0 2.0 1e-06 
0.0 -0.6878 0 2.0 1e-06 
0.0 -0.6877 0 2.0 1e-06 
0.0 -0.6876 0 2.0 1e-06 
0.0 -0.6875 0 2.0 1e-06 
0.0 -0.6874 0 2.0 1e-06 
0.0 -0.6873 0 2.0 1e-06 
0.0 -0.6872 0 2.0 1e-06 
0.0 -0.6871 0 2.0 1e-06 
0.0 -0.687 0 2.0 1e-06 
0.0 -0.6869 0 2.0 1e-06 
0.0 -0.6868 0 2.0 1e-06 
0.0 -0.6867 0 2.0 1e-06 
0.0 -0.6866 0 2.0 1e-06 
0.0 -0.6865 0 2.0 1e-06 
0.0 -0.6864 0 2.0 1e-06 
0.0 -0.6863 0 2.0 1e-06 
0.0 -0.6862 0 2.0 1e-06 
0.0 -0.6861 0 2.0 1e-06 
0.0 -0.686 0 2.0 1e-06 
0.0 -0.6859 0 2.0 1e-06 
0.0 -0.6858 0 2.0 1e-06 
0.0 -0.6857 0 2.0 1e-06 
0.0 -0.6856 0 2.0 1e-06 
0.0 -0.6855 0 2.0 1e-06 
0.0 -0.6854 0 2.0 1e-06 
0.0 -0.6853 0 2.0 1e-06 
0.0 -0.6852 0 2.0 1e-06 
0.0 -0.6851 0 2.0 1e-06 
0.0 -0.685 0 2.0 1e-06 
0.0 -0.6849 0 2.0 1e-06 
0.0 -0.6848 0 2.0 1e-06 
0.0 -0.6847 0 2.0 1e-06 
0.0 -0.6846 0 2.0 1e-06 
0.0 -0.6845 0 2.0 1e-06 
0.0 -0.6844 0 2.0 1e-06 
0.0 -0.6843 0 2.0 1e-06 
0.0 -0.6842 0 2.0 1e-06 
0.0 -0.6841 0 2.0 1e-06 
0.0 -0.684 0 2.0 1e-06 
0.0 -0.6839 0 2.0 1e-06 
0.0 -0.6838 0 2.0 1e-06 
0.0 -0.6837 0 2.0 1e-06 
0.0 -0.6836 0 2.0 1e-06 
0.0 -0.6835 0 2.0 1e-06 
0.0 -0.6834 0 2.0 1e-06 
0.0 -0.6833 0 2.0 1e-06 
0.0 -0.6832 0 2.0 1e-06 
0.0 -0.6831 0 2.0 1e-06 
0.0 -0.683 0 2.0 1e-06 
0.0 -0.6829 0 2.0 1e-06 
0.0 -0.6828 0 2.0 1e-06 
0.0 -0.6827 0 2.0 1e-06 
0.0 -0.6826 0 2.0 1e-06 
0.0 -0.6825 0 2.0 1e-06 
0.0 -0.6824 0 2.0 1e-06 
0.0 -0.6823 0 2.0 1e-06 
0.0 -0.6822 0 2.0 1e-06 
0.0 -0.6821 0 2.0 1e-06 
0.0 -0.682 0 2.0 1e-06 
0.0 -0.6819 0 2.0 1e-06 
0.0 -0.6818 0 2.0 1e-06 
0.0 -0.6817 0 2.0 1e-06 
0.0 -0.6816 0 2.0 1e-06 
0.0 -0.6815 0 2.0 1e-06 
0.0 -0.6814 0 2.0 1e-06 
0.0 -0.6813 0 2.0 1e-06 
0.0 -0.6812 0 2.0 1e-06 
0.0 -0.6811 0 2.0 1e-06 
0.0 -0.681 0 2.0 1e-06 
0.0 -0.6809 0 2.0 1e-06 
0.0 -0.6808 0 2.0 1e-06 
0.0 -0.6807 0 2.0 1e-06 
0.0 -0.6806 0 2.0 1e-06 
0.0 -0.6805 0 2.0 1e-06 
0.0 -0.6804 0 2.0 1e-06 
0.0 -0.6803 0 2.0 1e-06 
0.0 -0.6802 0 2.0 1e-06 
0.0 -0.6801 0 2.0 1e-06 
0.0 -0.68 0 2.0 1e-06 
0.0 -0.6799 0 2.0 1e-06 
0.0 -0.6798 0 2.0 1e-06 
0.0 -0.6797 0 2.0 1e-06 
0.0 -0.6796 0 2.0 1e-06 
0.0 -0.6795 0 2.0 1e-06 
0.0 -0.6794 0 2.0 1e-06 
0.0 -0.6793 0 2.0 1e-06 
0.0 -0.6792 0 2.0 1e-06 
0.0 -0.6791 0 2.0 1e-06 
0.0 -0.679 0 2.0 1e-06 
0.0 -0.6789 0 2.0 1e-06 
0.0 -0.6788 0 2.0 1e-06 
0.0 -0.6787 0 2.0 1e-06 
0.0 -0.6786 0 2.0 1e-06 
0.0 -0.6785 0 2.0 1e-06 
0.0 -0.6784 0 2.0 1e-06 
0.0 -0.6783 0 2.0 1e-06 
0.0 -0.6782 0 2.0 1e-06 
0.0 -0.6781 0 2.0 1e-06 
0.0 -0.678 0 2.0 1e-06 
0.0 -0.6779 0 2.0 1e-06 
0.0 -0.6778 0 2.0 1e-06 
0.0 -0.6777 0 2.0 1e-06 
0.0 -0.6776 0 2.0 1e-06 
0.0 -0.6775 0 2.0 1e-06 
0.0 -0.6774 0 2.0 1e-06 
0.0 -0.6773 0 2.0 1e-06 
0.0 -0.6772 0 2.0 1e-06 
0.0 -0.6771 0 2.0 1e-06 
0.0 -0.677 0 2.0 1e-06 
0.0 -0.6769 0 2.0 1e-06 
0.0 -0.6768 0 2.0 1e-06 
0.0 -0.6767 0 2.0 1e-06 
0.0 -0.6766 0 2.0 1e-06 
0.0 -0.6765 0 2.0 1e-06 
0.0 -0.6764 0 2.0 1e-06 
0.0 -0.6763 0 2.0 1e-06 
0.0 -0.6762 0 2.0 1e-06 
0.0 -0.6761 0 2.0 1e-06 
0.0 -0.676 0 2.0 1e-06 
0.0 -0.6759 0 2.0 1e-06 
0.0 -0.6758 0 2.0 1e-06 
0.0 -0.6757 0 2.0 1e-06 
0.0 -0.6756 0 2.0 1e-06 
0.0 -0.6755 0 2.0 1e-06 
0.0 -0.6754 0 2.0 1e-06 
0.0 -0.6753 0 2.0 1e-06 
0.0 -0.6752 0 2.0 1e-06 
0.0 -0.6751 0 2.0 1e-06 
0.0 -0.675 0 2.0 1e-06 
0.0 -0.6749 0 2.0 1e-06 
0.0 -0.6748 0 2.0 1e-06 
0.0 -0.6747 0 2.0 1e-06 
0.0 -0.6746 0 2.0 1e-06 
0.0 -0.6745 0 2.0 1e-06 
0.0 -0.6744 0 2.0 1e-06 
0.0 -0.6743 0 2.0 1e-06 
0.0 -0.6742 0 2.0 1e-06 
0.0 -0.6741 0 2.0 1e-06 
0.0 -0.674 0 2.0 1e-06 
0.0 -0.6739 0 2.0 1e-06 
0.0 -0.6738 0 2.0 1e-06 
0.0 -0.6737 0 2.0 1e-06 
0.0 -0.6736 0 2.0 1e-06 
0.0 -0.6735 0 2.0 1e-06 
0.0 -0.6734 0 2.0 1e-06 
0.0 -0.6733 0 2.0 1e-06 
0.0 -0.6732 0 2.0 1e-06 
0.0 -0.6731 0 2.0 1e-06 
0.0 -0.673 0 2.0 1e-06 
0.0 -0.6729 0 2.0 1e-06 
0.0 -0.6728 0 2.0 1e-06 
0.0 -0.6727 0 2.0 1e-06 
0.0 -0.6726 0 2.0 1e-06 
0.0 -0.6725 0 2.0 1e-06 
0.0 -0.6724 0 2.0 1e-06 
0.0 -0.6723 0 2.0 1e-06 
0.0 -0.6722 0 2.0 1e-06 
0.0 -0.6721 0 2.0 1e-06 
0.0 -0.672 0 2.0 1e-06 
0.0 -0.6719 0 2.0 1e-06 
0.0 -0.6718 0 2.0 1e-06 
0.0 -0.6717 0 2.0 1e-06 
0.0 -0.6716 0 2.0 1e-06 
0.0 -0.6715 0 2.0 1e-06 
0.0 -0.6714 0 2.0 1e-06 
0.0 -0.6713 0 2.0 1e-06 
0.0 -0.6712 0 2.0 1e-06 
0.0 -0.6711 0 2.0 1e-06 
0.0 -0.671 0 2.0 1e-06 
0.0 -0.6709 0 2.0 1e-06 
0.0 -0.6708 0 2.0 1e-06 
0.0 -0.6707 0 2.0 1e-06 
0.0 -0.6706 0 2.0 1e-06 
0.0 -0.6705 0 2.0 1e-06 
0.0 -0.6704 0 2.0 1e-06 
0.0 -0.6703 0 2.0 1e-06 
0.0 -0.6702 0 2.0 1e-06 
0.0 -0.6701 0 2.0 1e-06 
0.0 -0.67 0 2.0 1e-06 
0.0 -0.6699 0 2.0 1e-06 
0.0 -0.6698 0 2.0 1e-06 
0.0 -0.6697 0 2.0 1e-06 
0.0 -0.6696 0 2.0 1e-06 
0.0 -0.6695 0 2.0 1e-06 
0.0 -0.6694 0 2.0 1e-06 
0.0 -0.6693 0 2.0 1e-06 
0.0 -0.6692 0 2.0 1e-06 
0.0 -0.6691 0 2.0 1e-06 
0.0 -0.669 0 2.0 1e-06 
0.0 -0.6689 0 2.0 1e-06 
0.0 -0.6688 0 2.0 1e-06 
0.0 -0.6687 0 2.0 1e-06 
0.0 -0.6686 0 2.0 1e-06 
0.0 -0.6685 0 2.0 1e-06 
0.0 -0.6684 0 2.0 1e-06 
0.0 -0.6683 0 2.0 1e-06 
0.0 -0.6682 0 2.0 1e-06 
0.0 -0.6681 0 2.0 1e-06 
0.0 -0.668 0 2.0 1e-06 
0.0 -0.6679 0 2.0 1e-06 
0.0 -0.6678 0 2.0 1e-06 
0.0 -0.6677 0 2.0 1e-06 
0.0 -0.6676 0 2.0 1e-06 
0.0 -0.6675 0 2.0 1e-06 
0.0 -0.6674 0 2.0 1e-06 
0.0 -0.6673 0 2.0 1e-06 
0.0 -0.6672 0 2.0 1e-06 
0.0 -0.6671 0 2.0 1e-06 
0.0 -0.667 0 2.0 1e-06 
0.0 -0.6669 0 2.0 1e-06 
0.0 -0.6668 0 2.0 1e-06 
0.0 -0.6667 0 2.0 1e-06 
0.0 -0.6666 0 2.0 1e-06 
0.0 -0.6665 0 2.0 1e-06 
0.0 -0.6664 0 2.0 1e-06 
0.0 -0.6663 0 2.0 1e-06 
0.0 -0.6662 0 2.0 1e-06 
0.0 -0.6661 0 2.0 1e-06 
0.0 -0.666 0 2.0 1e-06 
0.0 -0.6659 0 2.0 1e-06 
0.0 -0.6658 0 2.0 1e-06 
0.0 -0.6657 0 2.0 1e-06 
0.0 -0.6656 0 2.0 1e-06 
0.0 -0.6655 0 2.0 1e-06 
0.0 -0.6654 0 2.0 1e-06 
0.0 -0.6653 0 2.0 1e-06 
0.0 -0.6652 0 2.0 1e-06 
0.0 -0.6651 0 2.0 1e-06 
0.0 -0.665 0 2.0 1e-06 
0.0 -0.6649 0 2.0 1e-06 
0.0 -0.6648 0 2.0 1e-06 
0.0 -0.6647 0 2.0 1e-06 
0.0 -0.6646 0 2.0 1e-06 
0.0 -0.6645 0 2.0 1e-06 
0.0 -0.6644 0 2.0 1e-06 
0.0 -0.6643 0 2.0 1e-06 
0.0 -0.6642 0 2.0 1e-06 
0.0 -0.6641 0 2.0 1e-06 
0.0 -0.664 0 2.0 1e-06 
0.0 -0.6639 0 2.0 1e-06 
0.0 -0.6638 0 2.0 1e-06 
0.0 -0.6637 0 2.0 1e-06 
0.0 -0.6636 0 2.0 1e-06 
0.0 -0.6635 0 2.0 1e-06 
0.0 -0.6634 0 2.0 1e-06 
0.0 -0.6633 0 2.0 1e-06 
0.0 -0.6632 0 2.0 1e-06 
0.0 -0.6631 0 2.0 1e-06 
0.0 -0.663 0 2.0 1e-06 
0.0 -0.6629 0 2.0 1e-06 
0.0 -0.6628 0 2.0 1e-06 
0.0 -0.6627 0 2.0 1e-06 
0.0 -0.6626 0 2.0 1e-06 
0.0 -0.6625 0 2.0 1e-06 
0.0 -0.6624 0 2.0 1e-06 
0.0 -0.6623 0 2.0 1e-06 
0.0 -0.6622 0 2.0 1e-06 
0.0 -0.6621 0 2.0 1e-06 
0.0 -0.662 0 2.0 1e-06 
0.0 -0.6619 0 2.0 1e-06 
0.0 -0.6618 0 2.0 1e-06 
0.0 -0.6617 0 2.0 1e-06 
0.0 -0.6616 0 2.0 1e-06 
0.0 -0.6615 0 2.0 1e-06 
0.0 -0.6614 0 2.0 1e-06 
0.0 -0.6613 0 2.0 1e-06 
0.0 -0.6612 0 2.0 1e-06 
0.0 -0.6611 0 2.0 1e-06 
0.0 -0.661 0 2.0 1e-06 
0.0 -0.6609 0 2.0 1e-06 
0.0 -0.6608 0 2.0 1e-06 
0.0 -0.6607 0 2.0 1e-06 
0.0 -0.6606 0 2.0 1e-06 
0.0 -0.6605 0 2.0 1e-06 
0.0 -0.6604 0 2.0 1e-06 
0.0 -0.6603 0 2.0 1e-06 
0.0 -0.6602 0 2.0 1e-06 
0.0 -0.6601 0 2.0 1e-06 
0.0 -0.66 0 2.0 1e-06 
0.0 -0.6599 0 2.0 1e-06 
0.0 -0.6598 0 2.0 1e-06 
0.0 -0.6597 0 2.0 1e-06 
0.0 -0.6596 0 2.0 1e-06 
0.0 -0.6595 0 2.0 1e-06 
0.0 -0.6594 0 2.0 1e-06 
0.0 -0.6593 0 2.0 1e-06 
0.0 -0.6592 0 2.0 1e-06 
0.0 -0.6591 0 2.0 1e-06 
0.0 -0.659 0 2.0 1e-06 
0.0 -0.6589 0 2.0 1e-06 
0.0 -0.6588 0 2.0 1e-06 
0.0 -0.6587 0 2.0 1e-06 
0.0 -0.6586 0 2.0 1e-06 
0.0 -0.6585 0 2.0 1e-06 
0.0 -0.6584 0 2.0 1e-06 
0.0 -0.6583 0 2.0 1e-06 
0.0 -0.6582 0 2.0 1e-06 
0.0 -0.6581 0 2.0 1e-06 
0.0 -0.658 0 2.0 1e-06 
0.0 -0.6579 0 2.0 1e-06 
0.0 -0.6578 0 2.0 1e-06 
0.0 -0.6577 0 2.0 1e-06 
0.0 -0.6576 0 2.0 1e-06 
0.0 -0.6575 0 2.0 1e-06 
0.0 -0.6574 0 2.0 1e-06 
0.0 -0.6573 0 2.0 1e-06 
0.0 -0.6572 0 2.0 1e-06 
0.0 -0.6571 0 2.0 1e-06 
0.0 -0.657 0 2.0 1e-06 
0.0 -0.6569 0 2.0 1e-06 
0.0 -0.6568 0 2.0 1e-06 
0.0 -0.6567 0 2.0 1e-06 
0.0 -0.6566 0 2.0 1e-06 
0.0 -0.6565 0 2.0 1e-06 
0.0 -0.6564 0 2.0 1e-06 
0.0 -0.6563 0 2.0 1e-06 
0.0 -0.6562 0 2.0 1e-06 
0.0 -0.6561 0 2.0 1e-06 
0.0 -0.656 0 2.0 1e-06 
0.0 -0.6559 0 2.0 1e-06 
0.0 -0.6558 0 2.0 1e-06 
0.0 -0.6557 0 2.0 1e-06 
0.0 -0.6556 0 2.0 1e-06 
0.0 -0.6555 0 2.0 1e-06 
0.0 -0.6554 0 2.0 1e-06 
0.0 -0.6553 0 2.0 1e-06 
0.0 -0.6552 0 2.0 1e-06 
0.0 -0.6551 0 2.0 1e-06 
0.0 -0.655 0 2.0 1e-06 
0.0 -0.6549 0 2.0 1e-06 
0.0 -0.6548 0 2.0 1e-06 
0.0 -0.6547 0 2.0 1e-06 
0.0 -0.6546 0 2.0 1e-06 
0.0 -0.6545 0 2.0 1e-06 
0.0 -0.6544 0 2.0 1e-06 
0.0 -0.6543 0 2.0 1e-06 
0.0 -0.6542 0 2.0 1e-06 
0.0 -0.6541 0 2.0 1e-06 
0.0 -0.654 0 2.0 1e-06 
0.0 -0.6539 0 2.0 1e-06 
0.0 -0.6538 0 2.0 1e-06 
0.0 -0.6537 0 2.0 1e-06 
0.0 -0.6536 0 2.0 1e-06 
0.0 -0.6535 0 2.0 1e-06 
0.0 -0.6534 0 2.0 1e-06 
0.0 -0.6533 0 2.0 1e-06 
0.0 -0.6532 0 2.0 1e-06 
0.0 -0.6531 0 2.0 1e-06 
0.0 -0.653 0 2.0 1e-06 
0.0 -0.6529 0 2.0 1e-06 
0.0 -0.6528 0 2.0 1e-06 
0.0 -0.6527 0 2.0 1e-06 
0.0 -0.6526 0 2.0 1e-06 
0.0 -0.6525 0 2.0 1e-06 
0.0 -0.6524 0 2.0 1e-06 
0.0 -0.6523 0 2.0 1e-06 
0.0 -0.6522 0 2.0 1e-06 
0.0 -0.6521 0 2.0 1e-06 
0.0 -0.652 0 2.0 1e-06 
0.0 -0.6519 0 2.0 1e-06 
0.0 -0.6518 0 2.0 1e-06 
0.0 -0.6517 0 2.0 1e-06 
0.0 -0.6516 0 2.0 1e-06 
0.0 -0.6515 0 2.0 1e-06 
0.0 -0.6514 0 2.0 1e-06 
0.0 -0.6513 0 2.0 1e-06 
0.0 -0.6512 0 2.0 1e-06 
0.0 -0.6511 0 2.0 1e-06 
0.0 -0.651 0 2.0 1e-06 
0.0 -0.6509 0 2.0 1e-06 
0.0 -0.6508 0 2.0 1e-06 
0.0 -0.6507 0 2.0 1e-06 
0.0 -0.6506 0 2.0 1e-06 
0.0 -0.6505 0 2.0 1e-06 
0.0 -0.6504 0 2.0 1e-06 
0.0 -0.6503 0 2.0 1e-06 
0.0 -0.6502 0 2.0 1e-06 
0.0 -0.6501 0 2.0 1e-06 
0.0 -0.65 0 2.0 1e-06 
0.0 -0.6499 0 2.0 1e-06 
0.0 -0.6498 0 2.0 1e-06 
0.0 -0.6497 0 2.0 1e-06 
0.0 -0.6496 0 2.0 1e-06 
0.0 -0.6495 0 2.0 1e-06 
0.0 -0.6494 0 2.0 1e-06 
0.0 -0.6493 0 2.0 1e-06 
0.0 -0.6492 0 2.0 1e-06 
0.0 -0.6491 0 2.0 1e-06 
0.0 -0.649 0 2.0 1e-06 
0.0 -0.6489 0 2.0 1e-06 
0.0 -0.6488 0 2.0 1e-06 
0.0 -0.6487 0 2.0 1e-06 
0.0 -0.6486 0 2.0 1e-06 
0.0 -0.6485 0 2.0 1e-06 
0.0 -0.6484 0 2.0 1e-06 
0.0 -0.6483 0 2.0 1e-06 
0.0 -0.6482 0 2.0 1e-06 
0.0 -0.6481 0 2.0 1e-06 
0.0 -0.648 0 2.0 1e-06 
0.0 -0.6479 0 2.0 1e-06 
0.0 -0.6478 0 2.0 1e-06 
0.0 -0.6477 0 2.0 1e-06 
0.0 -0.6476 0 2.0 1e-06 
0.0 -0.6475 0 2.0 1e-06 
0.0 -0.6474 0 2.0 1e-06 
0.0 -0.6473 0 2.0 1e-06 
0.0 -0.6472 0 2.0 1e-06 
0.0 -0.6471 0 2.0 1e-06 
0.0 -0.647 0 2.0 1e-06 
0.0 -0.6469 0 2.0 1e-06 
0.0 -0.6468 0 2.0 1e-06 
0.0 -0.6467 0 2.0 1e-06 
0.0 -0.6466 0 2.0 1e-06 
0.0 -0.6465 0 2.0 1e-06 
0.0 -0.6464 0 2.0 1e-06 
0.0 -0.6463 0 2.0 1e-06 
0.0 -0.6462 0 2.0 1e-06 
0.0 -0.6461 0 2.0 1e-06 
0.0 -0.646 0 2.0 1e-06 
0.0 -0.6459 0 2.0 1e-06 
0.0 -0.6458 0 2.0 1e-06 
0.0 -0.6457 0 2.0 1e-06 
0.0 -0.6456 0 2.0 1e-06 
0.0 -0.6455 0 2.0 1e-06 
0.0 -0.6454 0 2.0 1e-06 
0.0 -0.6453 0 2.0 1e-06 
0.0 -0.6452 0 2.0 1e-06 
0.0 -0.6451 0 2.0 1e-06 
0.0 -0.645 0 2.0 1e-06 
0.0 -0.6449 0 2.0 1e-06 
0.0 -0.6448 0 2.0 1e-06 
0.0 -0.6447 0 2.0 1e-06 
0.0 -0.6446 0 2.0 1e-06 
0.0 -0.6445 0 2.0 1e-06 
0.0 -0.6444 0 2.0 1e-06 
0.0 -0.6443 0 2.0 1e-06 
0.0 -0.6442 0 2.0 1e-06 
0.0 -0.6441 0 2.0 1e-06 
0.0 -0.644 0 2.0 1e-06 
0.0 -0.6439 0 2.0 1e-06 
0.0 -0.6438 0 2.0 1e-06 
0.0 -0.6437 0 2.0 1e-06 
0.0 -0.6436 0 2.0 1e-06 
0.0 -0.6435 0 2.0 1e-06 
0.0 -0.6434 0 2.0 1e-06 
0.0 -0.6433 0 2.0 1e-06 
0.0 -0.6432 0 2.0 1e-06 
0.0 -0.6431 0 2.0 1e-06 
0.0 -0.643 0 2.0 1e-06 
0.0 -0.6429 0 2.0 1e-06 
0.0 -0.6428 0 2.0 1e-06 
0.0 -0.6427 0 2.0 1e-06 
0.0 -0.6426 0 2.0 1e-06 
0.0 -0.6425 0 2.0 1e-06 
0.0 -0.6424 0 2.0 1e-06 
0.0 -0.6423 0 2.0 1e-06 
0.0 -0.6422 0 2.0 1e-06 
0.0 -0.6421 0 2.0 1e-06 
0.0 -0.642 0 2.0 1e-06 
0.0 -0.6419 0 2.0 1e-06 
0.0 -0.6418 0 2.0 1e-06 
0.0 -0.6417 0 2.0 1e-06 
0.0 -0.6416 0 2.0 1e-06 
0.0 -0.6415 0 2.0 1e-06 
0.0 -0.6414 0 2.0 1e-06 
0.0 -0.6413 0 2.0 1e-06 
0.0 -0.6412 0 2.0 1e-06 
0.0 -0.6411 0 2.0 1e-06 
0.0 -0.641 0 2.0 1e-06 
0.0 -0.6409 0 2.0 1e-06 
0.0 -0.6408 0 2.0 1e-06 
0.0 -0.6407 0 2.0 1e-06 
0.0 -0.6406 0 2.0 1e-06 
0.0 -0.6405 0 2.0 1e-06 
0.0 -0.6404 0 2.0 1e-06 
0.0 -0.6403 0 2.0 1e-06 
0.0 -0.6402 0 2.0 1e-06 
0.0 -0.6401 0 2.0 1e-06 
0.0 -0.64 0 2.0 1e-06 
0.0 -0.6399 0 2.0 1e-06 
0.0 -0.6398 0 2.0 1e-06 
0.0 -0.6397 0 2.0 1e-06 
0.0 -0.6396 0 2.0 1e-06 
0.0 -0.6395 0 2.0 1e-06 
0.0 -0.6394 0 2.0 1e-06 
0.0 -0.6393 0 2.0 1e-06 
0.0 -0.6392 0 2.0 1e-06 
0.0 -0.6391 0 2.0 1e-06 
0.0 -0.639 0 2.0 1e-06 
0.0 -0.6389 0 2.0 1e-06 
0.0 -0.6388 0 2.0 1e-06 
0.0 -0.6387 0 2.0 1e-06 
0.0 -0.6386 0 2.0 1e-06 
0.0 -0.6385 0 2.0 1e-06 
0.0 -0.6384 0 2.0 1e-06 
0.0 -0.6383 0 2.0 1e-06 
0.0 -0.6382 0 2.0 1e-06 
0.0 -0.6381 0 2.0 1e-06 
0.0 -0.638 0 2.0 1e-06 
0.0 -0.6379 0 2.0 1e-06 
0.0 -0.6378 0 2.0 1e-06 
0.0 -0.6377 0 2.0 1e-06 
0.0 -0.6376 0 2.0 1e-06 
0.0 -0.6375 0 2.0 1e-06 
0.0 -0.6374 0 2.0 1e-06 
0.0 -0.6373 0 2.0 1e-06 
0.0 -0.6372 0 2.0 1e-06 
0.0 -0.6371 0 2.0 1e-06 
0.0 -0.637 0 2.0 1e-06 
0.0 -0.6369 0 2.0 1e-06 
0.0 -0.6368 0 2.0 1e-06 
0.0 -0.6367 0 2.0 1e-06 
0.0 -0.6366 0 2.0 1e-06 
0.0 -0.6365 0 2.0 1e-06 
0.0 -0.6364 0 2.0 1e-06 
0.0 -0.6363 0 2.0 1e-06 
0.0 -0.6362 0 2.0 1e-06 
0.0 -0.6361 0 2.0 1e-06 
0.0 -0.636 0 2.0 1e-06 
0.0 -0.6359 0 2.0 1e-06 
0.0 -0.6358 0 2.0 1e-06 
0.0 -0.6357 0 2.0 1e-06 
0.0 -0.6356 0 2.0 1e-06 
0.0 -0.6355 0 2.0 1e-06 
0.0 -0.6354 0 2.0 1e-06 
0.0 -0.6353 0 2.0 1e-06 
0.0 -0.6352 0 2.0 1e-06 
0.0 -0.6351 0 2.0 1e-06 
0.0 -0.635 0 2.0 1e-06 
0.0 -0.6349 0 2.0 1e-06 
0.0 -0.6348 0 2.0 1e-06 
0.0 -0.6347 0 2.0 1e-06 
0.0 -0.6346 0 2.0 1e-06 
0.0 -0.6345 0 2.0 1e-06 
0.0 -0.6344 0 2.0 1e-06 
0.0 -0.6343 0 2.0 1e-06 
0.0 -0.6342 0 2.0 1e-06 
0.0 -0.6341 0 2.0 1e-06 
0.0 -0.634 0 2.0 1e-06 
0.0 -0.6339 0 2.0 1e-06 
0.0 -0.6338 0 2.0 1e-06 
0.0 -0.6337 0 2.0 1e-06 
0.0 -0.6336 0 2.0 1e-06 
0.0 -0.6335 0 2.0 1e-06 
0.0 -0.6334 0 2.0 1e-06 
0.0 -0.6333 0 2.0 1e-06 
0.0 -0.6332 0 2.0 1e-06 
0.0 -0.6331 0 2.0 1e-06 
0.0 -0.633 0 2.0 1e-06 
0.0 -0.6329 0 2.0 1e-06 
0.0 -0.6328 0 2.0 1e-06 
0.0 -0.6327 0 2.0 1e-06 
0.0 -0.6326 0 2.0 1e-06 
0.0 -0.6325 0 2.0 1e-06 
0.0 -0.6324 0 2.0 1e-06 
0.0 -0.6323 0 2.0 1e-06 
0.0 -0.6322 0 2.0 1e-06 
0.0 -0.6321 0 2.0 1e-06 
0.0 -0.632 0 2.0 1e-06 
0.0 -0.6319 0 2.0 1e-06 
0.0 -0.6318 0 2.0 1e-06 
0.0 -0.6317 0 2.0 1e-06 
0.0 -0.6316 0 2.0 1e-06 
0.0 -0.6315 0 2.0 1e-06 
0.0 -0.6314 0 2.0 1e-06 
0.0 -0.6313 0 2.0 1e-06 
0.0 -0.6312 0 2.0 1e-06 
0.0 -0.6311 0 2.0 1e-06 
0.0 -0.631 0 2.0 1e-06 
0.0 -0.6309 0 2.0 1e-06 
0.0 -0.6308 0 2.0 1e-06 
0.0 -0.6307 0 2.0 1e-06 
0.0 -0.6306 0 2.0 1e-06 
0.0 -0.6305 0 2.0 1e-06 
0.0 -0.6304 0 2.0 1e-06 
0.0 -0.6303 0 2.0 1e-06 
0.0 -0.6302 0 2.0 1e-06 
0.0 -0.6301 0 2.0 1e-06 
0.0 -0.63 0 2.0 1e-06 
0.0 -0.6299 0 2.0 1e-06 
0.0 -0.6298 0 2.0 1e-06 
0.0 -0.6297 0 2.0 1e-06 
0.0 -0.6296 0 2.0 1e-06 
0.0 -0.6295 0 2.0 1e-06 
0.0 -0.6294 0 2.0 1e-06 
0.0 -0.6293 0 2.0 1e-06 
0.0 -0.6292 0 2.0 1e-06 
0.0 -0.6291 0 2.0 1e-06 
0.0 -0.629 0 2.0 1e-06 
0.0 -0.6289 0 2.0 1e-06 
0.0 -0.6288 0 2.0 1e-06 
0.0 -0.6287 0 2.0 1e-06 
0.0 -0.6286 0 2.0 1e-06 
0.0 -0.6285 0 2.0 1e-06 
0.0 -0.6284 0 2.0 1e-06 
0.0 -0.6283 0 2.0 1e-06 
0.0 -0.6282 0 2.0 1e-06 
0.0 -0.6281 0 2.0 1e-06 
0.0 -0.628 0 2.0 1e-06 
0.0 -0.6279 0 2.0 1e-06 
0.0 -0.6278 0 2.0 1e-06 
0.0 -0.6277 0 2.0 1e-06 
0.0 -0.6276 0 2.0 1e-06 
0.0 -0.6275 0 2.0 1e-06 
0.0 -0.6274 0 2.0 1e-06 
0.0 -0.6273 0 2.0 1e-06 
0.0 -0.6272 0 2.0 1e-06 
0.0 -0.6271 0 2.0 1e-06 
0.0 -0.627 0 2.0 1e-06 
0.0 -0.6269 0 2.0 1e-06 
0.0 -0.6268 0 2.0 1e-06 
0.0 -0.6267 0 2.0 1e-06 
0.0 -0.6266 0 2.0 1e-06 
0.0 -0.6265 0 2.0 1e-06 
0.0 -0.6264 0 2.0 1e-06 
0.0 -0.6263 0 2.0 1e-06 
0.0 -0.6262 0 2.0 1e-06 
0.0 -0.6261 0 2.0 1e-06 
0.0 -0.626 0 2.0 1e-06 
0.0 -0.6259 0 2.0 1e-06 
0.0 -0.6258 0 2.0 1e-06 
0.0 -0.6257 0 2.0 1e-06 
0.0 -0.6256 0 2.0 1e-06 
0.0 -0.6255 0 2.0 1e-06 
0.0 -0.6254 0 2.0 1e-06 
0.0 -0.6253 0 2.0 1e-06 
0.0 -0.6252 0 2.0 1e-06 
0.0 -0.6251 0 2.0 1e-06 
0.0 -0.625 0 2.0 1e-06 
0.0 -0.6249 0 2.0 1e-06 
0.0 -0.6248 0 2.0 1e-06 
0.0 -0.6247 0 2.0 1e-06 
0.0 -0.6246 0 2.0 1e-06 
0.0 -0.6245 0 2.0 1e-06 
0.0 -0.6244 0 2.0 1e-06 
0.0 -0.6243 0 2.0 1e-06 
0.0 -0.6242 0 2.0 1e-06 
0.0 -0.6241 0 2.0 1e-06 
0.0 -0.624 0 2.0 1e-06 
0.0 -0.6239 0 2.0 1e-06 
0.0 -0.6238 0 2.0 1e-06 
0.0 -0.6237 0 2.0 1e-06 
0.0 -0.6236 0 2.0 1e-06 
0.0 -0.6235 0 2.0 1e-06 
0.0 -0.6234 0 2.0 1e-06 
0.0 -0.6233 0 2.0 1e-06 
0.0 -0.6232 0 2.0 1e-06 
0.0 -0.6231 0 2.0 1e-06 
0.0 -0.623 0 2.0 1e-06 
0.0 -0.6229 0 2.0 1e-06 
0.0 -0.6228 0 2.0 1e-06 
0.0 -0.6227 0 2.0 1e-06 
0.0 -0.6226 0 2.0 1e-06 
0.0 -0.6225 0 2.0 1e-06 
0.0 -0.6224 0 2.0 1e-06 
0.0 -0.6223 0 2.0 1e-06 
0.0 -0.6222 0 2.0 1e-06 
0.0 -0.6221 0 2.0 1e-06 
0.0 -0.622 0 2.0 1e-06 
0.0 -0.6219 0 2.0 1e-06 
0.0 -0.6218 0 2.0 1e-06 
0.0 -0.6217 0 2.0 1e-06 
0.0 -0.6216 0 2.0 1e-06 
0.0 -0.6215 0 2.0 1e-06 
0.0 -0.6214 0 2.0 1e-06 
0.0 -0.6213 0 2.0 1e-06 
0.0 -0.6212 0 2.0 1e-06 
0.0 -0.6211 0 2.0 1e-06 
0.0 -0.621 0 2.0 1e-06 
0.0 -0.6209 0 2.0 1e-06 
0.0 -0.6208 0 2.0 1e-06 
0.0 -0.6207 0 2.0 1e-06 
0.0 -0.6206 0 2.0 1e-06 
0.0 -0.6205 0 2.0 1e-06 
0.0 -0.6204 0 2.0 1e-06 
0.0 -0.6203 0 2.0 1e-06 
0.0 -0.6202 0 2.0 1e-06 
0.0 -0.6201 0 2.0 1e-06 
0.0 -0.62 0 2.0 1e-06 
0.0 -0.6199 0 2.0 1e-06 
0.0 -0.6198 0 2.0 1e-06 
0.0 -0.6197 0 2.0 1e-06 
0.0 -0.6196 0 2.0 1e-06 
0.0 -0.6195 0 2.0 1e-06 
0.0 -0.6194 0 2.0 1e-06 
0.0 -0.6193 0 2.0 1e-06 
0.0 -0.6192 0 2.0 1e-06 
0.0 -0.6191 0 2.0 1e-06 
0.0 -0.619 0 2.0 1e-06 
0.0 -0.6189 0 2.0 1e-06 
0.0 -0.6188 0 2.0 1e-06 
0.0 -0.6187 0 2.0 1e-06 
0.0 -0.6186 0 2.0 1e-06 
0.0 -0.6185 0 2.0 1e-06 
0.0 -0.6184 0 2.0 1e-06 
0.0 -0.6183 0 2.0 1e-06 
0.0 -0.6182 0 2.0 1e-06 
0.0 -0.6181 0 2.0 1e-06 
0.0 -0.618 0 2.0 1e-06 
0.0 -0.6179 0 2.0 1e-06 
0.0 -0.6178 0 2.0 1e-06 
0.0 -0.6177 0 2.0 1e-06 
0.0 -0.6176 0 2.0 1e-06 
0.0 -0.6175 0 2.0 1e-06 
0.0 -0.6174 0 2.0 1e-06 
0.0 -0.6173 0 2.0 1e-06 
0.0 -0.6172 0 2.0 1e-06 
0.0 -0.6171 0 2.0 1e-06 
0.0 -0.617 0 2.0 1e-06 
0.0 -0.6169 0 2.0 1e-06 
0.0 -0.6168 0 2.0 1e-06 
0.0 -0.6167 0 2.0 1e-06 
0.0 -0.6166 0 2.0 1e-06 
0.0 -0.6165 0 2.0 1e-06 
0.0 -0.6164 0 2.0 1e-06 
0.0 -0.6163 0 2.0 1e-06 
0.0 -0.6162 0 2.0 1e-06 
0.0 -0.6161 0 2.0 1e-06 
0.0 -0.616 0 2.0 1e-06 
0.0 -0.6159 0 2.0 1e-06 
0.0 -0.6158 0 2.0 1e-06 
0.0 -0.6157 0 2.0 1e-06 
0.0 -0.6156 0 2.0 1e-06 
0.0 -0.6155 0 2.0 1e-06 
0.0 -0.6154 0 2.0 1e-06 
0.0 -0.6153 0 2.0 1e-06 
0.0 -0.6152 0 2.0 1e-06 
0.0 -0.6151 0 2.0 1e-06 
0.0 -0.615 0 2.0 1e-06 
0.0 -0.6149 0 2.0 1e-06 
0.0 -0.6148 0 2.0 1e-06 
0.0 -0.6147 0 2.0 1e-06 
0.0 -0.6146 0 2.0 1e-06 
0.0 -0.6145 0 2.0 1e-06 
0.0 -0.6144 0 2.0 1e-06 
0.0 -0.6143 0 2.0 1e-06 
0.0 -0.6142 0 2.0 1e-06 
0.0 -0.6141 0 2.0 1e-06 
0.0 -0.614 0 2.0 1e-06 
0.0 -0.6139 0 2.0 1e-06 
0.0 -0.6138 0 2.0 1e-06 
0.0 -0.6137 0 2.0 1e-06 
0.0 -0.6136 0 2.0 1e-06 
0.0 -0.6135 0 2.0 1e-06 
0.0 -0.6134 0 2.0 1e-06 
0.0 -0.6133 0 2.0 1e-06 
0.0 -0.6132 0 2.0 1e-06 
0.0 -0.6131 0 2.0 1e-06 
0.0 -0.613 0 2.0 1e-06 
0.0 -0.6129 0 2.0 1e-06 
0.0 -0.6128 0 2.0 1e-06 
0.0 -0.6127 0 2.0 1e-06 
0.0 -0.6126 0 2.0 1e-06 
0.0 -0.6125 0 2.0 1e-06 
0.0 -0.6124 0 2.0 1e-06 
0.0 -0.6123 0 2.0 1e-06 
0.0 -0.6122 0 2.0 1e-06 
0.0 -0.6121 0 2.0 1e-06 
0.0 -0.612 0 2.0 1e-06 
0.0 -0.6119 0 2.0 1e-06 
0.0 -0.6118 0 2.0 1e-06 
0.0 -0.6117 0 2.0 1e-06 
0.0 -0.6116 0 2.0 1e-06 
0.0 -0.6115 0 2.0 1e-06 
0.0 -0.6114 0 2.0 1e-06 
0.0 -0.6113 0 2.0 1e-06 
0.0 -0.6112 0 2.0 1e-06 
0.0 -0.6111 0 2.0 1e-06 
0.0 -0.611 0 2.0 1e-06 
0.0 -0.6109 0 2.0 1e-06 
0.0 -0.6108 0 2.0 1e-06 
0.0 -0.6107 0 2.0 1e-06 
0.0 -0.6106 0 2.0 1e-06 
0.0 -0.6105 0 2.0 1e-06 
0.0 -0.6104 0 2.0 1e-06 
0.0 -0.6103 0 2.0 1e-06 
0.0 -0.6102 0 2.0 1e-06 
0.0 -0.6101 0 2.0 1e-06 
0.0 -0.61 0 2.0 1e-06 
0.0 -0.6099 0 2.0 1e-06 
0.0 -0.6098 0 2.0 1e-06 
0.0 -0.6097 0 2.0 1e-06 
0.0 -0.6096 0 2.0 1e-06 
0.0 -0.6095 0 2.0 1e-06 
0.0 -0.6094 0 2.0 1e-06 
0.0 -0.6093 0 2.0 1e-06 
0.0 -0.6092 0 2.0 1e-06 
0.0 -0.6091 0 2.0 1e-06 
0.0 -0.609 0 2.0 1e-06 
0.0 -0.6089 0 2.0 1e-06 
0.0 -0.6088 0 2.0 1e-06 
0.0 -0.6087 0 2.0 1e-06 
0.0 -0.6086 0 2.0 1e-06 
0.0 -0.6085 0 2.0 1e-06 
0.0 -0.6084 0 2.0 1e-06 
0.0 -0.6083 0 2.0 1e-06 
0.0 -0.6082 0 2.0 1e-06 
0.0 -0.6081 0 2.0 1e-06 
0.0 -0.608 0 2.0 1e-06 
0.0 -0.6079 0 2.0 1e-06 
0.0 -0.6078 0 2.0 1e-06 
0.0 -0.6077 0 2.0 1e-06 
0.0 -0.6076 0 2.0 1e-06 
0.0 -0.6075 0 2.0 1e-06 
0.0 -0.6074 0 2.0 1e-06 
0.0 -0.6073 0 2.0 1e-06 
0.0 -0.6072 0 2.0 1e-06 
0.0 -0.6071 0 2.0 1e-06 
0.0 -0.607 0 2.0 1e-06 
0.0 -0.6069 0 2.0 1e-06 
0.0 -0.6068 0 2.0 1e-06 
0.0 -0.6067 0 2.0 1e-06 
0.0 -0.6066 0 2.0 1e-06 
0.0 -0.6065 0 2.0 1e-06 
0.0 -0.6064 0 2.0 1e-06 
0.0 -0.6063 0 2.0 1e-06 
0.0 -0.6062 0 2.0 1e-06 
0.0 -0.6061 0 2.0 1e-06 
0.0 -0.606 0 2.0 1e-06 
0.0 -0.6059 0 2.0 1e-06 
0.0 -0.6058 0 2.0 1e-06 
0.0 -0.6057 0 2.0 1e-06 
0.0 -0.6056 0 2.0 1e-06 
0.0 -0.6055 0 2.0 1e-06 
0.0 -0.6054 0 2.0 1e-06 
0.0 -0.6053 0 2.0 1e-06 
0.0 -0.6052 0 2.0 1e-06 
0.0 -0.6051 0 2.0 1e-06 
0.0 -0.605 0 2.0 1e-06 
0.0 -0.6049 0 2.0 1e-06 
0.0 -0.6048 0 2.0 1e-06 
0.0 -0.6047 0 2.0 1e-06 
0.0 -0.6046 0 2.0 1e-06 
0.0 -0.6045 0 2.0 1e-06 
0.0 -0.6044 0 2.0 1e-06 
0.0 -0.6043 0 2.0 1e-06 
0.0 -0.6042 0 2.0 1e-06 
0.0 -0.6041 0 2.0 1e-06 
0.0 -0.604 0 2.0 1e-06 
0.0 -0.6039 0 2.0 1e-06 
0.0 -0.6038 0 2.0 1e-06 
0.0 -0.6037 0 2.0 1e-06 
0.0 -0.6036 0 2.0 1e-06 
0.0 -0.6035 0 2.0 1e-06 
0.0 -0.6034 0 2.0 1e-06 
0.0 -0.6033 0 2.0 1e-06 
0.0 -0.6032 0 2.0 1e-06 
0.0 -0.6031 0 2.0 1e-06 
0.0 -0.603 0 2.0 1e-06 
0.0 -0.6029 0 2.0 1e-06 
0.0 -0.6028 0 2.0 1e-06 
0.0 -0.6027 0 2.0 1e-06 
0.0 -0.6026 0 2.0 1e-06 
0.0 -0.6025 0 2.0 1e-06 
0.0 -0.6024 0 2.0 1e-06 
0.0 -0.6023 0 2.0 1e-06 
0.0 -0.6022 0 2.0 1e-06 
0.0 -0.6021 0 2.0 1e-06 
0.0 -0.602 0 2.0 1e-06 
0.0 -0.6019 0 2.0 1e-06 
0.0 -0.6018 0 2.0 1e-06 
0.0 -0.6017 0 2.0 1e-06 
0.0 -0.6016 0 2.0 1e-06 
0.0 -0.6015 0 2.0 1e-06 
0.0 -0.6014 0 2.0 1e-06 
0.0 -0.6013 0 2.0 1e-06 
0.0 -0.6012 0 2.0 1e-06 
0.0 -0.6011 0 2.0 1e-06 
0.0 -0.601 0 2.0 1e-06 
0.0 -0.6009 0 2.0 1e-06 
0.0 -0.6008 0 2.0 1e-06 
0.0 -0.6007 0 2.0 1e-06 
0.0 -0.6006 0 2.0 1e-06 
0.0 -0.6005 0 2.0 1e-06 
0.0 -0.6004 0 2.0 1e-06 
0.0 -0.6003 0 2.0 1e-06 
0.0 -0.6002 0 2.0 1e-06 
0.0 -0.6001 0 2.0 1e-06 
0.0 -0.6 0 2.0 1e-06 
0.0 -0.5999 0 2.0 1e-06 
0.0 -0.5998 0 2.0 1e-06 
0.0 -0.5997 0 2.0 1e-06 
0.0 -0.5996 0 2.0 1e-06 
0.0 -0.5995 0 2.0 1e-06 
0.0 -0.5994 0 2.0 1e-06 
0.0 -0.5993 0 2.0 1e-06 
0.0 -0.5992 0 2.0 1e-06 
0.0 -0.5991 0 2.0 1e-06 
0.0 -0.599 0 2.0 1e-06 
0.0 -0.5989 0 2.0 1e-06 
0.0 -0.5988 0 2.0 1e-06 
0.0 -0.5987 0 2.0 1e-06 
0.0 -0.5986 0 2.0 1e-06 
0.0 -0.5985 0 2.0 1e-06 
0.0 -0.5984 0 2.0 1e-06 
0.0 -0.5983 0 2.0 1e-06 
0.0 -0.5982 0 2.0 1e-06 
0.0 -0.5981 0 2.0 1e-06 
0.0 -0.598 0 2.0 1e-06 
0.0 -0.5979 0 2.0 1e-06 
0.0 -0.5978 0 2.0 1e-06 
0.0 -0.5977 0 2.0 1e-06 
0.0 -0.5976 0 2.0 1e-06 
0.0 -0.5975 0 2.0 1e-06 
0.0 -0.5974 0 2.0 1e-06 
0.0 -0.5973 0 2.0 1e-06 
0.0 -0.5972 0 2.0 1e-06 
0.0 -0.5971 0 2.0 1e-06 
0.0 -0.597 0 2.0 1e-06 
0.0 -0.5969 0 2.0 1e-06 
0.0 -0.5968 0 2.0 1e-06 
0.0 -0.5967 0 2.0 1e-06 
0.0 -0.5966 0 2.0 1e-06 
0.0 -0.5965 0 2.0 1e-06 
0.0 -0.5964 0 2.0 1e-06 
0.0 -0.5963 0 2.0 1e-06 
0.0 -0.5962 0 2.0 1e-06 
0.0 -0.5961 0 2.0 1e-06 
0.0 -0.596 0 2.0 1e-06 
0.0 -0.5959 0 2.0 1e-06 
0.0 -0.5958 0 2.0 1e-06 
0.0 -0.5957 0 2.0 1e-06 
0.0 -0.5956 0 2.0 1e-06 
0.0 -0.5955 0 2.0 1e-06 
0.0 -0.5954 0 2.0 1e-06 
0.0 -0.5953 0 2.0 1e-06 
0.0 -0.5952 0 2.0 1e-06 
0.0 -0.5951 0 2.0 1e-06 
0.0 -0.595 0 2.0 1e-06 
0.0 -0.5949 0 2.0 1e-06 
0.0 -0.5948 0 2.0 1e-06 
0.0 -0.5947 0 2.0 1e-06 
0.0 -0.5946 0 2.0 1e-06 
0.0 -0.5945 0 2.0 1e-06 
0.0 -0.5944 0 2.0 1e-06 
0.0 -0.5943 0 2.0 1e-06 
0.0 -0.5942 0 2.0 1e-06 
0.0 -0.5941 0 2.0 1e-06 
0.0 -0.594 0 2.0 1e-06 
0.0 -0.5939 0 2.0 1e-06 
0.0 -0.5938 0 2.0 1e-06 
0.0 -0.5937 0 2.0 1e-06 
0.0 -0.5936 0 2.0 1e-06 
0.0 -0.5935 0 2.0 1e-06 
0.0 -0.5934 0 2.0 1e-06 
0.0 -0.5933 0 2.0 1e-06 
0.0 -0.5932 0 2.0 1e-06 
0.0 -0.5931 0 2.0 1e-06 
0.0 -0.593 0 2.0 1e-06 
0.0 -0.5929 0 2.0 1e-06 
0.0 -0.5928 0 2.0 1e-06 
0.0 -0.5927 0 2.0 1e-06 
0.0 -0.5926 0 2.0 1e-06 
0.0 -0.5925 0 2.0 1e-06 
0.0 -0.5924 0 2.0 1e-06 
0.0 -0.5923 0 2.0 1e-06 
0.0 -0.5922 0 2.0 1e-06 
0.0 -0.5921 0 2.0 1e-06 
0.0 -0.592 0 2.0 1e-06 
0.0 -0.5919 0 2.0 1e-06 
0.0 -0.5918 0 2.0 1e-06 
0.0 -0.5917 0 2.0 1e-06 
0.0 -0.5916 0 2.0 1e-06 
0.0 -0.5915 0 2.0 1e-06 
0.0 -0.5914 0 2.0 1e-06 
0.0 -0.5913 0 2.0 1e-06 
0.0 -0.5912 0 2.0 1e-06 
0.0 -0.5911 0 2.0 1e-06 
0.0 -0.591 0 2.0 1e-06 
0.0 -0.5909 0 2.0 1e-06 
0.0 -0.5908 0 2.0 1e-06 
0.0 -0.5907 0 2.0 1e-06 
0.0 -0.5906 0 2.0 1e-06 
0.0 -0.5905 0 2.0 1e-06 
0.0 -0.5904 0 2.0 1e-06 
0.0 -0.5903 0 2.0 1e-06 
0.0 -0.5902 0 2.0 1e-06 
0.0 -0.5901 0 2.0 1e-06 
0.0 -0.59 0 2.0 1e-06 
0.0 -0.5899 0 2.0 1e-06 
0.0 -0.5898 0 2.0 1e-06 
0.0 -0.5897 0 2.0 1e-06 
0.0 -0.5896 0 2.0 1e-06 
0.0 -0.5895 0 2.0 1e-06 
0.0 -0.5894 0 2.0 1e-06 
0.0 -0.5893 0 2.0 1e-06 
0.0 -0.5892 0 2.0 1e-06 
0.0 -0.5891 0 2.0 1e-06 
0.0 -0.589 0 2.0 1e-06 
0.0 -0.5889 0 2.0 1e-06 
0.0 -0.5888 0 2.0 1e-06 
0.0 -0.5887 0 2.0 1e-06 
0.0 -0.5886 0 2.0 1e-06 
0.0 -0.5885 0 2.0 1e-06 
0.0 -0.5884 0 2.0 1e-06 
0.0 -0.5883 0 2.0 1e-06 
0.0 -0.5882 0 2.0 1e-06 
0.0 -0.5881 0 2.0 1e-06 
0.0 -0.588 0 2.0 1e-06 
0.0 -0.5879 0 2.0 1e-06 
0.0 -0.5878 0 2.0 1e-06 
0.0 -0.5877 0 2.0 1e-06 
0.0 -0.5876 0 2.0 1e-06 
0.0 -0.5875 0 2.0 1e-06 
0.0 -0.5874 0 2.0 1e-06 
0.0 -0.5873 0 2.0 1e-06 
0.0 -0.5872 0 2.0 1e-06 
0.0 -0.5871 0 2.0 1e-06 
0.0 -0.587 0 2.0 1e-06 
0.0 -0.5869 0 2.0 1e-06 
0.0 -0.5868 0 2.0 1e-06 
0.0 -0.5867 0 2.0 1e-06 
0.0 -0.5866 0 2.0 1e-06 
0.0 -0.5865 0 2.0 1e-06 
0.0 -0.5864 0 2.0 1e-06 
0.0 -0.5863 0 2.0 1e-06 
0.0 -0.5862 0 2.0 1e-06 
0.0 -0.5861 0 2.0 1e-06 
0.0 -0.586 0 2.0 1e-06 
0.0 -0.5859 0 2.0 1e-06 
0.0 -0.5858 0 2.0 1e-06 
0.0 -0.5857 0 2.0 1e-06 
0.0 -0.5856 0 2.0 1e-06 
0.0 -0.5855 0 2.0 1e-06 
0.0 -0.5854 0 2.0 1e-06 
0.0 -0.5853 0 2.0 1e-06 
0.0 -0.5852 0 2.0 1e-06 
0.0 -0.5851 0 2.0 1e-06 
0.0 -0.585 0 2.0 1e-06 
0.0 -0.5849 0 2.0 1e-06 
0.0 -0.5848 0 2.0 1e-06 
0.0 -0.5847 0 2.0 1e-06 
0.0 -0.5846 0 2.0 1e-06 
0.0 -0.5845 0 2.0 1e-06 
0.0 -0.5844 0 2.0 1e-06 
0.0 -0.5843 0 2.0 1e-06 
0.0 -0.5842 0 2.0 1e-06 
0.0 -0.5841 0 2.0 1e-06 
0.0 -0.584 0 2.0 1e-06 
0.0 -0.5839 0 2.0 1e-06 
0.0 -0.5838 0 2.0 1e-06 
0.0 -0.5837 0 2.0 1e-06 
0.0 -0.5836 0 2.0 1e-06 
0.0 -0.5835 0 2.0 1e-06 
0.0 -0.5834 0 2.0 1e-06 
0.0 -0.5833 0 2.0 1e-06 
0.0 -0.5832 0 2.0 1e-06 
0.0 -0.5831 0 2.0 1e-06 
0.0 -0.583 0 2.0 1e-06 
0.0 -0.5829 0 2.0 1e-06 
0.0 -0.5828 0 2.0 1e-06 
0.0 -0.5827 0 2.0 1e-06 
0.0 -0.5826 0 2.0 1e-06 
0.0 -0.5825 0 2.0 1e-06 
0.0 -0.5824 0 2.0 1e-06 
0.0 -0.5823 0 2.0 1e-06 
0.0 -0.5822 0 2.0 1e-06 
0.0 -0.5821 0 2.0 1e-06 
0.0 -0.582 0 2.0 1e-06 
0.0 -0.5819 0 2.0 1e-06 
0.0 -0.5818 0 2.0 1e-06 
0.0 -0.5817 0 2.0 1e-06 
0.0 -0.5816 0 2.0 1e-06 
0.0 -0.5815 0 2.0 1e-06 
0.0 -0.5814 0 2.0 1e-06 
0.0 -0.5813 0 2.0 1e-06 
0.0 -0.5812 0 2.0 1e-06 
0.0 -0.5811 0 2.0 1e-06 
0.0 -0.581 0 2.0 1e-06 
0.0 -0.5809 0 2.0 1e-06 
0.0 -0.5808 0 2.0 1e-06 
0.0 -0.5807 0 2.0 1e-06 
0.0 -0.5806 0 2.0 1e-06 
0.0 -0.5805 0 2.0 1e-06 
0.0 -0.5804 0 2.0 1e-06 
0.0 -0.5803 0 2.0 1e-06 
0.0 -0.5802 0 2.0 1e-06 
0.0 -0.5801 0 2.0 1e-06 
0.0 -0.58 0 2.0 1e-06 
0.0 -0.5799 0 2.0 1e-06 
0.0 -0.5798 0 2.0 1e-06 
0.0 -0.5797 0 2.0 1e-06 
0.0 -0.5796 0 2.0 1e-06 
0.0 -0.5795 0 2.0 1e-06 
0.0 -0.5794 0 2.0 1e-06 
0.0 -0.5793 0 2.0 1e-06 
0.0 -0.5792 0 2.0 1e-06 
0.0 -0.5791 0 2.0 1e-06 
0.0 -0.579 0 2.0 1e-06 
0.0 -0.5789 0 2.0 1e-06 
0.0 -0.5788 0 2.0 1e-06 
0.0 -0.5787 0 2.0 1e-06 
0.0 -0.5786 0 2.0 1e-06 
0.0 -0.5785 0 2.0 1e-06 
0.0 -0.5784 0 2.0 1e-06 
0.0 -0.5783 0 2.0 1e-06 
0.0 -0.5782 0 2.0 1e-06 
0.0 -0.5781 0 2.0 1e-06 
0.0 -0.578 0 2.0 1e-06 
0.0 -0.5779 0 2.0 1e-06 
0.0 -0.5778 0 2.0 1e-06 
0.0 -0.5777 0 2.0 1e-06 
0.0 -0.5776 0 2.0 1e-06 
0.0 -0.5775 0 2.0 1e-06 
0.0 -0.5774 0 2.0 1e-06 
0.0 -0.5773 0 2.0 1e-06 
0.0 -0.5772 0 2.0 1e-06 
0.0 -0.5771 0 2.0 1e-06 
0.0 -0.577 0 2.0 1e-06 
0.0 -0.5769 0 2.0 1e-06 
0.0 -0.5768 0 2.0 1e-06 
0.0 -0.5767 0 2.0 1e-06 
0.0 -0.5766 0 2.0 1e-06 
0.0 -0.5765 0 2.0 1e-06 
0.0 -0.5764 0 2.0 1e-06 
0.0 -0.5763 0 2.0 1e-06 
0.0 -0.5762 0 2.0 1e-06 
0.0 -0.5761 0 2.0 1e-06 
0.0 -0.576 0 2.0 1e-06 
0.0 -0.5759 0 2.0 1e-06 
0.0 -0.5758 0 2.0 1e-06 
0.0 -0.5757 0 2.0 1e-06 
0.0 -0.5756 0 2.0 1e-06 
0.0 -0.5755 0 2.0 1e-06 
0.0 -0.5754 0 2.0 1e-06 
0.0 -0.5753 0 2.0 1e-06 
0.0 -0.5752 0 2.0 1e-06 
0.0 -0.5751 0 2.0 1e-06 
0.0 -0.575 0 2.0 1e-06 
0.0 -0.5749 0 2.0 1e-06 
0.0 -0.5748 0 2.0 1e-06 
0.0 -0.5747 0 2.0 1e-06 
0.0 -0.5746 0 2.0 1e-06 
0.0 -0.5745 0 2.0 1e-06 
0.0 -0.5744 0 2.0 1e-06 
0.0 -0.5743 0 2.0 1e-06 
0.0 -0.5742 0 2.0 1e-06 
0.0 -0.5741 0 2.0 1e-06 
0.0 -0.574 0 2.0 1e-06 
0.0 -0.5739 0 2.0 1e-06 
0.0 -0.5738 0 2.0 1e-06 
0.0 -0.5737 0 2.0 1e-06 
0.0 -0.5736 0 2.0 1e-06 
0.0 -0.5735 0 2.0 1e-06 
0.0 -0.5734 0 2.0 1e-06 
0.0 -0.5733 0 2.0 1e-06 
0.0 -0.5732 0 2.0 1e-06 
0.0 -0.5731 0 2.0 1e-06 
0.0 -0.573 0 2.0 1e-06 
0.0 -0.5729 0 2.0 1e-06 
0.0 -0.5728 0 2.0 1e-06 
0.0 -0.5727 0 2.0 1e-06 
0.0 -0.5726 0 2.0 1e-06 
0.0 -0.5725 0 2.0 1e-06 
0.0 -0.5724 0 2.0 1e-06 
0.0 -0.5723 0 2.0 1e-06 
0.0 -0.5722 0 2.0 1e-06 
0.0 -0.5721 0 2.0 1e-06 
0.0 -0.572 0 2.0 1e-06 
0.0 -0.5719 0 2.0 1e-06 
0.0 -0.5718 0 2.0 1e-06 
0.0 -0.5717 0 2.0 1e-06 
0.0 -0.5716 0 2.0 1e-06 
0.0 -0.5715 0 2.0 1e-06 
0.0 -0.5714 0 2.0 1e-06 
0.0 -0.5713 0 2.0 1e-06 
0.0 -0.5712 0 2.0 1e-06 
0.0 -0.5711 0 2.0 1e-06 
0.0 -0.571 0 2.0 1e-06 
0.0 -0.5709 0 2.0 1e-06 
0.0 -0.5708 0 2.0 1e-06 
0.0 -0.5707 0 2.0 1e-06 
0.0 -0.5706 0 2.0 1e-06 
0.0 -0.5705 0 2.0 1e-06 
0.0 -0.5704 0 2.0 1e-06 
0.0 -0.5703 0 2.0 1e-06 
0.0 -0.5702 0 2.0 1e-06 
0.0 -0.5701 0 2.0 1e-06 
0.0 -0.57 0 2.0 1e-06 
0.0 -0.5699 0 2.0 1e-06 
0.0 -0.5698 0 2.0 1e-06 
0.0 -0.5697 0 2.0 1e-06 
0.0 -0.5696 0 2.0 1e-06 
0.0 -0.5695 0 2.0 1e-06 
0.0 -0.5694 0 2.0 1e-06 
0.0 -0.5693 0 2.0 1e-06 
0.0 -0.5692 0 2.0 1e-06 
0.0 -0.5691 0 2.0 1e-06 
0.0 -0.569 0 2.0 1e-06 
0.0 -0.5689 0 2.0 1e-06 
0.0 -0.5688 0 2.0 1e-06 
0.0 -0.5687 0 2.0 1e-06 
0.0 -0.5686 0 2.0 1e-06 
0.0 -0.5685 0 2.0 1e-06 
0.0 -0.5684 0 2.0 1e-06 
0.0 -0.5683 0 2.0 1e-06 
0.0 -0.5682 0 2.0 1e-06 
0.0 -0.5681 0 2.0 1e-06 
0.0 -0.568 0 2.0 1e-06 
0.0 -0.5679 0 2.0 1e-06 
0.0 -0.5678 0 2.0 1e-06 
0.0 -0.5677 0 2.0 1e-06 
0.0 -0.5676 0 2.0 1e-06 
0.0 -0.5675 0 2.0 1e-06 
0.0 -0.5674 0 2.0 1e-06 
0.0 -0.5673 0 2.0 1e-06 
0.0 -0.5672 0 2.0 1e-06 
0.0 -0.5671 0 2.0 1e-06 
0.0 -0.567 0 2.0 1e-06 
0.0 -0.5669 0 2.0 1e-06 
0.0 -0.5668 0 2.0 1e-06 
0.0 -0.5667 0 2.0 1e-06 
0.0 -0.5666 0 2.0 1e-06 
0.0 -0.5665 0 2.0 1e-06 
0.0 -0.5664 0 2.0 1e-06 
0.0 -0.5663 0 2.0 1e-06 
0.0 -0.5662 0 2.0 1e-06 
0.0 -0.5661 0 2.0 1e-06 
0.0 -0.566 0 2.0 1e-06 
0.0 -0.5659 0 2.0 1e-06 
0.0 -0.5658 0 2.0 1e-06 
0.0 -0.5657 0 2.0 1e-06 
0.0 -0.5656 0 2.0 1e-06 
0.0 -0.5655 0 2.0 1e-06 
0.0 -0.5654 0 2.0 1e-06 
0.0 -0.5653 0 2.0 1e-06 
0.0 -0.5652 0 2.0 1e-06 
0.0 -0.5651 0 2.0 1e-06 
0.0 -0.565 0 2.0 1e-06 
0.0 -0.5649 0 2.0 1e-06 
0.0 -0.5648 0 2.0 1e-06 
0.0 -0.5647 0 2.0 1e-06 
0.0 -0.5646 0 2.0 1e-06 
0.0 -0.5645 0 2.0 1e-06 
0.0 -0.5644 0 2.0 1e-06 
0.0 -0.5643 0 2.0 1e-06 
0.0 -0.5642 0 2.0 1e-06 
0.0 -0.5641 0 2.0 1e-06 
0.0 -0.564 0 2.0 1e-06 
0.0 -0.5639 0 2.0 1e-06 
0.0 -0.5638 0 2.0 1e-06 
0.0 -0.5637 0 2.0 1e-06 
0.0 -0.5636 0 2.0 1e-06 
0.0 -0.5635 0 2.0 1e-06 
0.0 -0.5634 0 2.0 1e-06 
0.0 -0.5633 0 2.0 1e-06 
0.0 -0.5632 0 2.0 1e-06 
0.0 -0.5631 0 2.0 1e-06 
0.0 -0.563 0 2.0 1e-06 
0.0 -0.5629 0 2.0 1e-06 
0.0 -0.5628 0 2.0 1e-06 
0.0 -0.5627 0 2.0 1e-06 
0.0 -0.5626 0 2.0 1e-06 
0.0 -0.5625 0 2.0 1e-06 
0.0 -0.5624 0 2.0 1e-06 
0.0 -0.5623 0 2.0 1e-06 
0.0 -0.5622 0 2.0 1e-06 
0.0 -0.5621 0 2.0 1e-06 
0.0 -0.562 0 2.0 1e-06 
0.0 -0.5619 0 2.0 1e-06 
0.0 -0.5618 0 2.0 1e-06 
0.0 -0.5617 0 2.0 1e-06 
0.0 -0.5616 0 2.0 1e-06 
0.0 -0.5615 0 2.0 1e-06 
0.0 -0.5614 0 2.0 1e-06 
0.0 -0.5613 0 2.0 1e-06 
0.0 -0.5612 0 2.0 1e-06 
0.0 -0.5611 0 2.0 1e-06 
0.0 -0.561 0 2.0 1e-06 
0.0 -0.5609 0 2.0 1e-06 
0.0 -0.5608 0 2.0 1e-06 
0.0 -0.5607 0 2.0 1e-06 
0.0 -0.5606 0 2.0 1e-06 
0.0 -0.5605 0 2.0 1e-06 
0.0 -0.5604 0 2.0 1e-06 
0.0 -0.5603 0 2.0 1e-06 
0.0 -0.5602 0 2.0 1e-06 
0.0 -0.5601 0 2.0 1e-06 
0.0 -0.56 0 2.0 1e-06 
0.0 -0.5599 0 2.0 1e-06 
0.0 -0.5598 0 2.0 1e-06 
0.0 -0.5597 0 2.0 1e-06 
0.0 -0.5596 0 2.0 1e-06 
0.0 -0.5595 0 2.0 1e-06 
0.0 -0.5594 0 2.0 1e-06 
0.0 -0.5593 0 2.0 1e-06 
0.0 -0.5592 0 2.0 1e-06 
0.0 -0.5591 0 2.0 1e-06 
0.0 -0.559 0 2.0 1e-06 
0.0 -0.5589 0 2.0 1e-06 
0.0 -0.5588 0 2.0 1e-06 
0.0 -0.5587 0 2.0 1e-06 
0.0 -0.5586 0 2.0 1e-06 
0.0 -0.5585 0 2.0 1e-06 
0.0 -0.5584 0 2.0 1e-06 
0.0 -0.5583 0 2.0 1e-06 
0.0 -0.5582 0 2.0 1e-06 
0.0 -0.5581 0 2.0 1e-06 
0.0 -0.558 0 2.0 1e-06 
0.0 -0.5579 0 2.0 1e-06 
0.0 -0.5578 0 2.0 1e-06 
0.0 -0.5577 0 2.0 1e-06 
0.0 -0.5576 0 2.0 1e-06 
0.0 -0.5575 0 2.0 1e-06 
0.0 -0.5574 0 2.0 1e-06 
0.0 -0.5573 0 2.0 1e-06 
0.0 -0.5572 0 2.0 1e-06 
0.0 -0.5571 0 2.0 1e-06 
0.0 -0.557 0 2.0 1e-06 
0.0 -0.5569 0 2.0 1e-06 
0.0 -0.5568 0 2.0 1e-06 
0.0 -0.5567 0 2.0 1e-06 
0.0 -0.5566 0 2.0 1e-06 
0.0 -0.5565 0 2.0 1e-06 
0.0 -0.5564 0 2.0 1e-06 
0.0 -0.5563 0 2.0 1e-06 
0.0 -0.5562 0 2.0 1e-06 
0.0 -0.5561 0 2.0 1e-06 
0.0 -0.556 0 2.0 1e-06 
0.0 -0.5559 0 2.0 1e-06 
0.0 -0.5558 0 2.0 1e-06 
0.0 -0.5557 0 2.0 1e-06 
0.0 -0.5556 0 2.0 1e-06 
0.0 -0.5555 0 2.0 1e-06 
0.0 -0.5554 0 2.0 1e-06 
0.0 -0.5553 0 2.0 1e-06 
0.0 -0.5552 0 2.0 1e-06 
0.0 -0.5551 0 2.0 1e-06 
0.0 -0.555 0 2.0 1e-06 
0.0 -0.5549 0 2.0 1e-06 
0.0 -0.5548 0 2.0 1e-06 
0.0 -0.5547 0 2.0 1e-06 
0.0 -0.5546 0 2.0 1e-06 
0.0 -0.5545 0 2.0 1e-06 
0.0 -0.5544 0 2.0 1e-06 
0.0 -0.5543 0 2.0 1e-06 
0.0 -0.5542 0 2.0 1e-06 
0.0 -0.5541 0 2.0 1e-06 
0.0 -0.554 0 2.0 1e-06 
0.0 -0.5539 0 2.0 1e-06 
0.0 -0.5538 0 2.0 1e-06 
0.0 -0.5537 0 2.0 1e-06 
0.0 -0.5536 0 2.0 1e-06 
0.0 -0.5535 0 2.0 1e-06 
0.0 -0.5534 0 2.0 1e-06 
0.0 -0.5533 0 2.0 1e-06 
0.0 -0.5532 0 2.0 1e-06 
0.0 -0.5531 0 2.0 1e-06 
0.0 -0.553 0 2.0 1e-06 
0.0 -0.5529 0 2.0 1e-06 
0.0 -0.5528 0 2.0 1e-06 
0.0 -0.5527 0 2.0 1e-06 
0.0 -0.5526 0 2.0 1e-06 
0.0 -0.5525 0 2.0 1e-06 
0.0 -0.5524 0 2.0 1e-06 
0.0 -0.5523 0 2.0 1e-06 
0.0 -0.5522 0 2.0 1e-06 
0.0 -0.5521 0 2.0 1e-06 
0.0 -0.552 0 2.0 1e-06 
0.0 -0.5519 0 2.0 1e-06 
0.0 -0.5518 0 2.0 1e-06 
0.0 -0.5517 0 2.0 1e-06 
0.0 -0.5516 0 2.0 1e-06 
0.0 -0.5515 0 2.0 1e-06 
0.0 -0.5514 0 2.0 1e-06 
0.0 -0.5513 0 2.0 1e-06 
0.0 -0.5512 0 2.0 1e-06 
0.0 -0.5511 0 2.0 1e-06 
0.0 -0.551 0 2.0 1e-06 
0.0 -0.5509 0 2.0 1e-06 
0.0 -0.5508 0 2.0 1e-06 
0.0 -0.5507 0 2.0 1e-06 
0.0 -0.5506 0 2.0 1e-06 
0.0 -0.5505 0 2.0 1e-06 
0.0 -0.5504 0 2.0 1e-06 
0.0 -0.5503 0 2.0 1e-06 
0.0 -0.5502 0 2.0 1e-06 
0.0 -0.5501 0 2.0 1e-06 
0.0 -0.55 0 2.0 1e-06 
0.0 -0.5499 0 2.0 1e-06 
0.0 -0.5498 0 2.0 1e-06 
0.0 -0.5497 0 2.0 1e-06 
0.0 -0.5496 0 2.0 1e-06 
0.0 -0.5495 0 2.0 1e-06 
0.0 -0.5494 0 2.0 1e-06 
0.0 -0.5493 0 2.0 1e-06 
0.0 -0.5492 0 2.0 1e-06 
0.0 -0.5491 0 2.0 1e-06 
0.0 -0.549 0 2.0 1e-06 
0.0 -0.5489 0 2.0 1e-06 
0.0 -0.5488 0 2.0 1e-06 
0.0 -0.5487 0 2.0 1e-06 
0.0 -0.5486 0 2.0 1e-06 
0.0 -0.5485 0 2.0 1e-06 
0.0 -0.5484 0 2.0 1e-06 
0.0 -0.5483 0 2.0 1e-06 
0.0 -0.5482 0 2.0 1e-06 
0.0 -0.5481 0 2.0 1e-06 
0.0 -0.548 0 2.0 1e-06 
0.0 -0.5479 0 2.0 1e-06 
0.0 -0.5478 0 2.0 1e-06 
0.0 -0.5477 0 2.0 1e-06 
0.0 -0.5476 0 2.0 1e-06 
0.0 -0.5475 0 2.0 1e-06 
0.0 -0.5474 0 2.0 1e-06 
0.0 -0.5473 0 2.0 1e-06 
0.0 -0.5472 0 2.0 1e-06 
0.0 -0.5471 0 2.0 1e-06 
0.0 -0.547 0 2.0 1e-06 
0.0 -0.5469 0 2.0 1e-06 
0.0 -0.5468 0 2.0 1e-06 
0.0 -0.5467 0 2.0 1e-06 
0.0 -0.5466 0 2.0 1e-06 
0.0 -0.5465 0 2.0 1e-06 
0.0 -0.5464 0 2.0 1e-06 
0.0 -0.5463 0 2.0 1e-06 
0.0 -0.5462 0 2.0 1e-06 
0.0 -0.5461 0 2.0 1e-06 
0.0 -0.546 0 2.0 1e-06 
0.0 -0.5459 0 2.0 1e-06 
0.0 -0.5458 0 2.0 1e-06 
0.0 -0.5457 0 2.0 1e-06 
0.0 -0.5456 0 2.0 1e-06 
0.0 -0.5455 0 2.0 1e-06 
0.0 -0.5454 0 2.0 1e-06 
0.0 -0.5453 0 2.0 1e-06 
0.0 -0.5452 0 2.0 1e-06 
0.0 -0.5451 0 2.0 1e-06 
0.0 -0.545 0 2.0 1e-06 
0.0 -0.5449 0 2.0 1e-06 
0.0 -0.5448 0 2.0 1e-06 
0.0 -0.5447 0 2.0 1e-06 
0.0 -0.5446 0 2.0 1e-06 
0.0 -0.5445 0 2.0 1e-06 
0.0 -0.5444 0 2.0 1e-06 
0.0 -0.5443 0 2.0 1e-06 
0.0 -0.5442 0 2.0 1e-06 
0.0 -0.5441 0 2.0 1e-06 
0.0 -0.544 0 2.0 1e-06 
0.0 -0.5439 0 2.0 1e-06 
0.0 -0.5438 0 2.0 1e-06 
0.0 -0.5437 0 2.0 1e-06 
0.0 -0.5436 0 2.0 1e-06 
0.0 -0.5435 0 2.0 1e-06 
0.0 -0.5434 0 2.0 1e-06 
0.0 -0.5433 0 2.0 1e-06 
0.0 -0.5432 0 2.0 1e-06 
0.0 -0.5431 0 2.0 1e-06 
0.0 -0.543 0 2.0 1e-06 
0.0 -0.5429 0 2.0 1e-06 
0.0 -0.5428 0 2.0 1e-06 
0.0 -0.5427 0 2.0 1e-06 
0.0 -0.5426 0 2.0 1e-06 
0.0 -0.5425 0 2.0 1e-06 
0.0 -0.5424 0 2.0 1e-06 
0.0 -0.5423 0 2.0 1e-06 
0.0 -0.5422 0 2.0 1e-06 
0.0 -0.5421 0 2.0 1e-06 
0.0 -0.542 0 2.0 1e-06 
0.0 -0.5419 0 2.0 1e-06 
0.0 -0.5418 0 2.0 1e-06 
0.0 -0.5417 0 2.0 1e-06 
0.0 -0.5416 0 2.0 1e-06 
0.0 -0.5415 0 2.0 1e-06 
0.0 -0.5414 0 2.0 1e-06 
0.0 -0.5413 0 2.0 1e-06 
0.0 -0.5412 0 2.0 1e-06 
0.0 -0.5411 0 2.0 1e-06 
0.0 -0.541 0 2.0 1e-06 
0.0 -0.5409 0 2.0 1e-06 
0.0 -0.5408 0 2.0 1e-06 
0.0 -0.5407 0 2.0 1e-06 
0.0 -0.5406 0 2.0 1e-06 
0.0 -0.5405 0 2.0 1e-06 
0.0 -0.5404 0 2.0 1e-06 
0.0 -0.5403 0 2.0 1e-06 
0.0 -0.5402 0 2.0 1e-06 
0.0 -0.5401 0 2.0 1e-06 
0.0 -0.54 0 2.0 1e-06 
0.0 -0.5399 0 2.0 1e-06 
0.0 -0.5398 0 2.0 1e-06 
0.0 -0.5397 0 2.0 1e-06 
0.0 -0.5396 0 2.0 1e-06 
0.0 -0.5395 0 2.0 1e-06 
0.0 -0.5394 0 2.0 1e-06 
0.0 -0.5393 0 2.0 1e-06 
0.0 -0.5392 0 2.0 1e-06 
0.0 -0.5391 0 2.0 1e-06 
0.0 -0.539 0 2.0 1e-06 
0.0 -0.5389 0 2.0 1e-06 
0.0 -0.5388 0 2.0 1e-06 
0.0 -0.5387 0 2.0 1e-06 
0.0 -0.5386 0 2.0 1e-06 
0.0 -0.5385 0 2.0 1e-06 
0.0 -0.5384 0 2.0 1e-06 
0.0 -0.5383 0 2.0 1e-06 
0.0 -0.5382 0 2.0 1e-06 
0.0 -0.5381 0 2.0 1e-06 
0.0 -0.538 0 2.0 1e-06 
0.0 -0.5379 0 2.0 1e-06 
0.0 -0.5378 0 2.0 1e-06 
0.0 -0.5377 0 2.0 1e-06 
0.0 -0.5376 0 2.0 1e-06 
0.0 -0.5375 0 2.0 1e-06 
0.0 -0.5374 0 2.0 1e-06 
0.0 -0.5373 0 2.0 1e-06 
0.0 -0.5372 0 2.0 1e-06 
0.0 -0.5371 0 2.0 1e-06 
0.0 -0.537 0 2.0 1e-06 
0.0 -0.5369 0 2.0 1e-06 
0.0 -0.5368 0 2.0 1e-06 
0.0 -0.5367 0 2.0 1e-06 
0.0 -0.5366 0 2.0 1e-06 
0.0 -0.5365 0 2.0 1e-06 
0.0 -0.5364 0 2.0 1e-06 
0.0 -0.5363 0 2.0 1e-06 
0.0 -0.5362 0 2.0 1e-06 
0.0 -0.5361 0 2.0 1e-06 
0.0 -0.536 0 2.0 1e-06 
0.0 -0.5359 0 2.0 1e-06 
0.0 -0.5358 0 2.0 1e-06 
0.0 -0.5357 0 2.0 1e-06 
0.0 -0.5356 0 2.0 1e-06 
0.0 -0.5355 0 2.0 1e-06 
0.0 -0.5354 0 2.0 1e-06 
0.0 -0.5353 0 2.0 1e-06 
0.0 -0.5352 0 2.0 1e-06 
0.0 -0.5351 0 2.0 1e-06 
0.0 -0.535 0 2.0 1e-06 
0.0 -0.5349 0 2.0 1e-06 
0.0 -0.5348 0 2.0 1e-06 
0.0 -0.5347 0 2.0 1e-06 
0.0 -0.5346 0 2.0 1e-06 
0.0 -0.5345 0 2.0 1e-06 
0.0 -0.5344 0 2.0 1e-06 
0.0 -0.5343 0 2.0 1e-06 
0.0 -0.5342 0 2.0 1e-06 
0.0 -0.5341 0 2.0 1e-06 
0.0 -0.534 0 2.0 1e-06 
0.0 -0.5339 0 2.0 1e-06 
0.0 -0.5338 0 2.0 1e-06 
0.0 -0.5337 0 2.0 1e-06 
0.0 -0.5336 0 2.0 1e-06 
0.0 -0.5335 0 2.0 1e-06 
0.0 -0.5334 0 2.0 1e-06 
0.0 -0.5333 0 2.0 1e-06 
0.0 -0.5332 0 2.0 1e-06 
0.0 -0.5331 0 2.0 1e-06 
0.0 -0.533 0 2.0 1e-06 
0.0 -0.5329 0 2.0 1e-06 
0.0 -0.5328 0 2.0 1e-06 
0.0 -0.5327 0 2.0 1e-06 
0.0 -0.5326 0 2.0 1e-06 
0.0 -0.5325 0 2.0 1e-06 
0.0 -0.5324 0 2.0 1e-06 
0.0 -0.5323 0 2.0 1e-06 
0.0 -0.5322 0 2.0 1e-06 
0.0 -0.5321 0 2.0 1e-06 
0.0 -0.532 0 2.0 1e-06 
0.0 -0.5319 0 2.0 1e-06 
0.0 -0.5318 0 2.0 1e-06 
0.0 -0.5317 0 2.0 1e-06 
0.0 -0.5316 0 2.0 1e-06 
0.0 -0.5315 0 2.0 1e-06 
0.0 -0.5314 0 2.0 1e-06 
0.0 -0.5313 0 2.0 1e-06 
0.0 -0.5312 0 2.0 1e-06 
0.0 -0.5311 0 2.0 1e-06 
0.0 -0.531 0 2.0 1e-06 
0.0 -0.5309 0 2.0 1e-06 
0.0 -0.5308 0 2.0 1e-06 
0.0 -0.5307 0 2.0 1e-06 
0.0 -0.5306 0 2.0 1e-06 
0.0 -0.5305 0 2.0 1e-06 
0.0 -0.5304 0 2.0 1e-06 
0.0 -0.5303 0 2.0 1e-06 
0.0 -0.5302 0 2.0 1e-06 
0.0 -0.5301 0 2.0 1e-06 
0.0 -0.53 0 2.0 1e-06 
0.0 -0.5299 0 2.0 1e-06 
0.0 -0.5298 0 2.0 1e-06 
0.0 -0.5297 0 2.0 1e-06 
0.0 -0.5296 0 2.0 1e-06 
0.0 -0.5295 0 2.0 1e-06 
0.0 -0.5294 0 2.0 1e-06 
0.0 -0.5293 0 2.0 1e-06 
0.0 -0.5292 0 2.0 1e-06 
0.0 -0.5291 0 2.0 1e-06 
0.0 -0.529 0 2.0 1e-06 
0.0 -0.5289 0 2.0 1e-06 
0.0 -0.5288 0 2.0 1e-06 
0.0 -0.5287 0 2.0 1e-06 
0.0 -0.5286 0 2.0 1e-06 
0.0 -0.5285 0 2.0 1e-06 
0.0 -0.5284 0 2.0 1e-06 
0.0 -0.5283 0 2.0 1e-06 
0.0 -0.5282 0 2.0 1e-06 
0.0 -0.5281 0 2.0 1e-06 
0.0 -0.528 0 2.0 1e-06 
0.0 -0.5279 0 2.0 1e-06 
0.0 -0.5278 0 2.0 1e-06 
0.0 -0.5277 0 2.0 1e-06 
0.0 -0.5276 0 2.0 1e-06 
0.0 -0.5275 0 2.0 1e-06 
0.0 -0.5274 0 2.0 1e-06 
0.0 -0.5273 0 2.0 1e-06 
0.0 -0.5272 0 2.0 1e-06 
0.0 -0.5271 0 2.0 1e-06 
0.0 -0.527 0 2.0 1e-06 
0.0 -0.5269 0 2.0 1e-06 
0.0 -0.5268 0 2.0 1e-06 
0.0 -0.5267 0 2.0 1e-06 
0.0 -0.5266 0 2.0 1e-06 
0.0 -0.5265 0 2.0 1e-06 
0.0 -0.5264 0 2.0 1e-06 
0.0 -0.5263 0 2.0 1e-06 
0.0 -0.5262 0 2.0 1e-06 
0.0 -0.5261 0 2.0 1e-06 
0.0 -0.526 0 2.0 1e-06 
0.0 -0.5259 0 2.0 1e-06 
0.0 -0.5258 0 2.0 1e-06 
0.0 -0.5257 0 2.0 1e-06 
0.0 -0.5256 0 2.0 1e-06 
0.0 -0.5255 0 2.0 1e-06 
0.0 -0.5254 0 2.0 1e-06 
0.0 -0.5253 0 2.0 1e-06 
0.0 -0.5252 0 2.0 1e-06 
0.0 -0.5251 0 2.0 1e-06 
0.0 -0.525 0 2.0 1e-06 
0.0 -0.5249 0 2.0 1e-06 
0.0 -0.5248 0 2.0 1e-06 
0.0 -0.5247 0 2.0 1e-06 
0.0 -0.5246 0 2.0 1e-06 
0.0 -0.5245 0 2.0 1e-06 
0.0 -0.5244 0 2.0 1e-06 
0.0 -0.5243 0 2.0 1e-06 
0.0 -0.5242 0 2.0 1e-06 
0.0 -0.5241 0 2.0 1e-06 
0.0 -0.524 0 2.0 1e-06 
0.0 -0.5239 0 2.0 1e-06 
0.0 -0.5238 0 2.0 1e-06 
0.0 -0.5237 0 2.0 1e-06 
0.0 -0.5236 0 2.0 1e-06 
0.0 -0.5235 0 2.0 1e-06 
0.0 -0.5234 0 2.0 1e-06 
0.0 -0.5233 0 2.0 1e-06 
0.0 -0.5232 0 2.0 1e-06 
0.0 -0.5231 0 2.0 1e-06 
0.0 -0.523 0 2.0 1e-06 
0.0 -0.5229 0 2.0 1e-06 
0.0 -0.5228 0 2.0 1e-06 
0.0 -0.5227 0 2.0 1e-06 
0.0 -0.5226 0 2.0 1e-06 
0.0 -0.5225 0 2.0 1e-06 
0.0 -0.5224 0 2.0 1e-06 
0.0 -0.5223 0 2.0 1e-06 
0.0 -0.5222 0 2.0 1e-06 
0.0 -0.5221 0 2.0 1e-06 
0.0 -0.522 0 2.0 1e-06 
0.0 -0.5219 0 2.0 1e-06 
0.0 -0.5218 0 2.0 1e-06 
0.0 -0.5217 0 2.0 1e-06 
0.0 -0.5216 0 2.0 1e-06 
0.0 -0.5215 0 2.0 1e-06 
0.0 -0.5214 0 2.0 1e-06 
0.0 -0.5213 0 2.0 1e-06 
0.0 -0.5212 0 2.0 1e-06 
0.0 -0.5211 0 2.0 1e-06 
0.0 -0.521 0 2.0 1e-06 
0.0 -0.5209 0 2.0 1e-06 
0.0 -0.5208 0 2.0 1e-06 
0.0 -0.5207 0 2.0 1e-06 
0.0 -0.5206 0 2.0 1e-06 
0.0 -0.5205 0 2.0 1e-06 
0.0 -0.5204 0 2.0 1e-06 
0.0 -0.5203 0 2.0 1e-06 
0.0 -0.5202 0 2.0 1e-06 
0.0 -0.5201 0 2.0 1e-06 
0.0 -0.52 0 2.0 1e-06 
0.0 -0.5199 0 2.0 1e-06 
0.0 -0.5198 0 2.0 1e-06 
0.0 -0.5197 0 2.0 1e-06 
0.0 -0.5196 0 2.0 1e-06 
0.0 -0.5195 0 2.0 1e-06 
0.0 -0.5194 0 2.0 1e-06 
0.0 -0.5193 0 2.0 1e-06 
0.0 -0.5192 0 2.0 1e-06 
0.0 -0.5191 0 2.0 1e-06 
0.0 -0.519 0 2.0 1e-06 
0.0 -0.5189 0 2.0 1e-06 
0.0 -0.5188 0 2.0 1e-06 
0.0 -0.5187 0 2.0 1e-06 
0.0 -0.5186 0 2.0 1e-06 
0.0 -0.5185 0 2.0 1e-06 
0.0 -0.5184 0 2.0 1e-06 
0.0 -0.5183 0 2.0 1e-06 
0.0 -0.5182 0 2.0 1e-06 
0.0 -0.5181 0 2.0 1e-06 
0.0 -0.518 0 2.0 1e-06 
0.0 -0.5179 0 2.0 1e-06 
0.0 -0.5178 0 2.0 1e-06 
0.0 -0.5177 0 2.0 1e-06 
0.0 -0.5176 0 2.0 1e-06 
0.0 -0.5175 0 2.0 1e-06 
0.0 -0.5174 0 2.0 1e-06 
0.0 -0.5173 0 2.0 1e-06 
0.0 -0.5172 0 2.0 1e-06 
0.0 -0.5171 0 2.0 1e-06 
0.0 -0.517 0 2.0 1e-06 
0.0 -0.5169 0 2.0 1e-06 
0.0 -0.5168 0 2.0 1e-06 
0.0 -0.5167 0 2.0 1e-06 
0.0 -0.5166 0 2.0 1e-06 
0.0 -0.5165 0 2.0 1e-06 
0.0 -0.5164 0 2.0 1e-06 
0.0 -0.5163 0 2.0 1e-06 
0.0 -0.5162 0 2.0 1e-06 
0.0 -0.5161 0 2.0 1e-06 
0.0 -0.516 0 2.0 1e-06 
0.0 -0.5159 0 2.0 1e-06 
0.0 -0.5158 0 2.0 1e-06 
0.0 -0.5157 0 2.0 1e-06 
0.0 -0.5156 0 2.0 1e-06 
0.0 -0.5155 0 2.0 1e-06 
0.0 -0.5154 0 2.0 1e-06 
0.0 -0.5153 0 2.0 1e-06 
0.0 -0.5152 0 2.0 1e-06 
0.0 -0.5151 0 2.0 1e-06 
0.0 -0.515 0 2.0 1e-06 
0.0 -0.5149 0 2.0 1e-06 
0.0 -0.5148 0 2.0 1e-06 
0.0 -0.5147 0 2.0 1e-06 
0.0 -0.5146 0 2.0 1e-06 
0.0 -0.5145 0 2.0 1e-06 
0.0 -0.5144 0 2.0 1e-06 
0.0 -0.5143 0 2.0 1e-06 
0.0 -0.5142 0 2.0 1e-06 
0.0 -0.5141 0 2.0 1e-06 
0.0 -0.514 0 2.0 1e-06 
0.0 -0.5139 0 2.0 1e-06 
0.0 -0.5138 0 2.0 1e-06 
0.0 -0.5137 0 2.0 1e-06 
0.0 -0.5136 0 2.0 1e-06 
0.0 -0.5135 0 2.0 1e-06 
0.0 -0.5134 0 2.0 1e-06 
0.0 -0.5133 0 2.0 1e-06 
0.0 -0.5132 0 2.0 1e-06 
0.0 -0.5131 0 2.0 1e-06 
0.0 -0.513 0 2.0 1e-06 
0.0 -0.5129 0 2.0 1e-06 
0.0 -0.5128 0 2.0 1e-06 
0.0 -0.5127 0 2.0 1e-06 
0.0 -0.5126 0 2.0 1e-06 
0.0 -0.5125 0 2.0 1e-06 
0.0 -0.5124 0 2.0 1e-06 
0.0 -0.5123 0 2.0 1e-06 
0.0 -0.5122 0 2.0 1e-06 
0.0 -0.5121 0 2.0 1e-06 
0.0 -0.512 0 2.0 1e-06 
0.0 -0.5119 0 2.0 1e-06 
0.0 -0.5118 0 2.0 1e-06 
0.0 -0.5117 0 2.0 1e-06 
0.0 -0.5116 0 2.0 1e-06 
0.0 -0.5115 0 2.0 1e-06 
0.0 -0.5114 0 2.0 1e-06 
0.0 -0.5113 0 2.0 1e-06 
0.0 -0.5112 0 2.0 1e-06 
0.0 -0.5111 0 2.0 1e-06 
0.0 -0.511 0 2.0 1e-06 
0.0 -0.5109 0 2.0 1e-06 
0.0 -0.5108 0 2.0 1e-06 
0.0 -0.5107 0 2.0 1e-06 
0.0 -0.5106 0 2.0 1e-06 
0.0 -0.5105 0 2.0 1e-06 
0.0 -0.5104 0 2.0 1e-06 
0.0 -0.5103 0 2.0 1e-06 
0.0 -0.5102 0 2.0 1e-06 
0.0 -0.5101 0 2.0 1e-06 
0.0 -0.51 0 2.0 1e-06 
0.0 -0.5099 0 2.0 1e-06 
0.0 -0.5098 0 2.0 1e-06 
0.0 -0.5097 0 2.0 1e-06 
0.0 -0.5096 0 2.0 1e-06 
0.0 -0.5095 0 2.0 1e-06 
0.0 -0.5094 0 2.0 1e-06 
0.0 -0.5093 0 2.0 1e-06 
0.0 -0.5092 0 2.0 1e-06 
0.0 -0.5091 0 2.0 1e-06 
0.0 -0.509 0 2.0 1e-06 
0.0 -0.5089 0 2.0 1e-06 
0.0 -0.5088 0 2.0 1e-06 
0.0 -0.5087 0 2.0 1e-06 
0.0 -0.5086 0 2.0 1e-06 
0.0 -0.5085 0 2.0 1e-06 
0.0 -0.5084 0 2.0 1e-06 
0.0 -0.5083 0 2.0 1e-06 
0.0 -0.5082 0 2.0 1e-06 
0.0 -0.5081 0 2.0 1e-06 
0.0 -0.508 0 2.0 1e-06 
0.0 -0.5079 0 2.0 1e-06 
0.0 -0.5078 0 2.0 1e-06 
0.0 -0.5077 0 2.0 1e-06 
0.0 -0.5076 0 2.0 1e-06 
0.0 -0.5075 0 2.0 1e-06 
0.0 -0.5074 0 2.0 1e-06 
0.0 -0.5073 0 2.0 1e-06 
0.0 -0.5072 0 2.0 1e-06 
0.0 -0.5071 0 2.0 1e-06 
0.0 -0.507 0 2.0 1e-06 
0.0 -0.5069 0 2.0 1e-06 
0.0 -0.5068 0 2.0 1e-06 
0.0 -0.5067 0 2.0 1e-06 
0.0 -0.5066 0 2.0 1e-06 
0.0 -0.5065 0 2.0 1e-06 
0.0 -0.5064 0 2.0 1e-06 
0.0 -0.5063 0 2.0 1e-06 
0.0 -0.5062 0 2.0 1e-06 
0.0 -0.5061 0 2.0 1e-06 
0.0 -0.506 0 2.0 1e-06 
0.0 -0.5059 0 2.0 1e-06 
0.0 -0.5058 0 2.0 1e-06 
0.0 -0.5057 0 2.0 1e-06 
0.0 -0.5056 0 2.0 1e-06 
0.0 -0.5055 0 2.0 1e-06 
0.0 -0.5054 0 2.0 1e-06 
0.0 -0.5053 0 2.0 1e-06 
0.0 -0.5052 0 2.0 1e-06 
0.0 -0.5051 0 2.0 1e-06 
0.0 -0.505 0 2.0 1e-06 
0.0 -0.5049 0 2.0 1e-06 
0.0 -0.5048 0 2.0 1e-06 
0.0 -0.5047 0 2.0 1e-06 
0.0 -0.5046 0 2.0 1e-06 
0.0 -0.5045 0 2.0 1e-06 
0.0 -0.5044 0 2.0 1e-06 
0.0 -0.5043 0 2.0 1e-06 
0.0 -0.5042 0 2.0 1e-06 
0.0 -0.5041 0 2.0 1e-06 
0.0 -0.504 0 2.0 1e-06 
0.0 -0.5039 0 2.0 1e-06 
0.0 -0.5038 0 2.0 1e-06 
0.0 -0.5037 0 2.0 1e-06 
0.0 -0.5036 0 2.0 1e-06 
0.0 -0.5035 0 2.0 1e-06 
0.0 -0.5034 0 2.0 1e-06 
0.0 -0.5033 0 2.0 1e-06 
0.0 -0.5032 0 2.0 1e-06 
0.0 -0.5031 0 2.0 1e-06 
0.0 -0.503 0 2.0 1e-06 
0.0 -0.5029 0 2.0 1e-06 
0.0 -0.5028 0 2.0 1e-06 
0.0 -0.5027 0 2.0 1e-06 
0.0 -0.5026 0 2.0 1e-06 
0.0 -0.5025 0 2.0 1e-06 
0.0 -0.5024 0 2.0 1e-06 
0.0 -0.5023 0 2.0 1e-06 
0.0 -0.5022 0 2.0 1e-06 
0.0 -0.5021 0 2.0 1e-06 
0.0 -0.502 0 2.0 1e-06 
0.0 -0.5019 0 2.0 1e-06 
0.0 -0.5018 0 2.0 1e-06 
0.0 -0.5017 0 2.0 1e-06 
0.0 -0.5016 0 2.0 1e-06 
0.0 -0.5015 0 2.0 1e-06 
0.0 -0.5014 0 2.0 1e-06 
0.0 -0.5013 0 2.0 1e-06 
0.0 -0.5012 0 2.0 1e-06 
0.0 -0.5011 0 2.0 1e-06 
0.0 -0.501 0 2.0 1e-06 
0.0 -0.5009 0 2.0 1e-06 
0.0 -0.5008 0 2.0 1e-06 
0.0 -0.5007 0 2.0 1e-06 
0.0 -0.5006 0 2.0 1e-06 
0.0 -0.5005 0 2.0 1e-06 
0.0 -0.5004 0 2.0 1e-06 
0.0 -0.5003 0 2.0 1e-06 
0.0 -0.5002 0 2.0 1e-06 
0.0 -0.5001 0 2.0 1e-06 
0.0 -0.5 0 2.0 1e-06 
0.0 -0.4999 0 2.0 1e-06 
0.0 -0.4998 0 2.0 1e-06 
0.0 -0.4997 0 2.0 1e-06 
0.0 -0.4996 0 2.0 1e-06 
0.0 -0.4995 0 2.0 1e-06 
0.0 -0.4994 0 2.0 1e-06 
0.0 -0.4993 0 2.0 1e-06 
0.0 -0.4992 0 2.0 1e-06 
0.0 -0.4991 0 2.0 1e-06 
0.0 -0.499 0 2.0 1e-06 
0.0 -0.4989 0 2.0 1e-06 
0.0 -0.4988 0 2.0 1e-06 
0.0 -0.4987 0 2.0 1e-06 
0.0 -0.4986 0 2.0 1e-06 
0.0 -0.4985 0 2.0 1e-06 
0.0 -0.4984 0 2.0 1e-06 
0.0 -0.4983 0 2.0 1e-06 
0.0 -0.4982 0 2.0 1e-06 
0.0 -0.4981 0 2.0 1e-06 
0.0 -0.498 0 2.0 1e-06 
0.0 -0.4979 0 2.0 1e-06 
0.0 -0.4978 0 2.0 1e-06 
0.0 -0.4977 0 2.0 1e-06 
0.0 -0.4976 0 2.0 1e-06 
0.0 -0.4975 0 2.0 1e-06 
0.0 -0.4974 0 2.0 1e-06 
0.0 -0.4973 0 2.0 1e-06 
0.0 -0.4972 0 2.0 1e-06 
0.0 -0.4971 0 2.0 1e-06 
0.0 -0.497 0 2.0 1e-06 
0.0 -0.4969 0 2.0 1e-06 
0.0 -0.4968 0 2.0 1e-06 
0.0 -0.4967 0 2.0 1e-06 
0.0 -0.4966 0 2.0 1e-06 
0.0 -0.4965 0 2.0 1e-06 
0.0 -0.4964 0 2.0 1e-06 
0.0 -0.4963 0 2.0 1e-06 
0.0 -0.4962 0 2.0 1e-06 
0.0 -0.4961 0 2.0 1e-06 
0.0 -0.496 0 2.0 1e-06 
0.0 -0.4959 0 2.0 1e-06 
0.0 -0.4958 0 2.0 1e-06 
0.0 -0.4957 0 2.0 1e-06 
0.0 -0.4956 0 2.0 1e-06 
0.0 -0.4955 0 2.0 1e-06 
0.0 -0.4954 0 2.0 1e-06 
0.0 -0.4953 0 2.0 1e-06 
0.0 -0.4952 0 2.0 1e-06 
0.0 -0.4951 0 2.0 1e-06 
0.0 -0.495 0 2.0 1e-06 
0.0 -0.4949 0 2.0 1e-06 
0.0 -0.4948 0 2.0 1e-06 
0.0 -0.4947 0 2.0 1e-06 
0.0 -0.4946 0 2.0 1e-06 
0.0 -0.4945 0 2.0 1e-06 
0.0 -0.4944 0 2.0 1e-06 
0.0 -0.4943 0 2.0 1e-06 
0.0 -0.4942 0 2.0 1e-06 
0.0 -0.4941 0 2.0 1e-06 
0.0 -0.494 0 2.0 1e-06 
0.0 -0.4939 0 2.0 1e-06 
0.0 -0.4938 0 2.0 1e-06 
0.0 -0.4937 0 2.0 1e-06 
0.0 -0.4936 0 2.0 1e-06 
0.0 -0.4935 0 2.0 1e-06 
0.0 -0.4934 0 2.0 1e-06 
0.0 -0.4933 0 2.0 1e-06 
0.0 -0.4932 0 2.0 1e-06 
0.0 -0.4931 0 2.0 1e-06 
0.0 -0.493 0 2.0 1e-06 
0.0 -0.4929 0 2.0 1e-06 
0.0 -0.4928 0 2.0 1e-06 
0.0 -0.4927 0 2.0 1e-06 
0.0 -0.4926 0 2.0 1e-06 
0.0 -0.4925 0 2.0 1e-06 
0.0 -0.4924 0 2.0 1e-06 
0.0 -0.4923 0 2.0 1e-06 
0.0 -0.4922 0 2.0 1e-06 
0.0 -0.4921 0 2.0 1e-06 
0.0 -0.492 0 2.0 1e-06 
0.0 -0.4919 0 2.0 1e-06 
0.0 -0.4918 0 2.0 1e-06 
0.0 -0.4917 0 2.0 1e-06 
0.0 -0.4916 0 2.0 1e-06 
0.0 -0.4915 0 2.0 1e-06 
0.0 -0.4914 0 2.0 1e-06 
0.0 -0.4913 0 2.0 1e-06 
0.0 -0.4912 0 2.0 1e-06 
0.0 -0.4911 0 2.0 1e-06 
0.0 -0.491 0 2.0 1e-06 
0.0 -0.4909 0 2.0 1e-06 
0.0 -0.4908 0 2.0 1e-06 
0.0 -0.4907 0 2.0 1e-06 
0.0 -0.4906 0 2.0 1e-06 
0.0 -0.4905 0 2.0 1e-06 
0.0 -0.4904 0 2.0 1e-06 
0.0 -0.4903 0 2.0 1e-06 
0.0 -0.4902 0 2.0 1e-06 
0.0 -0.4901 0 2.0 1e-06 
0.0 -0.49 0 2.0 1e-06 
0.0 -0.4899 0 2.0 1e-06 
0.0 -0.4898 0 2.0 1e-06 
0.0 -0.4897 0 2.0 1e-06 
0.0 -0.4896 0 2.0 1e-06 
0.0 -0.4895 0 2.0 1e-06 
0.0 -0.4894 0 2.0 1e-06 
0.0 -0.4893 0 2.0 1e-06 
0.0 -0.4892 0 2.0 1e-06 
0.0 -0.4891 0 2.0 1e-06 
0.0 -0.489 0 2.0 1e-06 
0.0 -0.4889 0 2.0 1e-06 
0.0 -0.4888 0 2.0 1e-06 
0.0 -0.4887 0 2.0 1e-06 
0.0 -0.4886 0 2.0 1e-06 
0.0 -0.4885 0 2.0 1e-06 
0.0 -0.4884 0 2.0 1e-06 
0.0 -0.4883 0 2.0 1e-06 
0.0 -0.4882 0 2.0 1e-06 
0.0 -0.4881 0 2.0 1e-06 
0.0 -0.488 0 2.0 1e-06 
0.0 -0.4879 0 2.0 1e-06 
0.0 -0.4878 0 2.0 1e-06 
0.0 -0.4877 0 2.0 1e-06 
0.0 -0.4876 0 2.0 1e-06 
0.0 -0.4875 0 2.0 1e-06 
0.0 -0.4874 0 2.0 1e-06 
0.0 -0.4873 0 2.0 1e-06 
0.0 -0.4872 0 2.0 1e-06 
0.0 -0.4871 0 2.0 1e-06 
0.0 -0.487 0 2.0 1e-06 
0.0 -0.4869 0 2.0 1e-06 
0.0 -0.4868 0 2.0 1e-06 
0.0 -0.4867 0 2.0 1e-06 
0.0 -0.4866 0 2.0 1e-06 
0.0 -0.4865 0 2.0 1e-06 
0.0 -0.4864 0 2.0 1e-06 
0.0 -0.4863 0 2.0 1e-06 
0.0 -0.4862 0 2.0 1e-06 
0.0 -0.4861 0 2.0 1e-06 
0.0 -0.486 0 2.0 1e-06 
0.0 -0.4859 0 2.0 1e-06 
0.0 -0.4858 0 2.0 1e-06 
0.0 -0.4857 0 2.0 1e-06 
0.0 -0.4856 0 2.0 1e-06 
0.0 -0.4855 0 2.0 1e-06 
0.0 -0.4854 0 2.0 1e-06 
0.0 -0.4853 0 2.0 1e-06 
0.0 -0.4852 0 2.0 1e-06 
0.0 -0.4851 0 2.0 1e-06 
0.0 -0.485 0 2.0 1e-06 
0.0 -0.4849 0 2.0 1e-06 
0.0 -0.4848 0 2.0 1e-06 
0.0 -0.4847 0 2.0 1e-06 
0.0 -0.4846 0 2.0 1e-06 
0.0 -0.4845 0 2.0 1e-06 
0.0 -0.4844 0 2.0 1e-06 
0.0 -0.4843 0 2.0 1e-06 
0.0 -0.4842 0 2.0 1e-06 
0.0 -0.4841 0 2.0 1e-06 
0.0 -0.484 0 2.0 1e-06 
0.0 -0.4839 0 2.0 1e-06 
0.0 -0.4838 0 2.0 1e-06 
0.0 -0.4837 0 2.0 1e-06 
0.0 -0.4836 0 2.0 1e-06 
0.0 -0.4835 0 2.0 1e-06 
0.0 -0.4834 0 2.0 1e-06 
0.0 -0.4833 0 2.0 1e-06 
0.0 -0.4832 0 2.0 1e-06 
0.0 -0.4831 0 2.0 1e-06 
0.0 -0.483 0 2.0 1e-06 
0.0 -0.4829 0 2.0 1e-06 
0.0 -0.4828 0 2.0 1e-06 
0.0 -0.4827 0 2.0 1e-06 
0.0 -0.4826 0 2.0 1e-06 
0.0 -0.4825 0 2.0 1e-06 
0.0 -0.4824 0 2.0 1e-06 
0.0 -0.4823 0 2.0 1e-06 
0.0 -0.4822 0 2.0 1e-06 
0.0 -0.4821 0 2.0 1e-06 
0.0 -0.482 0 2.0 1e-06 
0.0 -0.4819 0 2.0 1e-06 
0.0 -0.4818 0 2.0 1e-06 
0.0 -0.4817 0 2.0 1e-06 
0.0 -0.4816 0 2.0 1e-06 
0.0 -0.4815 0 2.0 1e-06 
0.0 -0.4814 0 2.0 1e-06 
0.0 -0.4813 0 2.0 1e-06 
0.0 -0.4812 0 2.0 1e-06 
0.0 -0.4811 0 2.0 1e-06 
0.0 -0.481 0 2.0 1e-06 
0.0 -0.4809 0 2.0 1e-06 
0.0 -0.4808 0 2.0 1e-06 
0.0 -0.4807 0 2.0 1e-06 
0.0 -0.4806 0 2.0 1e-06 
0.0 -0.4805 0 2.0 1e-06 
0.0 -0.4804 0 2.0 1e-06 
0.0 -0.4803 0 2.0 1e-06 
0.0 -0.4802 0 2.0 1e-06 
0.0 -0.4801 0 2.0 1e-06 
0.0 -0.48 0 2.0 1e-06 
0.0 -0.4799 0 2.0 1e-06 
0.0 -0.4798 0 2.0 1e-06 
0.0 -0.4797 0 2.0 1e-06 
0.0 -0.4796 0 2.0 1e-06 
0.0 -0.4795 0 2.0 1e-06 
0.0 -0.4794 0 2.0 1e-06 
0.0 -0.4793 0 2.0 1e-06 
0.0 -0.4792 0 2.0 1e-06 
0.0 -0.4791 0 2.0 1e-06 
0.0 -0.479 0 2.0 1e-06 
0.0 -0.4789 0 2.0 1e-06 
0.0 -0.4788 0 2.0 1e-06 
0.0 -0.4787 0 2.0 1e-06 
0.0 -0.4786 0 2.0 1e-06 
0.0 -0.4785 0 2.0 1e-06 
0.0 -0.4784 0 2.0 1e-06 
0.0 -0.4783 0 2.0 1e-06 
0.0 -0.4782 0 2.0 1e-06 
0.0 -0.4781 0 2.0 1e-06 
0.0 -0.478 0 2.0 1e-06 
0.0 -0.4779 0 2.0 1e-06 
0.0 -0.4778 0 2.0 1e-06 
0.0 -0.4777 0 2.0 1e-06 
0.0 -0.4776 0 2.0 1e-06 
0.0 -0.4775 0 2.0 1e-06 
0.0 -0.4774 0 2.0 1e-06 
0.0 -0.4773 0 2.0 1e-06 
0.0 -0.4772 0 2.0 1e-06 
0.0 -0.4771 0 2.0 1e-06 
0.0 -0.477 0 2.0 1e-06 
0.0 -0.4769 0 2.0 1e-06 
0.0 -0.4768 0 2.0 1e-06 
0.0 -0.4767 0 2.0 1e-06 
0.0 -0.4766 0 2.0 1e-06 
0.0 -0.4765 0 2.0 1e-06 
0.0 -0.4764 0 2.0 1e-06 
0.0 -0.4763 0 2.0 1e-06 
0.0 -0.4762 0 2.0 1e-06 
0.0 -0.4761 0 2.0 1e-06 
0.0 -0.476 0 2.0 1e-06 
0.0 -0.4759 0 2.0 1e-06 
0.0 -0.4758 0 2.0 1e-06 
0.0 -0.4757 0 2.0 1e-06 
0.0 -0.4756 0 2.0 1e-06 
0.0 -0.4755 0 2.0 1e-06 
0.0 -0.4754 0 2.0 1e-06 
0.0 -0.4753 0 2.0 1e-06 
0.0 -0.4752 0 2.0 1e-06 
0.0 -0.4751 0 2.0 1e-06 
0.0 -0.475 0 2.0 1e-06 
0.0 -0.4749 0 2.0 1e-06 
0.0 -0.4748 0 2.0 1e-06 
0.0 -0.4747 0 2.0 1e-06 
0.0 -0.4746 0 2.0 1e-06 
0.0 -0.4745 0 2.0 1e-06 
0.0 -0.4744 0 2.0 1e-06 
0.0 -0.4743 0 2.0 1e-06 
0.0 -0.4742 0 2.0 1e-06 
0.0 -0.4741 0 2.0 1e-06 
0.0 -0.474 0 2.0 1e-06 
0.0 -0.4739 0 2.0 1e-06 
0.0 -0.4738 0 2.0 1e-06 
0.0 -0.4737 0 2.0 1e-06 
0.0 -0.4736 0 2.0 1e-06 
0.0 -0.4735 0 2.0 1e-06 
0.0 -0.4734 0 2.0 1e-06 
0.0 -0.4733 0 2.0 1e-06 
0.0 -0.4732 0 2.0 1e-06 
0.0 -0.4731 0 2.0 1e-06 
0.0 -0.473 0 2.0 1e-06 
0.0 -0.4729 0 2.0 1e-06 
0.0 -0.4728 0 2.0 1e-06 
0.0 -0.4727 0 2.0 1e-06 
0.0 -0.4726 0 2.0 1e-06 
0.0 -0.4725 0 2.0 1e-06 
0.0 -0.4724 0 2.0 1e-06 
0.0 -0.4723 0 2.0 1e-06 
0.0 -0.4722 0 2.0 1e-06 
0.0 -0.4721 0 2.0 1e-06 
0.0 -0.472 0 2.0 1e-06 
0.0 -0.4719 0 2.0 1e-06 
0.0 -0.4718 0 2.0 1e-06 
0.0 -0.4717 0 2.0 1e-06 
0.0 -0.4716 0 2.0 1e-06 
0.0 -0.4715 0 2.0 1e-06 
0.0 -0.4714 0 2.0 1e-06 
0.0 -0.4713 0 2.0 1e-06 
0.0 -0.4712 0 2.0 1e-06 
0.0 -0.4711 0 2.0 1e-06 
0.0 -0.471 0 2.0 1e-06 
0.0 -0.4709 0 2.0 1e-06 
0.0 -0.4708 0 2.0 1e-06 
0.0 -0.4707 0 2.0 1e-06 
0.0 -0.4706 0 2.0 1e-06 
0.0 -0.4705 0 2.0 1e-06 
0.0 -0.4704 0 2.0 1e-06 
0.0 -0.4703 0 2.0 1e-06 
0.0 -0.4702 0 2.0 1e-06 
0.0 -0.4701 0 2.0 1e-06 
0.0 -0.47 0 2.0 1e-06 
0.0 -0.4699 0 2.0 1e-06 
0.0 -0.4698 0 2.0 1e-06 
0.0 -0.4697 0 2.0 1e-06 
0.0 -0.4696 0 2.0 1e-06 
0.0 -0.4695 0 2.0 1e-06 
0.0 -0.4694 0 2.0 1e-06 
0.0 -0.4693 0 2.0 1e-06 
0.0 -0.4692 0 2.0 1e-06 
0.0 -0.4691 0 2.0 1e-06 
0.0 -0.469 0 2.0 1e-06 
0.0 -0.4689 0 2.0 1e-06 
0.0 -0.4688 0 2.0 1e-06 
0.0 -0.4687 0 2.0 1e-06 
0.0 -0.4686 0 2.0 1e-06 
0.0 -0.4685 0 2.0 1e-06 
0.0 -0.4684 0 2.0 1e-06 
0.0 -0.4683 0 2.0 1e-06 
0.0 -0.4682 0 2.0 1e-06 
0.0 -0.4681 0 2.0 1e-06 
0.0 -0.468 0 2.0 1e-06 
0.0 -0.4679 0 2.0 1e-06 
0.0 -0.4678 0 2.0 1e-06 
0.0 -0.4677 0 2.0 1e-06 
0.0 -0.4676 0 2.0 1e-06 
0.0 -0.4675 0 2.0 1e-06 
0.0 -0.4674 0 2.0 1e-06 
0.0 -0.4673 0 2.0 1e-06 
0.0 -0.4672 0 2.0 1e-06 
0.0 -0.4671 0 2.0 1e-06 
0.0 -0.467 0 2.0 1e-06 
0.0 -0.4669 0 2.0 1e-06 
0.0 -0.4668 0 2.0 1e-06 
0.0 -0.4667 0 2.0 1e-06 
0.0 -0.4666 0 2.0 1e-06 
0.0 -0.4665 0 2.0 1e-06 
0.0 -0.4664 0 2.0 1e-06 
0.0 -0.4663 0 2.0 1e-06 
0.0 -0.4662 0 2.0 1e-06 
0.0 -0.4661 0 2.0 1e-06 
0.0 -0.466 0 2.0 1e-06 
0.0 -0.4659 0 2.0 1e-06 
0.0 -0.4658 0 2.0 1e-06 
0.0 -0.4657 0 2.0 1e-06 
0.0 -0.4656 0 2.0 1e-06 
0.0 -0.4655 0 2.0 1e-06 
0.0 -0.4654 0 2.0 1e-06 
0.0 -0.4653 0 2.0 1e-06 
0.0 -0.4652 0 2.0 1e-06 
0.0 -0.4651 0 2.0 1e-06 
0.0 -0.465 0 2.0 1e-06 
0.0 -0.4649 0 2.0 1e-06 
0.0 -0.4648 0 2.0 1e-06 
0.0 -0.4647 0 2.0 1e-06 
0.0 -0.4646 0 2.0 1e-06 
0.0 -0.4645 0 2.0 1e-06 
0.0 -0.4644 0 2.0 1e-06 
0.0 -0.4643 0 2.0 1e-06 
0.0 -0.4642 0 2.0 1e-06 
0.0 -0.4641 0 2.0 1e-06 
0.0 -0.464 0 2.0 1e-06 
0.0 -0.4639 0 2.0 1e-06 
0.0 -0.4638 0 2.0 1e-06 
0.0 -0.4637 0 2.0 1e-06 
0.0 -0.4636 0 2.0 1e-06 
0.0 -0.4635 0 2.0 1e-06 
0.0 -0.4634 0 2.0 1e-06 
0.0 -0.4633 0 2.0 1e-06 
0.0 -0.4632 0 2.0 1e-06 
0.0 -0.4631 0 2.0 1e-06 
0.0 -0.463 0 2.0 1e-06 
0.0 -0.4629 0 2.0 1e-06 
0.0 -0.4628 0 2.0 1e-06 
0.0 -0.4627 0 2.0 1e-06 
0.0 -0.4626 0 2.0 1e-06 
0.0 -0.4625 0 2.0 1e-06 
0.0 -0.4624 0 2.0 1e-06 
0.0 -0.4623 0 2.0 1e-06 
0.0 -0.4622 0 2.0 1e-06 
0.0 -0.4621 0 2.0 1e-06 
0.0 -0.462 0 2.0 1e-06 
0.0 -0.4619 0 2.0 1e-06 
0.0 -0.4618 0 2.0 1e-06 
0.0 -0.4617 0 2.0 1e-06 
0.0 -0.4616 0 2.0 1e-06 
0.0 -0.4615 0 2.0 1e-06 
0.0 -0.4614 0 2.0 1e-06 
0.0 -0.4613 0 2.0 1e-06 
0.0 -0.4612 0 2.0 1e-06 
0.0 -0.4611 0 2.0 1e-06 
0.0 -0.461 0 2.0 1e-06 
0.0 -0.4609 0 2.0 1e-06 
0.0 -0.4608 0 2.0 1e-06 
0.0 -0.4607 0 2.0 1e-06 
0.0 -0.4606 0 2.0 1e-06 
0.0 -0.4605 0 2.0 1e-06 
0.0 -0.4604 0 2.0 1e-06 
0.0 -0.4603 0 2.0 1e-06 
0.0 -0.4602 0 2.0 1e-06 
0.0 -0.4601 0 2.0 1e-06 
0.0 -0.46 0 2.0 1e-06 
0.0 -0.4599 0 2.0 1e-06 
0.0 -0.4598 0 2.0 1e-06 
0.0 -0.4597 0 2.0 1e-06 
0.0 -0.4596 0 2.0 1e-06 
0.0 -0.4595 0 2.0 1e-06 
0.0 -0.4594 0 2.0 1e-06 
0.0 -0.4593 0 2.0 1e-06 
0.0 -0.4592 0 2.0 1e-06 
0.0 -0.4591 0 2.0 1e-06 
0.0 -0.459 0 2.0 1e-06 
0.0 -0.4589 0 2.0 1e-06 
0.0 -0.4588 0 2.0 1e-06 
0.0 -0.4587 0 2.0 1e-06 
0.0 -0.4586 0 2.0 1e-06 
0.0 -0.4585 0 2.0 1e-06 
0.0 -0.4584 0 2.0 1e-06 
0.0 -0.4583 0 2.0 1e-06 
0.0 -0.4582 0 2.0 1e-06 
0.0 -0.4581 0 2.0 1e-06 
0.0 -0.458 0 2.0 1e-06 
0.0 -0.4579 0 2.0 1e-06 
0.0 -0.4578 0 2.0 1e-06 
0.0 -0.4577 0 2.0 1e-06 
0.0 -0.4576 0 2.0 1e-06 
0.0 -0.4575 0 2.0 1e-06 
0.0 -0.4574 0 2.0 1e-06 
0.0 -0.4573 0 2.0 1e-06 
0.0 -0.4572 0 2.0 1e-06 
0.0 -0.4571 0 2.0 1e-06 
0.0 -0.457 0 2.0 1e-06 
0.0 -0.4569 0 2.0 1e-06 
0.0 -0.4568 0 2.0 1e-06 
0.0 -0.4567 0 2.0 1e-06 
0.0 -0.4566 0 2.0 1e-06 
0.0 -0.4565 0 2.0 1e-06 
0.0 -0.4564 0 2.0 1e-06 
0.0 -0.4563 0 2.0 1e-06 
0.0 -0.4562 0 2.0 1e-06 
0.0 -0.4561 0 2.0 1e-06 
0.0 -0.456 0 2.0 1e-06 
0.0 -0.4559 0 2.0 1e-06 
0.0 -0.4558 0 2.0 1e-06 
0.0 -0.4557 0 2.0 1e-06 
0.0 -0.4556 0 2.0 1e-06 
0.0 -0.4555 0 2.0 1e-06 
0.0 -0.4554 0 2.0 1e-06 
0.0 -0.4553 0 2.0 1e-06 
0.0 -0.4552 0 2.0 1e-06 
0.0 -0.4551 0 2.0 1e-06 
0.0 -0.455 0 2.0 1e-06 
0.0 -0.4549 0 2.0 1e-06 
0.0 -0.4548 0 2.0 1e-06 
0.0 -0.4547 0 2.0 1e-06 
0.0 -0.4546 0 2.0 1e-06 
0.0 -0.4545 0 2.0 1e-06 
0.0 -0.4544 0 2.0 1e-06 
0.0 -0.4543 0 2.0 1e-06 
0.0 -0.4542 0 2.0 1e-06 
0.0 -0.4541 0 2.0 1e-06 
0.0 -0.454 0 2.0 1e-06 
0.0 -0.4539 0 2.0 1e-06 
0.0 -0.4538 0 2.0 1e-06 
0.0 -0.4537 0 2.0 1e-06 
0.0 -0.4536 0 2.0 1e-06 
0.0 -0.4535 0 2.0 1e-06 
0.0 -0.4534 0 2.0 1e-06 
0.0 -0.4533 0 2.0 1e-06 
0.0 -0.4532 0 2.0 1e-06 
0.0 -0.4531 0 2.0 1e-06 
0.0 -0.453 0 2.0 1e-06 
0.0 -0.4529 0 2.0 1e-06 
0.0 -0.4528 0 2.0 1e-06 
0.0 -0.4527 0 2.0 1e-06 
0.0 -0.4526 0 2.0 1e-06 
0.0 -0.4525 0 2.0 1e-06 
0.0 -0.4524 0 2.0 1e-06 
0.0 -0.4523 0 2.0 1e-06 
0.0 -0.4522 0 2.0 1e-06 
0.0 -0.4521 0 2.0 1e-06 
0.0 -0.452 0 2.0 1e-06 
0.0 -0.4519 0 2.0 1e-06 
0.0 -0.4518 0 2.0 1e-06 
0.0 -0.4517 0 2.0 1e-06 
0.0 -0.4516 0 2.0 1e-06 
0.0 -0.4515 0 2.0 1e-06 
0.0 -0.4514 0 2.0 1e-06 
0.0 -0.4513 0 2.0 1e-06 
0.0 -0.4512 0 2.0 1e-06 
0.0 -0.4511 0 2.0 1e-06 
0.0 -0.451 0 2.0 1e-06 
0.0 -0.4509 0 2.0 1e-06 
0.0 -0.4508 0 2.0 1e-06 
0.0 -0.4507 0 2.0 1e-06 
0.0 -0.4506 0 2.0 1e-06 
0.0 -0.4505 0 2.0 1e-06 
0.0 -0.4504 0 2.0 1e-06 
0.0 -0.4503 0 2.0 1e-06 
0.0 -0.4502 0 2.0 1e-06 
0.0 -0.4501 0 2.0 1e-06 
0.0 -0.45 0 2.0 1e-06 
0.0 -0.4499 0 2.0 1e-06 
0.0 -0.4498 0 2.0 1e-06 
0.0 -0.4497 0 2.0 1e-06 
0.0 -0.4496 0 2.0 1e-06 
0.0 -0.4495 0 2.0 1e-06 
0.0 -0.4494 0 2.0 1e-06 
0.0 -0.4493 0 2.0 1e-06 
0.0 -0.4492 0 2.0 1e-06 
0.0 -0.4491 0 2.0 1e-06 
0.0 -0.449 0 2.0 1e-06 
0.0 -0.4489 0 2.0 1e-06 
0.0 -0.4488 0 2.0 1e-06 
0.0 -0.4487 0 2.0 1e-06 
0.0 -0.4486 0 2.0 1e-06 
0.0 -0.4485 0 2.0 1e-06 
0.0 -0.4484 0 2.0 1e-06 
0.0 -0.4483 0 2.0 1e-06 
0.0 -0.4482 0 2.0 1e-06 
0.0 -0.4481 0 2.0 1e-06 
0.0 -0.448 0 2.0 1e-06 
0.0 -0.4479 0 2.0 1e-06 
0.0 -0.4478 0 2.0 1e-06 
0.0 -0.4477 0 2.0 1e-06 
0.0 -0.4476 0 2.0 1e-06 
0.0 -0.4475 0 2.0 1e-06 
0.0 -0.4474 0 2.0 1e-06 
0.0 -0.4473 0 2.0 1e-06 
0.0 -0.4472 0 2.0 1e-06 
0.0 -0.4471 0 2.0 1e-06 
0.0 -0.447 0 2.0 1e-06 
0.0 -0.4469 0 2.0 1e-06 
0.0 -0.4468 0 2.0 1e-06 
0.0 -0.4467 0 2.0 1e-06 
0.0 -0.4466 0 2.0 1e-06 
0.0 -0.4465 0 2.0 1e-06 
0.0 -0.4464 0 2.0 1e-06 
0.0 -0.4463 0 2.0 1e-06 
0.0 -0.4462 0 2.0 1e-06 
0.0 -0.4461 0 2.0 1e-06 
0.0 -0.446 0 2.0 1e-06 
0.0 -0.4459 0 2.0 1e-06 
0.0 -0.4458 0 2.0 1e-06 
0.0 -0.4457 0 2.0 1e-06 
0.0 -0.4456 0 2.0 1e-06 
0.0 -0.4455 0 2.0 1e-06 
0.0 -0.4454 0 2.0 1e-06 
0.0 -0.4453 0 2.0 1e-06 
0.0 -0.4452 0 2.0 1e-06 
0.0 -0.4451 0 2.0 1e-06 
0.0 -0.445 0 2.0 1e-06 
0.0 -0.4449 0 2.0 1e-06 
0.0 -0.4448 0 2.0 1e-06 
0.0 -0.4447 0 2.0 1e-06 
0.0 -0.4446 0 2.0 1e-06 
0.0 -0.4445 0 2.0 1e-06 
0.0 -0.4444 0 2.0 1e-06 
0.0 -0.4443 0 2.0 1e-06 
0.0 -0.4442 0 2.0 1e-06 
0.0 -0.4441 0 2.0 1e-06 
0.0 -0.444 0 2.0 1e-06 
0.0 -0.4439 0 2.0 1e-06 
0.0 -0.4438 0 2.0 1e-06 
0.0 -0.4437 0 2.0 1e-06 
0.0 -0.4436 0 2.0 1e-06 
0.0 -0.4435 0 2.0 1e-06 
0.0 -0.4434 0 2.0 1e-06 
0.0 -0.4433 0 2.0 1e-06 
0.0 -0.4432 0 2.0 1e-06 
0.0 -0.4431 0 2.0 1e-06 
0.0 -0.443 0 2.0 1e-06 
0.0 -0.4429 0 2.0 1e-06 
0.0 -0.4428 0 2.0 1e-06 
0.0 -0.4427 0 2.0 1e-06 
0.0 -0.4426 0 2.0 1e-06 
0.0 -0.4425 0 2.0 1e-06 
0.0 -0.4424 0 2.0 1e-06 
0.0 -0.4423 0 2.0 1e-06 
0.0 -0.4422 0 2.0 1e-06 
0.0 -0.4421 0 2.0 1e-06 
0.0 -0.442 0 2.0 1e-06 
0.0 -0.4419 0 2.0 1e-06 
0.0 -0.4418 0 2.0 1e-06 
0.0 -0.4417 0 2.0 1e-06 
0.0 -0.4416 0 2.0 1e-06 
0.0 -0.4415 0 2.0 1e-06 
0.0 -0.4414 0 2.0 1e-06 
0.0 -0.4413 0 2.0 1e-06 
0.0 -0.4412 0 2.0 1e-06 
0.0 -0.4411 0 2.0 1e-06 
0.0 -0.441 0 2.0 1e-06 
0.0 -0.4409 0 2.0 1e-06 
0.0 -0.4408 0 2.0 1e-06 
0.0 -0.4407 0 2.0 1e-06 
0.0 -0.4406 0 2.0 1e-06 
0.0 -0.4405 0 2.0 1e-06 
0.0 -0.4404 0 2.0 1e-06 
0.0 -0.4403 0 2.0 1e-06 
0.0 -0.4402 0 2.0 1e-06 
0.0 -0.4401 0 2.0 1e-06 
0.0 -0.44 0 2.0 1e-06 
0.0 -0.4399 0 2.0 1e-06 
0.0 -0.4398 0 2.0 1e-06 
0.0 -0.4397 0 2.0 1e-06 
0.0 -0.4396 0 2.0 1e-06 
0.0 -0.4395 0 2.0 1e-06 
0.0 -0.4394 0 2.0 1e-06 
0.0 -0.4393 0 2.0 1e-06 
0.0 -0.4392 0 2.0 1e-06 
0.0 -0.4391 0 2.0 1e-06 
0.0 -0.439 0 2.0 1e-06 
0.0 -0.4389 0 2.0 1e-06 
0.0 -0.4388 0 2.0 1e-06 
0.0 -0.4387 0 2.0 1e-06 
0.0 -0.4386 0 2.0 1e-06 
0.0 -0.4385 0 2.0 1e-06 
0.0 -0.4384 0 2.0 1e-06 
0.0 -0.4383 0 2.0 1e-06 
0.0 -0.4382 0 2.0 1e-06 
0.0 -0.4381 0 2.0 1e-06 
0.0 -0.438 0 2.0 1e-06 
0.0 -0.4379 0 2.0 1e-06 
0.0 -0.4378 0 2.0 1e-06 
0.0 -0.4377 0 2.0 1e-06 
0.0 -0.4376 0 2.0 1e-06 
0.0 -0.4375 0 2.0 1e-06 
0.0 -0.4374 0 2.0 1e-06 
0.0 -0.4373 0 2.0 1e-06 
0.0 -0.4372 0 2.0 1e-06 
0.0 -0.4371 0 2.0 1e-06 
0.0 -0.437 0 2.0 1e-06 
0.0 -0.4369 0 2.0 1e-06 
0.0 -0.4368 0 2.0 1e-06 
0.0 -0.4367 0 2.0 1e-06 
0.0 -0.4366 0 2.0 1e-06 
0.0 -0.4365 0 2.0 1e-06 
0.0 -0.4364 0 2.0 1e-06 
0.0 -0.4363 0 2.0 1e-06 
0.0 -0.4362 0 2.0 1e-06 
0.0 -0.4361 0 2.0 1e-06 
0.0 -0.436 0 2.0 1e-06 
0.0 -0.4359 0 2.0 1e-06 
0.0 -0.4358 0 2.0 1e-06 
0.0 -0.4357 0 2.0 1e-06 
0.0 -0.4356 0 2.0 1e-06 
0.0 -0.4355 0 2.0 1e-06 
0.0 -0.4354 0 2.0 1e-06 
0.0 -0.4353 0 2.0 1e-06 
0.0 -0.4352 0 2.0 1e-06 
0.0 -0.4351 0 2.0 1e-06 
0.0 -0.435 0 2.0 1e-06 
0.0 -0.4349 0 2.0 1e-06 
0.0 -0.4348 0 2.0 1e-06 
0.0 -0.4347 0 2.0 1e-06 
0.0 -0.4346 0 2.0 1e-06 
0.0 -0.4345 0 2.0 1e-06 
0.0 -0.4344 0 2.0 1e-06 
0.0 -0.4343 0 2.0 1e-06 
0.0 -0.4342 0 2.0 1e-06 
0.0 -0.4341 0 2.0 1e-06 
0.0 -0.434 0 2.0 1e-06 
0.0 -0.4339 0 2.0 1e-06 
0.0 -0.4338 0 2.0 1e-06 
0.0 -0.4337 0 2.0 1e-06 
0.0 -0.4336 0 2.0 1e-06 
0.0 -0.4335 0 2.0 1e-06 
0.0 -0.4334 0 2.0 1e-06 
0.0 -0.4333 0 2.0 1e-06 
0.0 -0.4332 0 2.0 1e-06 
0.0 -0.4331 0 2.0 1e-06 
0.0 -0.433 0 2.0 1e-06 
0.0 -0.4329 0 2.0 1e-06 
0.0 -0.4328 0 2.0 1e-06 
0.0 -0.4327 0 2.0 1e-06 
0.0 -0.4326 0 2.0 1e-06 
0.0 -0.4325 0 2.0 1e-06 
0.0 -0.4324 0 2.0 1e-06 
0.0 -0.4323 0 2.0 1e-06 
0.0 -0.4322 0 2.0 1e-06 
0.0 -0.4321 0 2.0 1e-06 
0.0 -0.432 0 2.0 1e-06 
0.0 -0.4319 0 2.0 1e-06 
0.0 -0.4318 0 2.0 1e-06 
0.0 -0.4317 0 2.0 1e-06 
0.0 -0.4316 0 2.0 1e-06 
0.0 -0.4315 0 2.0 1e-06 
0.0 -0.4314 0 2.0 1e-06 
0.0 -0.4313 0 2.0 1e-06 
0.0 -0.4312 0 2.0 1e-06 
0.0 -0.4311 0 2.0 1e-06 
0.0 -0.431 0 2.0 1e-06 
0.0 -0.4309 0 2.0 1e-06 
0.0 -0.4308 0 2.0 1e-06 
0.0 -0.4307 0 2.0 1e-06 
0.0 -0.4306 0 2.0 1e-06 
0.0 -0.4305 0 2.0 1e-06 
0.0 -0.4304 0 2.0 1e-06 
0.0 -0.4303 0 2.0 1e-06 
0.0 -0.4302 0 2.0 1e-06 
0.0 -0.4301 0 2.0 1e-06 
0.0 -0.43 0 2.0 1e-06 
0.0 -0.4299 0 2.0 1e-06 
0.0 -0.4298 0 2.0 1e-06 
0.0 -0.4297 0 2.0 1e-06 
0.0 -0.4296 0 2.0 1e-06 
0.0 -0.4295 0 2.0 1e-06 
0.0 -0.4294 0 2.0 1e-06 
0.0 -0.4293 0 2.0 1e-06 
0.0 -0.4292 0 2.0 1e-06 
0.0 -0.4291 0 2.0 1e-06 
0.0 -0.429 0 2.0 1e-06 
0.0 -0.4289 0 2.0 1e-06 
0.0 -0.4288 0 2.0 1e-06 
0.0 -0.4287 0 2.0 1e-06 
0.0 -0.4286 0 2.0 1e-06 
0.0 -0.4285 0 2.0 1e-06 
0.0 -0.4284 0 2.0 1e-06 
0.0 -0.4283 0 2.0 1e-06 
0.0 -0.4282 0 2.0 1e-06 
0.0 -0.4281 0 2.0 1e-06 
0.0 -0.428 0 2.0 1e-06 
0.0 -0.4279 0 2.0 1e-06 
0.0 -0.4278 0 2.0 1e-06 
0.0 -0.4277 0 2.0 1e-06 
0.0 -0.4276 0 2.0 1e-06 
0.0 -0.4275 0 2.0 1e-06 
0.0 -0.4274 0 2.0 1e-06 
0.0 -0.4273 0 2.0 1e-06 
0.0 -0.4272 0 2.0 1e-06 
0.0 -0.4271 0 2.0 1e-06 
0.0 -0.427 0 2.0 1e-06 
0.0 -0.4269 0 2.0 1e-06 
0.0 -0.4268 0 2.0 1e-06 
0.0 -0.4267 0 2.0 1e-06 
0.0 -0.4266 0 2.0 1e-06 
0.0 -0.4265 0 2.0 1e-06 
0.0 -0.4264 0 2.0 1e-06 
0.0 -0.4263 0 2.0 1e-06 
0.0 -0.4262 0 2.0 1e-06 
0.0 -0.4261 0 2.0 1e-06 
0.0 -0.426 0 2.0 1e-06 
0.0 -0.4259 0 2.0 1e-06 
0.0 -0.4258 0 2.0 1e-06 
0.0 -0.4257 0 2.0 1e-06 
0.0 -0.4256 0 2.0 1e-06 
0.0 -0.4255 0 2.0 1e-06 
0.0 -0.4254 0 2.0 1e-06 
0.0 -0.4253 0 2.0 1e-06 
0.0 -0.4252 0 2.0 1e-06 
0.0 -0.4251 0 2.0 1e-06 
0.0 -0.425 0 2.0 1e-06 
0.0 -0.4249 0 2.0 1e-06 
0.0 -0.4248 0 2.0 1e-06 
0.0 -0.4247 0 2.0 1e-06 
0.0 -0.4246 0 2.0 1e-06 
0.0 -0.4245 0 2.0 1e-06 
0.0 -0.4244 0 2.0 1e-06 
0.0 -0.4243 0 2.0 1e-06 
0.0 -0.4242 0 2.0 1e-06 
0.0 -0.4241 0 2.0 1e-06 
0.0 -0.424 0 2.0 1e-06 
0.0 -0.4239 0 2.0 1e-06 
0.0 -0.4238 0 2.0 1e-06 
0.0 -0.4237 0 2.0 1e-06 
0.0 -0.4236 0 2.0 1e-06 
0.0 -0.4235 0 2.0 1e-06 
0.0 -0.4234 0 2.0 1e-06 
0.0 -0.4233 0 2.0 1e-06 
0.0 -0.4232 0 2.0 1e-06 
0.0 -0.4231 0 2.0 1e-06 
0.0 -0.423 0 2.0 1e-06 
0.0 -0.4229 0 2.0 1e-06 
0.0 -0.4228 0 2.0 1e-06 
0.0 -0.4227 0 2.0 1e-06 
0.0 -0.4226 0 2.0 1e-06 
0.0 -0.4225 0 2.0 1e-06 
0.0 -0.4224 0 2.0 1e-06 
0.0 -0.4223 0 2.0 1e-06 
0.0 -0.4222 0 2.0 1e-06 
0.0 -0.4221 0 2.0 1e-06 
0.0 -0.422 0 2.0 1e-06 
0.0 -0.4219 0 2.0 1e-06 
0.0 -0.4218 0 2.0 1e-06 
0.0 -0.4217 0 2.0 1e-06 
0.0 -0.4216 0 2.0 1e-06 
0.0 -0.4215 0 2.0 1e-06 
0.0 -0.4214 0 2.0 1e-06 
0.0 -0.4213 0 2.0 1e-06 
0.0 -0.4212 0 2.0 1e-06 
0.0 -0.4211 0 2.0 1e-06 
0.0 -0.421 0 2.0 1e-06 
0.0 -0.4209 0 2.0 1e-06 
0.0 -0.4208 0 2.0 1e-06 
0.0 -0.4207 0 2.0 1e-06 
0.0 -0.4206 0 2.0 1e-06 
0.0 -0.4205 0 2.0 1e-06 
0.0 -0.4204 0 2.0 1e-06 
0.0 -0.4203 0 2.0 1e-06 
0.0 -0.4202 0 2.0 1e-06 
0.0 -0.4201 0 2.0 1e-06 
0.0 -0.42 0 2.0 1e-06 
0.0 -0.4199 0 2.0 1e-06 
0.0 -0.4198 0 2.0 1e-06 
0.0 -0.4197 0 2.0 1e-06 
0.0 -0.4196 0 2.0 1e-06 
0.0 -0.4195 0 2.0 1e-06 
0.0 -0.4194 0 2.0 1e-06 
0.0 -0.4193 0 2.0 1e-06 
0.0 -0.4192 0 2.0 1e-06 
0.0 -0.4191 0 2.0 1e-06 
0.0 -0.419 0 2.0 1e-06 
0.0 -0.4189 0 2.0 1e-06 
0.0 -0.4188 0 2.0 1e-06 
0.0 -0.4187 0 2.0 1e-06 
0.0 -0.4186 0 2.0 1e-06 
0.0 -0.4185 0 2.0 1e-06 
0.0 -0.4184 0 2.0 1e-06 
0.0 -0.4183 0 2.0 1e-06 
0.0 -0.4182 0 2.0 1e-06 
0.0 -0.4181 0 2.0 1e-06 
0.0 -0.418 0 2.0 1e-06 
0.0 -0.4179 0 2.0 1e-06 
0.0 -0.4178 0 2.0 1e-06 
0.0 -0.4177 0 2.0 1e-06 
0.0 -0.4176 0 2.0 1e-06 
0.0 -0.4175 0 2.0 1e-06 
0.0 -0.4174 0 2.0 1e-06 
0.0 -0.4173 0 2.0 1e-06 
0.0 -0.4172 0 2.0 1e-06 
0.0 -0.4171 0 2.0 1e-06 
0.0 -0.417 0 2.0 1e-06 
0.0 -0.4169 0 2.0 1e-06 
0.0 -0.4168 0 2.0 1e-06 
0.0 -0.4167 0 2.0 1e-06 
0.0 -0.4166 0 2.0 1e-06 
0.0 -0.4165 0 2.0 1e-06 
0.0 -0.4164 0 2.0 1e-06 
0.0 -0.4163 0 2.0 1e-06 
0.0 -0.4162 0 2.0 1e-06 
0.0 -0.4161 0 2.0 1e-06 
0.0 -0.416 0 2.0 1e-06 
0.0 -0.4159 0 2.0 1e-06 
0.0 -0.4158 0 2.0 1e-06 
0.0 -0.4157 0 2.0 1e-06 
0.0 -0.4156 0 2.0 1e-06 
0.0 -0.4155 0 2.0 1e-06 
0.0 -0.4154 0 2.0 1e-06 
0.0 -0.4153 0 2.0 1e-06 
0.0 -0.4152 0 2.0 1e-06 
0.0 -0.4151 0 2.0 1e-06 
0.0 -0.415 0 2.0 1e-06 
0.0 -0.4149 0 2.0 1e-06 
0.0 -0.4148 0 2.0 1e-06 
0.0 -0.4147 0 2.0 1e-06 
0.0 -0.4146 0 2.0 1e-06 
0.0 -0.4145 0 2.0 1e-06 
0.0 -0.4144 0 2.0 1e-06 
0.0 -0.4143 0 2.0 1e-06 
0.0 -0.4142 0 2.0 1e-06 
0.0 -0.4141 0 2.0 1e-06 
0.0 -0.414 0 2.0 1e-06 
0.0 -0.4139 0 2.0 1e-06 
0.0 -0.4138 0 2.0 1e-06 
0.0 -0.4137 0 2.0 1e-06 
0.0 -0.4136 0 2.0 1e-06 
0.0 -0.4135 0 2.0 1e-06 
0.0 -0.4134 0 2.0 1e-06 
0.0 -0.4133 0 2.0 1e-06 
0.0 -0.4132 0 2.0 1e-06 
0.0 -0.4131 0 2.0 1e-06 
0.0 -0.413 0 2.0 1e-06 
0.0 -0.4129 0 2.0 1e-06 
0.0 -0.4128 0 2.0 1e-06 
0.0 -0.4127 0 2.0 1e-06 
0.0 -0.4126 0 2.0 1e-06 
0.0 -0.4125 0 2.0 1e-06 
0.0 -0.4124 0 2.0 1e-06 
0.0 -0.4123 0 2.0 1e-06 
0.0 -0.4122 0 2.0 1e-06 
0.0 -0.4121 0 2.0 1e-06 
0.0 -0.412 0 2.0 1e-06 
0.0 -0.4119 0 2.0 1e-06 
0.0 -0.4118 0 2.0 1e-06 
0.0 -0.4117 0 2.0 1e-06 
0.0 -0.4116 0 2.0 1e-06 
0.0 -0.4115 0 2.0 1e-06 
0.0 -0.4114 0 2.0 1e-06 
0.0 -0.4113 0 2.0 1e-06 
0.0 -0.4112 0 2.0 1e-06 
0.0 -0.4111 0 2.0 1e-06 
0.0 -0.411 0 2.0 1e-06 
0.0 -0.4109 0 2.0 1e-06 
0.0 -0.4108 0 2.0 1e-06 
0.0 -0.4107 0 2.0 1e-06 
0.0 -0.4106 0 2.0 1e-06 
0.0 -0.4105 0 2.0 1e-06 
0.0 -0.4104 0 2.0 1e-06 
0.0 -0.4103 0 2.0 1e-06 
0.0 -0.4102 0 2.0 1e-06 
0.0 -0.4101 0 2.0 1e-06 
0.0 -0.41 0 2.0 1e-06 
0.0 -0.4099 0 2.0 1e-06 
0.0 -0.4098 0 2.0 1e-06 
0.0 -0.4097 0 2.0 1e-06 
0.0 -0.4096 0 2.0 1e-06 
0.0 -0.4095 0 2.0 1e-06 
0.0 -0.4094 0 2.0 1e-06 
0.0 -0.4093 0 2.0 1e-06 
0.0 -0.4092 0 2.0 1e-06 
0.0 -0.4091 0 2.0 1e-06 
0.0 -0.409 0 2.0 1e-06 
0.0 -0.4089 0 2.0 1e-06 
0.0 -0.4088 0 2.0 1e-06 
0.0 -0.4087 0 2.0 1e-06 
0.0 -0.4086 0 2.0 1e-06 
0.0 -0.4085 0 2.0 1e-06 
0.0 -0.4084 0 2.0 1e-06 
0.0 -0.4083 0 2.0 1e-06 
0.0 -0.4082 0 2.0 1e-06 
0.0 -0.4081 0 2.0 1e-06 
0.0 -0.408 0 2.0 1e-06 
0.0 -0.4079 0 2.0 1e-06 
0.0 -0.4078 0 2.0 1e-06 
0.0 -0.4077 0 2.0 1e-06 
0.0 -0.4076 0 2.0 1e-06 
0.0 -0.4075 0 2.0 1e-06 
0.0 -0.4074 0 2.0 1e-06 
0.0 -0.4073 0 2.0 1e-06 
0.0 -0.4072 0 2.0 1e-06 
0.0 -0.4071 0 2.0 1e-06 
0.0 -0.407 0 2.0 1e-06 
0.0 -0.4069 0 2.0 1e-06 
0.0 -0.4068 0 2.0 1e-06 
0.0 -0.4067 0 2.0 1e-06 
0.0 -0.4066 0 2.0 1e-06 
0.0 -0.4065 0 2.0 1e-06 
0.0 -0.4064 0 2.0 1e-06 
0.0 -0.4063 0 2.0 1e-06 
0.0 -0.4062 0 2.0 1e-06 
0.0 -0.4061 0 2.0 1e-06 
0.0 -0.406 0 2.0 1e-06 
0.0 -0.4059 0 2.0 1e-06 
0.0 -0.4058 0 2.0 1e-06 
0.0 -0.4057 0 2.0 1e-06 
0.0 -0.4056 0 2.0 1e-06 
0.0 -0.4055 0 2.0 1e-06 
0.0 -0.4054 0 2.0 1e-06 
0.0 -0.4053 0 2.0 1e-06 
0.0 -0.4052 0 2.0 1e-06 
0.0 -0.4051 0 2.0 1e-06 
0.0 -0.405 0 2.0 1e-06 
0.0 -0.4049 0 2.0 1e-06 
0.0 -0.4048 0 2.0 1e-06 
0.0 -0.4047 0 2.0 1e-06 
0.0 -0.4046 0 2.0 1e-06 
0.0 -0.4045 0 2.0 1e-06 
0.0 -0.4044 0 2.0 1e-06 
0.0 -0.4043 0 2.0 1e-06 
0.0 -0.4042 0 2.0 1e-06 
0.0 -0.4041 0 2.0 1e-06 
0.0 -0.404 0 2.0 1e-06 
0.0 -0.4039 0 2.0 1e-06 
0.0 -0.4038 0 2.0 1e-06 
0.0 -0.4037 0 2.0 1e-06 
0.0 -0.4036 0 2.0 1e-06 
0.0 -0.4035 0 2.0 1e-06 
0.0 -0.4034 0 2.0 1e-06 
0.0 -0.4033 0 2.0 1e-06 
0.0 -0.4032 0 2.0 1e-06 
0.0 -0.4031 0 2.0 1e-06 
0.0 -0.403 0 2.0 1e-06 
0.0 -0.4029 0 2.0 1e-06 
0.0 -0.4028 0 2.0 1e-06 
0.0 -0.4027 0 2.0 1e-06 
0.0 -0.4026 0 2.0 1e-06 
0.0 -0.4025 0 2.0 1e-06 
0.0 -0.4024 0 2.0 1e-06 
0.0 -0.4023 0 2.0 1e-06 
0.0 -0.4022 0 2.0 1e-06 
0.0 -0.4021 0 2.0 1e-06 
0.0 -0.402 0 2.0 1e-06 
0.0 -0.4019 0 2.0 1e-06 
0.0 -0.4018 0 2.0 1e-06 
0.0 -0.4017 0 2.0 1e-06 
0.0 -0.4016 0 2.0 1e-06 
0.0 -0.4015 0 2.0 1e-06 
0.0 -0.4014 0 2.0 1e-06 
0.0 -0.4013 0 2.0 1e-06 
0.0 -0.4012 0 2.0 1e-06 
0.0 -0.4011 0 2.0 1e-06 
0.0 -0.401 0 2.0 1e-06 
0.0 -0.4009 0 2.0 1e-06 
0.0 -0.4008 0 2.0 1e-06 
0.0 -0.4007 0 2.0 1e-06 
0.0 -0.4006 0 2.0 1e-06 
0.0 -0.4005 0 2.0 1e-06 
0.0 -0.4004 0 2.0 1e-06 
0.0 -0.4003 0 2.0 1e-06 
0.0 -0.4002 0 2.0 1e-06 
0.0 -0.4001 0 2.0 1e-06 
0.0 -0.4 0 2.0 1e-06 
0.0 -0.3999 0 2.0 1e-06 
0.0 -0.3998 0 2.0 1e-06 
0.0 -0.3997 0 2.0 1e-06 
0.0 -0.3996 0 2.0 1e-06 
0.0 -0.3995 0 2.0 1e-06 
0.0 -0.3994 0 2.0 1e-06 
0.0 -0.3993 0 2.0 1e-06 
0.0 -0.3992 0 2.0 1e-06 
0.0 -0.3991 0 2.0 1e-06 
0.0 -0.399 0 2.0 1e-06 
0.0 -0.3989 0 2.0 1e-06 
0.0 -0.3988 0 2.0 1e-06 
0.0 -0.3987 0 2.0 1e-06 
0.0 -0.3986 0 2.0 1e-06 
0.0 -0.3985 0 2.0 1e-06 
0.0 -0.3984 0 2.0 1e-06 
0.0 -0.3983 0 2.0 1e-06 
0.0 -0.3982 0 2.0 1e-06 
0.0 -0.3981 0 2.0 1e-06 
0.0 -0.398 0 2.0 1e-06 
0.0 -0.3979 0 2.0 1e-06 
0.0 -0.3978 0 2.0 1e-06 
0.0 -0.3977 0 2.0 1e-06 
0.0 -0.3976 0 2.0 1e-06 
0.0 -0.3975 0 2.0 1e-06 
0.0 -0.3974 0 2.0 1e-06 
0.0 -0.3973 0 2.0 1e-06 
0.0 -0.3972 0 2.0 1e-06 
0.0 -0.3971 0 2.0 1e-06 
0.0 -0.397 0 2.0 1e-06 
0.0 -0.3969 0 2.0 1e-06 
0.0 -0.3968 0 2.0 1e-06 
0.0 -0.3967 0 2.0 1e-06 
0.0 -0.3966 0 2.0 1e-06 
0.0 -0.3965 0 2.0 1e-06 
0.0 -0.3964 0 2.0 1e-06 
0.0 -0.3963 0 2.0 1e-06 
0.0 -0.3962 0 2.0 1e-06 
0.0 -0.3961 0 2.0 1e-06 
0.0 -0.396 0 2.0 1e-06 
0.0 -0.3959 0 2.0 1e-06 
0.0 -0.3958 0 2.0 1e-06 
0.0 -0.3957 0 2.0 1e-06 
0.0 -0.3956 0 2.0 1e-06 
0.0 -0.3955 0 2.0 1e-06 
0.0 -0.3954 0 2.0 1e-06 
0.0 -0.3953 0 2.0 1e-06 
0.0 -0.3952 0 2.0 1e-06 
0.0 -0.3951 0 2.0 1e-06 
0.0 -0.395 0 2.0 1e-06 
0.0 -0.3949 0 2.0 1e-06 
0.0 -0.3948 0 2.0 1e-06 
0.0 -0.3947 0 2.0 1e-06 
0.0 -0.3946 0 2.0 1e-06 
0.0 -0.3945 0 2.0 1e-06 
0.0 -0.3944 0 2.0 1e-06 
0.0 -0.3943 0 2.0 1e-06 
0.0 -0.3942 0 2.0 1e-06 
0.0 -0.3941 0 2.0 1e-06 
0.0 -0.394 0 2.0 1e-06 
0.0 -0.3939 0 2.0 1e-06 
0.0 -0.3938 0 2.0 1e-06 
0.0 -0.3937 0 2.0 1e-06 
0.0 -0.3936 0 2.0 1e-06 
0.0 -0.3935 0 2.0 1e-06 
0.0 -0.3934 0 2.0 1e-06 
0.0 -0.3933 0 2.0 1e-06 
0.0 -0.3932 0 2.0 1e-06 
0.0 -0.3931 0 2.0 1e-06 
0.0 -0.393 0 2.0 1e-06 
0.0 -0.3929 0 2.0 1e-06 
0.0 -0.3928 0 2.0 1e-06 
0.0 -0.3927 0 2.0 1e-06 
0.0 -0.3926 0 2.0 1e-06 
0.0 -0.3925 0 2.0 1e-06 
0.0 -0.3924 0 2.0 1e-06 
0.0 -0.3923 0 2.0 1e-06 
0.0 -0.3922 0 2.0 1e-06 
0.0 -0.3921 0 2.0 1e-06 
0.0 -0.392 0 2.0 1e-06 
0.0 -0.3919 0 2.0 1e-06 
0.0 -0.3918 0 2.0 1e-06 
0.0 -0.3917 0 2.0 1e-06 
0.0 -0.3916 0 2.0 1e-06 
0.0 -0.3915 0 2.0 1e-06 
0.0 -0.3914 0 2.0 1e-06 
0.0 -0.3913 0 2.0 1e-06 
0.0 -0.3912 0 2.0 1e-06 
0.0 -0.3911 0 2.0 1e-06 
0.0 -0.391 0 2.0 1e-06 
0.0 -0.3909 0 2.0 1e-06 
0.0 -0.3908 0 2.0 1e-06 
0.0 -0.3907 0 2.0 1e-06 
0.0 -0.3906 0 2.0 1e-06 
0.0 -0.3905 0 2.0 1e-06 
0.0 -0.3904 0 2.0 1e-06 
0.0 -0.3903 0 2.0 1e-06 
0.0 -0.3902 0 2.0 1e-06 
0.0 -0.3901 0 2.0 1e-06 
0.0 -0.39 0 2.0 1e-06 
0.0 -0.3899 0 2.0 1e-06 
0.0 -0.3898 0 2.0 1e-06 
0.0 -0.3897 0 2.0 1e-06 
0.0 -0.3896 0 2.0 1e-06 
0.0 -0.3895 0 2.0 1e-06 
0.0 -0.3894 0 2.0 1e-06 
0.0 -0.3893 0 2.0 1e-06 
0.0 -0.3892 0 2.0 1e-06 
0.0 -0.3891 0 2.0 1e-06 
0.0 -0.389 0 2.0 1e-06 
0.0 -0.3889 0 2.0 1e-06 
0.0 -0.3888 0 2.0 1e-06 
0.0 -0.3887 0 2.0 1e-06 
0.0 -0.3886 0 2.0 1e-06 
0.0 -0.3885 0 2.0 1e-06 
0.0 -0.3884 0 2.0 1e-06 
0.0 -0.3883 0 2.0 1e-06 
0.0 -0.3882 0 2.0 1e-06 
0.0 -0.3881 0 2.0 1e-06 
0.0 -0.388 0 2.0 1e-06 
0.0 -0.3879 0 2.0 1e-06 
0.0 -0.3878 0 2.0 1e-06 
0.0 -0.3877 0 2.0 1e-06 
0.0 -0.3876 0 2.0 1e-06 
0.0 -0.3875 0 2.0 1e-06 
0.0 -0.3874 0 2.0 1e-06 
0.0 -0.3873 0 2.0 1e-06 
0.0 -0.3872 0 2.0 1e-06 
0.0 -0.3871 0 2.0 1e-06 
0.0 -0.387 0 2.0 1e-06 
0.0 -0.3869 0 2.0 1e-06 
0.0 -0.3868 0 2.0 1e-06 
0.0 -0.3867 0 2.0 1e-06 
0.0 -0.3866 0 2.0 1e-06 
0.0 -0.3865 0 2.0 1e-06 
0.0 -0.3864 0 2.0 1e-06 
0.0 -0.3863 0 2.0 1e-06 
0.0 -0.3862 0 2.0 1e-06 
0.0 -0.3861 0 2.0 1e-06 
0.0 -0.386 0 2.0 1e-06 
0.0 -0.3859 0 2.0 1e-06 
0.0 -0.3858 0 2.0 1e-06 
0.0 -0.3857 0 2.0 1e-06 
0.0 -0.3856 0 2.0 1e-06 
0.0 -0.3855 0 2.0 1e-06 
0.0 -0.3854 0 2.0 1e-06 
0.0 -0.3853 0 2.0 1e-06 
0.0 -0.3852 0 2.0 1e-06 
0.0 -0.3851 0 2.0 1e-06 
0.0 -0.385 0 2.0 1e-06 
0.0 -0.3849 0 2.0 1e-06 
0.0 -0.3848 0 2.0 1e-06 
0.0 -0.3847 0 2.0 1e-06 
0.0 -0.3846 0 2.0 1e-06 
0.0 -0.3845 0 2.0 1e-06 
0.0 -0.3844 0 2.0 1e-06 
0.0 -0.3843 0 2.0 1e-06 
0.0 -0.3842 0 2.0 1e-06 
0.0 -0.3841 0 2.0 1e-06 
0.0 -0.384 0 2.0 1e-06 
0.0 -0.3839 0 2.0 1e-06 
0.0 -0.3838 0 2.0 1e-06 
0.0 -0.3837 0 2.0 1e-06 
0.0 -0.3836 0 2.0 1e-06 
0.0 -0.3835 0 2.0 1e-06 
0.0 -0.3834 0 2.0 1e-06 
0.0 -0.3833 0 2.0 1e-06 
0.0 -0.3832 0 2.0 1e-06 
0.0 -0.3831 0 2.0 1e-06 
0.0 -0.383 0 2.0 1e-06 
0.0 -0.3829 0 2.0 1e-06 
0.0 -0.3828 0 2.0 1e-06 
0.0 -0.3827 0 2.0 1e-06 
0.0 -0.3826 0 2.0 1e-06 
0.0 -0.3825 0 2.0 1e-06 
0.0 -0.3824 0 2.0 1e-06 
0.0 -0.3823 0 2.0 1e-06 
0.0 -0.3822 0 2.0 1e-06 
0.0 -0.3821 0 2.0 1e-06 
0.0 -0.382 0 2.0 1e-06 
0.0 -0.3819 0 2.0 1e-06 
0.0 -0.3818 0 2.0 1e-06 
0.0 -0.3817 0 2.0 1e-06 
0.0 -0.3816 0 2.0 1e-06 
0.0 -0.3815 0 2.0 1e-06 
0.0 -0.3814 0 2.0 1e-06 
0.0 -0.3813 0 2.0 1e-06 
0.0 -0.3812 0 2.0 1e-06 
0.0 -0.3811 0 2.0 1e-06 
0.0 -0.381 0 2.0 1e-06 
0.0 -0.3809 0 2.0 1e-06 
0.0 -0.3808 0 2.0 1e-06 
0.0 -0.3807 0 2.0 1e-06 
0.0 -0.3806 0 2.0 1e-06 
0.0 -0.3805 0 2.0 1e-06 
0.0 -0.3804 0 2.0 1e-06 
0.0 -0.3803 0 2.0 1e-06 
0.0 -0.3802 0 2.0 1e-06 
0.0 -0.3801 0 2.0 1e-06 
0.0 -0.38 0 2.0 1e-06 
0.0 -0.3799 0 2.0 1e-06 
0.0 -0.3798 0 2.0 1e-06 
0.0 -0.3797 0 2.0 1e-06 
0.0 -0.3796 0 2.0 1e-06 
0.0 -0.3795 0 2.0 1e-06 
0.0 -0.3794 0 2.0 1e-06 
0.0 -0.3793 0 2.0 1e-06 
0.0 -0.3792 0 2.0 1e-06 
0.0 -0.3791 0 2.0 1e-06 
0.0 -0.379 0 2.0 1e-06 
0.0 -0.3789 0 2.0 1e-06 
0.0 -0.3788 0 2.0 1e-06 
0.0 -0.3787 0 2.0 1e-06 
0.0 -0.3786 0 2.0 1e-06 
0.0 -0.3785 0 2.0 1e-06 
0.0 -0.3784 0 2.0 1e-06 
0.0 -0.3783 0 2.0 1e-06 
0.0 -0.3782 0 2.0 1e-06 
0.0 -0.3781 0 2.0 1e-06 
0.0 -0.378 0 2.0 1e-06 
0.0 -0.3779 0 2.0 1e-06 
0.0 -0.3778 0 2.0 1e-06 
0.0 -0.3777 0 2.0 1e-06 
0.0 -0.3776 0 2.0 1e-06 
0.0 -0.3775 0 2.0 1e-06 
0.0 -0.3774 0 2.0 1e-06 
0.0 -0.3773 0 2.0 1e-06 
0.0 -0.3772 0 2.0 1e-06 
0.0 -0.3771 0 2.0 1e-06 
0.0 -0.377 0 2.0 1e-06 
0.0 -0.3769 0 2.0 1e-06 
0.0 -0.3768 0 2.0 1e-06 
0.0 -0.3767 0 2.0 1e-06 
0.0 -0.3766 0 2.0 1e-06 
0.0 -0.3765 0 2.0 1e-06 
0.0 -0.3764 0 2.0 1e-06 
0.0 -0.3763 0 2.0 1e-06 
0.0 -0.3762 0 2.0 1e-06 
0.0 -0.3761 0 2.0 1e-06 
0.0 -0.376 0 2.0 1e-06 
0.0 -0.3759 0 2.0 1e-06 
0.0 -0.3758 0 2.0 1e-06 
0.0 -0.3757 0 2.0 1e-06 
0.0 -0.3756 0 2.0 1e-06 
0.0 -0.3755 0 2.0 1e-06 
0.0 -0.3754 0 2.0 1e-06 
0.0 -0.3753 0 2.0 1e-06 
0.0 -0.3752 0 2.0 1e-06 
0.0 -0.3751 0 2.0 1e-06 
0.0 -0.375 0 2.0 1e-06 
0.0 -0.3749 0 2.0 1e-06 
0.0 -0.3748 0 2.0 1e-06 
0.0 -0.3747 0 2.0 1e-06 
0.0 -0.3746 0 2.0 1e-06 
0.0 -0.3745 0 2.0 1e-06 
0.0 -0.3744 0 2.0 1e-06 
0.0 -0.3743 0 2.0 1e-06 
0.0 -0.3742 0 2.0 1e-06 
0.0 -0.3741 0 2.0 1e-06 
0.0 -0.374 0 2.0 1e-06 
0.0 -0.3739 0 2.0 1e-06 
0.0 -0.3738 0 2.0 1e-06 
0.0 -0.3737 0 2.0 1e-06 
0.0 -0.3736 0 2.0 1e-06 
0.0 -0.3735 0 2.0 1e-06 
0.0 -0.3734 0 2.0 1e-06 
0.0 -0.3733 0 2.0 1e-06 
0.0 -0.3732 0 2.0 1e-06 
0.0 -0.3731 0 2.0 1e-06 
0.0 -0.373 0 2.0 1e-06 
0.0 -0.3729 0 2.0 1e-06 
0.0 -0.3728 0 2.0 1e-06 
0.0 -0.3727 0 2.0 1e-06 
0.0 -0.3726 0 2.0 1e-06 
0.0 -0.3725 0 2.0 1e-06 
0.0 -0.3724 0 2.0 1e-06 
0.0 -0.3723 0 2.0 1e-06 
0.0 -0.3722 0 2.0 1e-06 
0.0 -0.3721 0 2.0 1e-06 
0.0 -0.372 0 2.0 1e-06 
0.0 -0.3719 0 2.0 1e-06 
0.0 -0.3718 0 2.0 1e-06 
0.0 -0.3717 0 2.0 1e-06 
0.0 -0.3716 0 2.0 1e-06 
0.0 -0.3715 0 2.0 1e-06 
0.0 -0.3714 0 2.0 1e-06 
0.0 -0.3713 0 2.0 1e-06 
0.0 -0.3712 0 2.0 1e-06 
0.0 -0.3711 0 2.0 1e-06 
0.0 -0.371 0 2.0 1e-06 
0.0 -0.3709 0 2.0 1e-06 
0.0 -0.3708 0 2.0 1e-06 
0.0 -0.3707 0 2.0 1e-06 
0.0 -0.3706 0 2.0 1e-06 
0.0 -0.3705 0 2.0 1e-06 
0.0 -0.3704 0 2.0 1e-06 
0.0 -0.3703 0 2.0 1e-06 
0.0 -0.3702 0 2.0 1e-06 
0.0 -0.3701 0 2.0 1e-06 
0.0 -0.37 0 2.0 1e-06 
0.0 -0.3699 0 2.0 1e-06 
0.0 -0.3698 0 2.0 1e-06 
0.0 -0.3697 0 2.0 1e-06 
0.0 -0.3696 0 2.0 1e-06 
0.0 -0.3695 0 2.0 1e-06 
0.0 -0.3694 0 2.0 1e-06 
0.0 -0.3693 0 2.0 1e-06 
0.0 -0.3692 0 2.0 1e-06 
0.0 -0.3691 0 2.0 1e-06 
0.0 -0.369 0 2.0 1e-06 
0.0 -0.3689 0 2.0 1e-06 
0.0 -0.3688 0 2.0 1e-06 
0.0 -0.3687 0 2.0 1e-06 
0.0 -0.3686 0 2.0 1e-06 
0.0 -0.3685 0 2.0 1e-06 
0.0 -0.3684 0 2.0 1e-06 
0.0 -0.3683 0 2.0 1e-06 
0.0 -0.3682 0 2.0 1e-06 
0.0 -0.3681 0 2.0 1e-06 
0.0 -0.368 0 2.0 1e-06 
0.0 -0.3679 0 2.0 1e-06 
0.0 -0.3678 0 2.0 1e-06 
0.0 -0.3677 0 2.0 1e-06 
0.0 -0.3676 0 2.0 1e-06 
0.0 -0.3675 0 2.0 1e-06 
0.0 -0.3674 0 2.0 1e-06 
0.0 -0.3673 0 2.0 1e-06 
0.0 -0.3672 0 2.0 1e-06 
0.0 -0.3671 0 2.0 1e-06 
0.0 -0.367 0 2.0 1e-06 
0.0 -0.3669 0 2.0 1e-06 
0.0 -0.3668 0 2.0 1e-06 
0.0 -0.3667 0 2.0 1e-06 
0.0 -0.3666 0 2.0 1e-06 
0.0 -0.3665 0 2.0 1e-06 
0.0 -0.3664 0 2.0 1e-06 
0.0 -0.3663 0 2.0 1e-06 
0.0 -0.3662 0 2.0 1e-06 
0.0 -0.3661 0 2.0 1e-06 
0.0 -0.366 0 2.0 1e-06 
0.0 -0.3659 0 2.0 1e-06 
0.0 -0.3658 0 2.0 1e-06 
0.0 -0.3657 0 2.0 1e-06 
0.0 -0.3656 0 2.0 1e-06 
0.0 -0.3655 0 2.0 1e-06 
0.0 -0.3654 0 2.0 1e-06 
0.0 -0.3653 0 2.0 1e-06 
0.0 -0.3652 0 2.0 1e-06 
0.0 -0.3651 0 2.0 1e-06 
0.0 -0.365 0 2.0 1e-06 
0.0 -0.3649 0 2.0 1e-06 
0.0 -0.3648 0 2.0 1e-06 
0.0 -0.3647 0 2.0 1e-06 
0.0 -0.3646 0 2.0 1e-06 
0.0 -0.3645 0 2.0 1e-06 
0.0 -0.3644 0 2.0 1e-06 
0.0 -0.3643 0 2.0 1e-06 
0.0 -0.3642 0 2.0 1e-06 
0.0 -0.3641 0 2.0 1e-06 
0.0 -0.364 0 2.0 1e-06 
0.0 -0.3639 0 2.0 1e-06 
0.0 -0.3638 0 2.0 1e-06 
0.0 -0.3637 0 2.0 1e-06 
0.0 -0.3636 0 2.0 1e-06 
0.0 -0.3635 0 2.0 1e-06 
0.0 -0.3634 0 2.0 1e-06 
0.0 -0.3633 0 2.0 1e-06 
0.0 -0.3632 0 2.0 1e-06 
0.0 -0.3631 0 2.0 1e-06 
0.0 -0.363 0 2.0 1e-06 
0.0 -0.3629 0 2.0 1e-06 
0.0 -0.3628 0 2.0 1e-06 
0.0 -0.3627 0 2.0 1e-06 
0.0 -0.3626 0 2.0 1e-06 
0.0 -0.3625 0 2.0 1e-06 
0.0 -0.3624 0 2.0 1e-06 
0.0 -0.3623 0 2.0 1e-06 
0.0 -0.3622 0 2.0 1e-06 
0.0 -0.3621 0 2.0 1e-06 
0.0 -0.362 0 2.0 1e-06 
0.0 -0.3619 0 2.0 1e-06 
0.0 -0.3618 0 2.0 1e-06 
0.0 -0.3617 0 2.0 1e-06 
0.0 -0.3616 0 2.0 1e-06 
0.0 -0.3615 0 2.0 1e-06 
0.0 -0.3614 0 2.0 1e-06 
0.0 -0.3613 0 2.0 1e-06 
0.0 -0.3612 0 2.0 1e-06 
0.0 -0.3611 0 2.0 1e-06 
0.0 -0.361 0 2.0 1e-06 
0.0 -0.3609 0 2.0 1e-06 
0.0 -0.3608 0 2.0 1e-06 
0.0 -0.3607 0 2.0 1e-06 
0.0 -0.3606 0 2.0 1e-06 
0.0 -0.3605 0 2.0 1e-06 
0.0 -0.3604 0 2.0 1e-06 
0.0 -0.3603 0 2.0 1e-06 
0.0 -0.3602 0 2.0 1e-06 
0.0 -0.3601 0 2.0 1e-06 
0.0 -0.36 0 2.0 1e-06 
0.0 -0.3599 0 2.0 1e-06 
0.0 -0.3598 0 2.0 1e-06 
0.0 -0.3597 0 2.0 1e-06 
0.0 -0.3596 0 2.0 1e-06 
0.0 -0.3595 0 2.0 1e-06 
0.0 -0.3594 0 2.0 1e-06 
0.0 -0.3593 0 2.0 1e-06 
0.0 -0.3592 0 2.0 1e-06 
0.0 -0.3591 0 2.0 1e-06 
0.0 -0.359 0 2.0 1e-06 
0.0 -0.3589 0 2.0 1e-06 
0.0 -0.3588 0 2.0 1e-06 
0.0 -0.3587 0 2.0 1e-06 
0.0 -0.3586 0 2.0 1e-06 
0.0 -0.3585 0 2.0 1e-06 
0.0 -0.3584 0 2.0 1e-06 
0.0 -0.3583 0 2.0 1e-06 
0.0 -0.3582 0 2.0 1e-06 
0.0 -0.3581 0 2.0 1e-06 
0.0 -0.358 0 2.0 1e-06 
0.0 -0.3579 0 2.0 1e-06 
0.0 -0.3578 0 2.0 1e-06 
0.0 -0.3577 0 2.0 1e-06 
0.0 -0.3576 0 2.0 1e-06 
0.0 -0.3575 0 2.0 1e-06 
0.0 -0.3574 0 2.0 1e-06 
0.0 -0.3573 0 2.0 1e-06 
0.0 -0.3572 0 2.0 1e-06 
0.0 -0.3571 0 2.0 1e-06 
0.0 -0.357 0 2.0 1e-06 
0.0 -0.3569 0 2.0 1e-06 
0.0 -0.3568 0 2.0 1e-06 
0.0 -0.3567 0 2.0 1e-06 
0.0 -0.3566 0 2.0 1e-06 
0.0 -0.3565 0 2.0 1e-06 
0.0 -0.3564 0 2.0 1e-06 
0.0 -0.3563 0 2.0 1e-06 
0.0 -0.3562 0 2.0 1e-06 
0.0 -0.3561 0 2.0 1e-06 
0.0 -0.356 0 2.0 1e-06 
0.0 -0.3559 0 2.0 1e-06 
0.0 -0.3558 0 2.0 1e-06 
0.0 -0.3557 0 2.0 1e-06 
0.0 -0.3556 0 2.0 1e-06 
0.0 -0.3555 0 2.0 1e-06 
0.0 -0.3554 0 2.0 1e-06 
0.0 -0.3553 0 2.0 1e-06 
0.0 -0.3552 0 2.0 1e-06 
0.0 -0.3551 0 2.0 1e-06 
0.0 -0.355 0 2.0 1e-06 
0.0 -0.3549 0 2.0 1e-06 
0.0 -0.3548 0 2.0 1e-06 
0.0 -0.3547 0 2.0 1e-06 
0.0 -0.3546 0 2.0 1e-06 
0.0 -0.3545 0 2.0 1e-06 
0.0 -0.3544 0 2.0 1e-06 
0.0 -0.3543 0 2.0 1e-06 
0.0 -0.3542 0 2.0 1e-06 
0.0 -0.3541 0 2.0 1e-06 
0.0 -0.354 0 2.0 1e-06 
0.0 -0.3539 0 2.0 1e-06 
0.0 -0.3538 0 2.0 1e-06 
0.0 -0.3537 0 2.0 1e-06 
0.0 -0.3536 0 2.0 1e-06 
0.0 -0.3535 0 2.0 1e-06 
0.0 -0.3534 0 2.0 1e-06 
0.0 -0.3533 0 2.0 1e-06 
0.0 -0.3532 0 2.0 1e-06 
0.0 -0.3531 0 2.0 1e-06 
0.0 -0.353 0 2.0 1e-06 
0.0 -0.3529 0 2.0 1e-06 
0.0 -0.3528 0 2.0 1e-06 
0.0 -0.3527 0 2.0 1e-06 
0.0 -0.3526 0 2.0 1e-06 
0.0 -0.3525 0 2.0 1e-06 
0.0 -0.3524 0 2.0 1e-06 
0.0 -0.3523 0 2.0 1e-06 
0.0 -0.3522 0 2.0 1e-06 
0.0 -0.3521 0 2.0 1e-06 
0.0 -0.352 0 2.0 1e-06 
0.0 -0.3519 0 2.0 1e-06 
0.0 -0.3518 0 2.0 1e-06 
0.0 -0.3517 0 2.0 1e-06 
0.0 -0.3516 0 2.0 1e-06 
0.0 -0.3515 0 2.0 1e-06 
0.0 -0.3514 0 2.0 1e-06 
0.0 -0.3513 0 2.0 1e-06 
0.0 -0.3512 0 2.0 1e-06 
0.0 -0.3511 0 2.0 1e-06 
0.0 -0.351 0 2.0 1e-06 
0.0 -0.3509 0 2.0 1e-06 
0.0 -0.3508 0 2.0 1e-06 
0.0 -0.3507 0 2.0 1e-06 
0.0 -0.3506 0 2.0 1e-06 
0.0 -0.3505 0 2.0 1e-06 
0.0 -0.3504 0 2.0 1e-06 
0.0 -0.3503 0 2.0 1e-06 
0.0 -0.3502 0 2.0 1e-06 
0.0 -0.3501 0 2.0 1e-06 
0.0 -0.35 0 2.0 1e-06 
0.0 -0.3499 0 2.0 1e-06 
0.0 -0.3498 0 2.0 1e-06 
0.0 -0.3497 0 2.0 1e-06 
0.0 -0.3496 0 2.0 1e-06 
0.0 -0.3495 0 2.0 1e-06 
0.0 -0.3494 0 2.0 1e-06 
0.0 -0.3493 0 2.0 1e-06 
0.0 -0.3492 0 2.0 1e-06 
0.0 -0.3491 0 2.0 1e-06 
0.0 -0.349 0 2.0 1e-06 
0.0 -0.3489 0 2.0 1e-06 
0.0 -0.3488 0 2.0 1e-06 
0.0 -0.3487 0 2.0 1e-06 
0.0 -0.3486 0 2.0 1e-06 
0.0 -0.3485 0 2.0 1e-06 
0.0 -0.3484 0 2.0 1e-06 
0.0 -0.3483 0 2.0 1e-06 
0.0 -0.3482 0 2.0 1e-06 
0.0 -0.3481 0 2.0 1e-06 
0.0 -0.348 0 2.0 1e-06 
0.0 -0.3479 0 2.0 1e-06 
0.0 -0.3478 0 2.0 1e-06 
0.0 -0.3477 0 2.0 1e-06 
0.0 -0.3476 0 2.0 1e-06 
0.0 -0.3475 0 2.0 1e-06 
0.0 -0.3474 0 2.0 1e-06 
0.0 -0.3473 0 2.0 1e-06 
0.0 -0.3472 0 2.0 1e-06 
0.0 -0.3471 0 2.0 1e-06 
0.0 -0.347 0 2.0 1e-06 
0.0 -0.3469 0 2.0 1e-06 
0.0 -0.3468 0 2.0 1e-06 
0.0 -0.3467 0 2.0 1e-06 
0.0 -0.3466 0 2.0 1e-06 
0.0 -0.3465 0 2.0 1e-06 
0.0 -0.3464 0 2.0 1e-06 
0.0 -0.3463 0 2.0 1e-06 
0.0 -0.3462 0 2.0 1e-06 
0.0 -0.3461 0 2.0 1e-06 
0.0 -0.346 0 2.0 1e-06 
0.0 -0.3459 0 2.0 1e-06 
0.0 -0.3458 0 2.0 1e-06 
0.0 -0.3457 0 2.0 1e-06 
0.0 -0.3456 0 2.0 1e-06 
0.0 -0.3455 0 2.0 1e-06 
0.0 -0.3454 0 2.0 1e-06 
0.0 -0.3453 0 2.0 1e-06 
0.0 -0.3452 0 2.0 1e-06 
0.0 -0.3451 0 2.0 1e-06 
0.0 -0.345 0 2.0 1e-06 
0.0 -0.3449 0 2.0 1e-06 
0.0 -0.3448 0 2.0 1e-06 
0.0 -0.3447 0 2.0 1e-06 
0.0 -0.3446 0 2.0 1e-06 
0.0 -0.3445 0 2.0 1e-06 
0.0 -0.3444 0 2.0 1e-06 
0.0 -0.3443 0 2.0 1e-06 
0.0 -0.3442 0 2.0 1e-06 
0.0 -0.3441 0 2.0 1e-06 
0.0 -0.344 0 2.0 1e-06 
0.0 -0.3439 0 2.0 1e-06 
0.0 -0.3438 0 2.0 1e-06 
0.0 -0.3437 0 2.0 1e-06 
0.0 -0.3436 0 2.0 1e-06 
0.0 -0.3435 0 2.0 1e-06 
0.0 -0.3434 0 2.0 1e-06 
0.0 -0.3433 0 2.0 1e-06 
0.0 -0.3432 0 2.0 1e-06 
0.0 -0.3431 0 2.0 1e-06 
0.0 -0.343 0 2.0 1e-06 
0.0 -0.3429 0 2.0 1e-06 
0.0 -0.3428 0 2.0 1e-06 
0.0 -0.3427 0 2.0 1e-06 
0.0 -0.3426 0 2.0 1e-06 
0.0 -0.3425 0 2.0 1e-06 
0.0 -0.3424 0 2.0 1e-06 
0.0 -0.3423 0 2.0 1e-06 
0.0 -0.3422 0 2.0 1e-06 
0.0 -0.3421 0 2.0 1e-06 
0.0 -0.342 0 2.0 1e-06 
0.0 -0.3419 0 2.0 1e-06 
0.0 -0.3418 0 2.0 1e-06 
0.0 -0.3417 0 2.0 1e-06 
0.0 -0.3416 0 2.0 1e-06 
0.0 -0.3415 0 2.0 1e-06 
0.0 -0.3414 0 2.0 1e-06 
0.0 -0.3413 0 2.0 1e-06 
0.0 -0.3412 0 2.0 1e-06 
0.0 -0.3411 0 2.0 1e-06 
0.0 -0.341 0 2.0 1e-06 
0.0 -0.3409 0 2.0 1e-06 
0.0 -0.3408 0 2.0 1e-06 
0.0 -0.3407 0 2.0 1e-06 
0.0 -0.3406 0 2.0 1e-06 
0.0 -0.3405 0 2.0 1e-06 
0.0 -0.3404 0 2.0 1e-06 
0.0 -0.3403 0 2.0 1e-06 
0.0 -0.3402 0 2.0 1e-06 
0.0 -0.3401 0 2.0 1e-06 
0.0 -0.34 0 2.0 1e-06 
0.0 -0.3399 0 2.0 1e-06 
0.0 -0.3398 0 2.0 1e-06 
0.0 -0.3397 0 2.0 1e-06 
0.0 -0.3396 0 2.0 1e-06 
0.0 -0.3395 0 2.0 1e-06 
0.0 -0.3394 0 2.0 1e-06 
0.0 -0.3393 0 2.0 1e-06 
0.0 -0.3392 0 2.0 1e-06 
0.0 -0.3391 0 2.0 1e-06 
0.0 -0.339 0 2.0 1e-06 
0.0 -0.3389 0 2.0 1e-06 
0.0 -0.3388 0 2.0 1e-06 
0.0 -0.3387 0 2.0 1e-06 
0.0 -0.3386 0 2.0 1e-06 
0.0 -0.3385 0 2.0 1e-06 
0.0 -0.3384 0 2.0 1e-06 
0.0 -0.3383 0 2.0 1e-06 
0.0 -0.3382 0 2.0 1e-06 
0.0 -0.3381 0 2.0 1e-06 
0.0 -0.338 0 2.0 1e-06 
0.0 -0.3379 0 2.0 1e-06 
0.0 -0.3378 0 2.0 1e-06 
0.0 -0.3377 0 2.0 1e-06 
0.0 -0.3376 0 2.0 1e-06 
0.0 -0.3375 0 2.0 1e-06 
0.0 -0.3374 0 2.0 1e-06 
0.0 -0.3373 0 2.0 1e-06 
0.0 -0.3372 0 2.0 1e-06 
0.0 -0.3371 0 2.0 1e-06 
0.0 -0.337 0 2.0 1e-06 
0.0 -0.3369 0 2.0 1e-06 
0.0 -0.3368 0 2.0 1e-06 
0.0 -0.3367 0 2.0 1e-06 
0.0 -0.3366 0 2.0 1e-06 
0.0 -0.3365 0 2.0 1e-06 
0.0 -0.3364 0 2.0 1e-06 
0.0 -0.3363 0 2.0 1e-06 
0.0 -0.3362 0 2.0 1e-06 
0.0 -0.3361 0 2.0 1e-06 
0.0 -0.336 0 2.0 1e-06 
0.0 -0.3359 0 2.0 1e-06 
0.0 -0.3358 0 2.0 1e-06 
0.0 -0.3357 0 2.0 1e-06 
0.0 -0.3356 0 2.0 1e-06 
0.0 -0.3355 0 2.0 1e-06 
0.0 -0.3354 0 2.0 1e-06 
0.0 -0.3353 0 2.0 1e-06 
0.0 -0.3352 0 2.0 1e-06 
0.0 -0.3351 0 2.0 1e-06 
0.0 -0.335 0 2.0 1e-06 
0.0 -0.3349 0 2.0 1e-06 
0.0 -0.3348 0 2.0 1e-06 
0.0 -0.3347 0 2.0 1e-06 
0.0 -0.3346 0 2.0 1e-06 
0.0 -0.3345 0 2.0 1e-06 
0.0 -0.3344 0 2.0 1e-06 
0.0 -0.3343 0 2.0 1e-06 
0.0 -0.3342 0 2.0 1e-06 
0.0 -0.3341 0 2.0 1e-06 
0.0 -0.334 0 2.0 1e-06 
0.0 -0.3339 0 2.0 1e-06 
0.0 -0.3338 0 2.0 1e-06 
0.0 -0.3337 0 2.0 1e-06 
0.0 -0.3336 0 2.0 1e-06 
0.0 -0.3335 0 2.0 1e-06 
0.0 -0.3334 0 2.0 1e-06 
0.0 -0.3333 0 2.0 1e-06 
0.0 -0.3332 0 2.0 1e-06 
0.0 -0.3331 0 2.0 1e-06 
0.0 -0.333 0 2.0 1e-06 
0.0 -0.3329 0 2.0 1e-06 
0.0 -0.3328 0 2.0 1e-06 
0.0 -0.3327 0 2.0 1e-06 
0.0 -0.3326 0 2.0 1e-06 
0.0 -0.3325 0 2.0 1e-06 
0.0 -0.3324 0 2.0 1e-06 
0.0 -0.3323 0 2.0 1e-06 
0.0 -0.3322 0 2.0 1e-06 
0.0 -0.3321 0 2.0 1e-06 
0.0 -0.332 0 2.0 1e-06 
0.0 -0.3319 0 2.0 1e-06 
0.0 -0.3318 0 2.0 1e-06 
0.0 -0.3317 0 2.0 1e-06 
0.0 -0.3316 0 2.0 1e-06 
0.0 -0.3315 0 2.0 1e-06 
0.0 -0.3314 0 2.0 1e-06 
0.0 -0.3313 0 2.0 1e-06 
0.0 -0.3312 0 2.0 1e-06 
0.0 -0.3311 0 2.0 1e-06 
0.0 -0.331 0 2.0 1e-06 
0.0 -0.3309 0 2.0 1e-06 
0.0 -0.3308 0 2.0 1e-06 
0.0 -0.3307 0 2.0 1e-06 
0.0 -0.3306 0 2.0 1e-06 
0.0 -0.3305 0 2.0 1e-06 
0.0 -0.3304 0 2.0 1e-06 
0.0 -0.3303 0 2.0 1e-06 
0.0 -0.3302 0 2.0 1e-06 
0.0 -0.3301 0 2.0 1e-06 
0.0 -0.33 0 2.0 1e-06 
0.0 -0.3299 0 2.0 1e-06 
0.0 -0.3298 0 2.0 1e-06 
0.0 -0.3297 0 2.0 1e-06 
0.0 -0.3296 0 2.0 1e-06 
0.0 -0.3295 0 2.0 1e-06 
0.0 -0.3294 0 2.0 1e-06 
0.0 -0.3293 0 2.0 1e-06 
0.0 -0.3292 0 2.0 1e-06 
0.0 -0.3291 0 2.0 1e-06 
0.0 -0.329 0 2.0 1e-06 
0.0 -0.3289 0 2.0 1e-06 
0.0 -0.3288 0 2.0 1e-06 
0.0 -0.3287 0 2.0 1e-06 
0.0 -0.3286 0 2.0 1e-06 
0.0 -0.3285 0 2.0 1e-06 
0.0 -0.3284 0 2.0 1e-06 
0.0 -0.3283 0 2.0 1e-06 
0.0 -0.3282 0 2.0 1e-06 
0.0 -0.3281 0 2.0 1e-06 
0.0 -0.328 0 2.0 1e-06 
0.0 -0.3279 0 2.0 1e-06 
0.0 -0.3278 0 2.0 1e-06 
0.0 -0.3277 0 2.0 1e-06 
0.0 -0.3276 0 2.0 1e-06 
0.0 -0.3275 0 2.0 1e-06 
0.0 -0.3274 0 2.0 1e-06 
0.0 -0.3273 0 2.0 1e-06 
0.0 -0.3272 0 2.0 1e-06 
0.0 -0.3271 0 2.0 1e-06 
0.0 -0.327 0 2.0 1e-06 
0.0 -0.3269 0 2.0 1e-06 
0.0 -0.3268 0 2.0 1e-06 
0.0 -0.3267 0 2.0 1e-06 
0.0 -0.3266 0 2.0 1e-06 
0.0 -0.3265 0 2.0 1e-06 
0.0 -0.3264 0 2.0 1e-06 
0.0 -0.3263 0 2.0 1e-06 
0.0 -0.3262 0 2.0 1e-06 
0.0 -0.3261 0 2.0 1e-06 
0.0 -0.326 0 2.0 1e-06 
0.0 -0.3259 0 2.0 1e-06 
0.0 -0.3258 0 2.0 1e-06 
0.0 -0.3257 0 2.0 1e-06 
0.0 -0.3256 0 2.0 1e-06 
0.0 -0.3255 0 2.0 1e-06 
0.0 -0.3254 0 2.0 1e-06 
0.0 -0.3253 0 2.0 1e-06 
0.0 -0.3252 0 2.0 1e-06 
0.0 -0.3251 0 2.0 1e-06 
0.0 -0.325 0 2.0 1e-06 
0.0 -0.3249 0 2.0 1e-06 
0.0 -0.3248 0 2.0 1e-06 
0.0 -0.3247 0 2.0 1e-06 
0.0 -0.3246 0 2.0 1e-06 
0.0 -0.3245 0 2.0 1e-06 
0.0 -0.3244 0 2.0 1e-06 
0.0 -0.3243 0 2.0 1e-06 
0.0 -0.3242 0 2.0 1e-06 
0.0 -0.3241 0 2.0 1e-06 
0.0 -0.324 0 2.0 1e-06 
0.0 -0.3239 0 2.0 1e-06 
0.0 -0.3238 0 2.0 1e-06 
0.0 -0.3237 0 2.0 1e-06 
0.0 -0.3236 0 2.0 1e-06 
0.0 -0.3235 0 2.0 1e-06 
0.0 -0.3234 0 2.0 1e-06 
0.0 -0.3233 0 2.0 1e-06 
0.0 -0.3232 0 2.0 1e-06 
0.0 -0.3231 0 2.0 1e-06 
0.0 -0.323 0 2.0 1e-06 
0.0 -0.3229 0 2.0 1e-06 
0.0 -0.3228 0 2.0 1e-06 
0.0 -0.3227 0 2.0 1e-06 
0.0 -0.3226 0 2.0 1e-06 
0.0 -0.3225 0 2.0 1e-06 
0.0 -0.3224 0 2.0 1e-06 
0.0 -0.3223 0 2.0 1e-06 
0.0 -0.3222 0 2.0 1e-06 
0.0 -0.3221 0 2.0 1e-06 
0.0 -0.322 0 2.0 1e-06 
0.0 -0.3219 0 2.0 1e-06 
0.0 -0.3218 0 2.0 1e-06 
0.0 -0.3217 0 2.0 1e-06 
0.0 -0.3216 0 2.0 1e-06 
0.0 -0.3215 0 2.0 1e-06 
0.0 -0.3214 0 2.0 1e-06 
0.0 -0.3213 0 2.0 1e-06 
0.0 -0.3212 0 2.0 1e-06 
0.0 -0.3211 0 2.0 1e-06 
0.0 -0.321 0 2.0 1e-06 
0.0 -0.3209 0 2.0 1e-06 
0.0 -0.3208 0 2.0 1e-06 
0.0 -0.3207 0 2.0 1e-06 
0.0 -0.3206 0 2.0 1e-06 
0.0 -0.3205 0 2.0 1e-06 
0.0 -0.3204 0 2.0 1e-06 
0.0 -0.3203 0 2.0 1e-06 
0.0 -0.3202 0 2.0 1e-06 
0.0 -0.3201 0 2.0 1e-06 
0.0 -0.32 0 2.0 1e-06 
0.0 -0.3199 0 2.0 1e-06 
0.0 -0.3198 0 2.0 1e-06 
0.0 -0.3197 0 2.0 1e-06 
0.0 -0.3196 0 2.0 1e-06 
0.0 -0.3195 0 2.0 1e-06 
0.0 -0.3194 0 2.0 1e-06 
0.0 -0.3193 0 2.0 1e-06 
0.0 -0.3192 0 2.0 1e-06 
0.0 -0.3191 0 2.0 1e-06 
0.0 -0.319 0 2.0 1e-06 
0.0 -0.3189 0 2.0 1e-06 
0.0 -0.3188 0 2.0 1e-06 
0.0 -0.3187 0 2.0 1e-06 
0.0 -0.3186 0 2.0 1e-06 
0.0 -0.3185 0 2.0 1e-06 
0.0 -0.3184 0 2.0 1e-06 
0.0 -0.3183 0 2.0 1e-06 
0.0 -0.3182 0 2.0 1e-06 
0.0 -0.3181 0 2.0 1e-06 
0.0 -0.318 0 2.0 1e-06 
0.0 -0.3179 0 2.0 1e-06 
0.0 -0.3178 0 2.0 1e-06 
0.0 -0.3177 0 2.0 1e-06 
0.0 -0.3176 0 2.0 1e-06 
0.0 -0.3175 0 2.0 1e-06 
0.0 -0.3174 0 2.0 1e-06 
0.0 -0.3173 0 2.0 1e-06 
0.0 -0.3172 0 2.0 1e-06 
0.0 -0.3171 0 2.0 1e-06 
0.0 -0.317 0 2.0 1e-06 
0.0 -0.3169 0 2.0 1e-06 
0.0 -0.3168 0 2.0 1e-06 
0.0 -0.3167 0 2.0 1e-06 
0.0 -0.3166 0 2.0 1e-06 
0.0 -0.3165 0 2.0 1e-06 
0.0 -0.3164 0 2.0 1e-06 
0.0 -0.3163 0 2.0 1e-06 
0.0 -0.3162 0 2.0 1e-06 
0.0 -0.3161 0 2.0 1e-06 
0.0 -0.316 0 2.0 1e-06 
0.0 -0.3159 0 2.0 1e-06 
0.0 -0.3158 0 2.0 1e-06 
0.0 -0.3157 0 2.0 1e-06 
0.0 -0.3156 0 2.0 1e-06 
0.0 -0.3155 0 2.0 1e-06 
0.0 -0.3154 0 2.0 1e-06 
0.0 -0.3153 0 2.0 1e-06 
0.0 -0.3152 0 2.0 1e-06 
0.0 -0.3151 0 2.0 1e-06 
0.0 -0.315 0 2.0 1e-06 
0.0 -0.3149 0 2.0 1e-06 
0.0 -0.3148 0 2.0 1e-06 
0.0 -0.3147 0 2.0 1e-06 
0.0 -0.3146 0 2.0 1e-06 
0.0 -0.3145 0 2.0 1e-06 
0.0 -0.3144 0 2.0 1e-06 
0.0 -0.3143 0 2.0 1e-06 
0.0 -0.3142 0 2.0 1e-06 
0.0 -0.3141 0 2.0 1e-06 
0.0 -0.314 0 2.0 1e-06 
0.0 -0.3139 0 2.0 1e-06 
0.0 -0.3138 0 2.0 1e-06 
0.0 -0.3137 0 2.0 1e-06 
0.0 -0.3136 0 2.0 1e-06 
0.0 -0.3135 0 2.0 1e-06 
0.0 -0.3134 0 2.0 1e-06 
0.0 -0.3133 0 2.0 1e-06 
0.0 -0.3132 0 2.0 1e-06 
0.0 -0.3131 0 2.0 1e-06 
0.0 -0.313 0 2.0 1e-06 
0.0 -0.3129 0 2.0 1e-06 
0.0 -0.3128 0 2.0 1e-06 
0.0 -0.3127 0 2.0 1e-06 
0.0 -0.3126 0 2.0 1e-06 
0.0 -0.3125 0 2.0 1e-06 
0.0 -0.3124 0 2.0 1e-06 
0.0 -0.3123 0 2.0 1e-06 
0.0 -0.3122 0 2.0 1e-06 
0.0 -0.3121 0 2.0 1e-06 
0.0 -0.312 0 2.0 1e-06 
0.0 -0.3119 0 2.0 1e-06 
0.0 -0.3118 0 2.0 1e-06 
0.0 -0.3117 0 2.0 1e-06 
0.0 -0.3116 0 2.0 1e-06 
0.0 -0.3115 0 2.0 1e-06 
0.0 -0.3114 0 2.0 1e-06 
0.0 -0.3113 0 2.0 1e-06 
0.0 -0.3112 0 2.0 1e-06 
0.0 -0.3111 0 2.0 1e-06 
0.0 -0.311 0 2.0 1e-06 
0.0 -0.3109 0 2.0 1e-06 
0.0 -0.3108 0 2.0 1e-06 
0.0 -0.3107 0 2.0 1e-06 
0.0 -0.3106 0 2.0 1e-06 
0.0 -0.3105 0 2.0 1e-06 
0.0 -0.3104 0 2.0 1e-06 
0.0 -0.3103 0 2.0 1e-06 
0.0 -0.3102 0 2.0 1e-06 
0.0 -0.3101 0 2.0 1e-06 
0.0 -0.31 0 2.0 1e-06 
0.0 -0.3099 0 2.0 1e-06 
0.0 -0.3098 0 2.0 1e-06 
0.0 -0.3097 0 2.0 1e-06 
0.0 -0.3096 0 2.0 1e-06 
0.0 -0.3095 0 2.0 1e-06 
0.0 -0.3094 0 2.0 1e-06 
0.0 -0.3093 0 2.0 1e-06 
0.0 -0.3092 0 2.0 1e-06 
0.0 -0.3091 0 2.0 1e-06 
0.0 -0.309 0 2.0 1e-06 
0.0 -0.3089 0 2.0 1e-06 
0.0 -0.3088 0 2.0 1e-06 
0.0 -0.3087 0 2.0 1e-06 
0.0 -0.3086 0 2.0 1e-06 
0.0 -0.3085 0 2.0 1e-06 
0.0 -0.3084 0 2.0 1e-06 
0.0 -0.3083 0 2.0 1e-06 
0.0 -0.3082 0 2.0 1e-06 
0.0 -0.3081 0 2.0 1e-06 
0.0 -0.308 0 2.0 1e-06 
0.0 -0.3079 0 2.0 1e-06 
0.0 -0.3078 0 2.0 1e-06 
0.0 -0.3077 0 2.0 1e-06 
0.0 -0.3076 0 2.0 1e-06 
0.0 -0.3075 0 2.0 1e-06 
0.0 -0.3074 0 2.0 1e-06 
0.0 -0.3073 0 2.0 1e-06 
0.0 -0.3072 0 2.0 1e-06 
0.0 -0.3071 0 2.0 1e-06 
0.0 -0.307 0 2.0 1e-06 
0.0 -0.3069 0 2.0 1e-06 
0.0 -0.3068 0 2.0 1e-06 
0.0 -0.3067 0 2.0 1e-06 
0.0 -0.3066 0 2.0 1e-06 
0.0 -0.3065 0 2.0 1e-06 
0.0 -0.3064 0 2.0 1e-06 
0.0 -0.3063 0 2.0 1e-06 
0.0 -0.3062 0 2.0 1e-06 
0.0 -0.3061 0 2.0 1e-06 
0.0 -0.306 0 2.0 1e-06 
0.0 -0.3059 0 2.0 1e-06 
0.0 -0.3058 0 2.0 1e-06 
0.0 -0.3057 0 2.0 1e-06 
0.0 -0.3056 0 2.0 1e-06 
0.0 -0.3055 0 2.0 1e-06 
0.0 -0.3054 0 2.0 1e-06 
0.0 -0.3053 0 2.0 1e-06 
0.0 -0.3052 0 2.0 1e-06 
0.0 -0.3051 0 2.0 1e-06 
0.0 -0.305 0 2.0 1e-06 
0.0 -0.3049 0 2.0 1e-06 
0.0 -0.3048 0 2.0 1e-06 
0.0 -0.3047 0 2.0 1e-06 
0.0 -0.3046 0 2.0 1e-06 
0.0 -0.3045 0 2.0 1e-06 
0.0 -0.3044 0 2.0 1e-06 
0.0 -0.3043 0 2.0 1e-06 
0.0 -0.3042 0 2.0 1e-06 
0.0 -0.3041 0 2.0 1e-06 
0.0 -0.304 0 2.0 1e-06 
0.0 -0.3039 0 2.0 1e-06 
0.0 -0.3038 0 2.0 1e-06 
0.0 -0.3037 0 2.0 1e-06 
0.0 -0.3036 0 2.0 1e-06 
0.0 -0.3035 0 2.0 1e-06 
0.0 -0.3034 0 2.0 1e-06 
0.0 -0.3033 0 2.0 1e-06 
0.0 -0.3032 0 2.0 1e-06 
0.0 -0.3031 0 2.0 1e-06 
0.0 -0.303 0 2.0 1e-06 
0.0 -0.3029 0 2.0 1e-06 
0.0 -0.3028 0 2.0 1e-06 
0.0 -0.3027 0 2.0 1e-06 
0.0 -0.3026 0 2.0 1e-06 
0.0 -0.3025 0 2.0 1e-06 
0.0 -0.3024 0 2.0 1e-06 
0.0 -0.3023 0 2.0 1e-06 
0.0 -0.3022 0 2.0 1e-06 
0.0 -0.3021 0 2.0 1e-06 
0.0 -0.302 0 2.0 1e-06 
0.0 -0.3019 0 2.0 1e-06 
0.0 -0.3018 0 2.0 1e-06 
0.0 -0.3017 0 2.0 1e-06 
0.0 -0.3016 0 2.0 1e-06 
0.0 -0.3015 0 2.0 1e-06 
0.0 -0.3014 0 2.0 1e-06 
0.0 -0.3013 0 2.0 1e-06 
0.0 -0.3012 0 2.0 1e-06 
0.0 -0.3011 0 2.0 1e-06 
0.0 -0.301 0 2.0 1e-06 
0.0 -0.3009 0 2.0 1e-06 
0.0 -0.3008 0 2.0 1e-06 
0.0 -0.3007 0 2.0 1e-06 
0.0 -0.3006 0 2.0 1e-06 
0.0 -0.3005 0 2.0 1e-06 
0.0 -0.3004 0 2.0 1e-06 
0.0 -0.3003 0 2.0 1e-06 
0.0 -0.3002 0 2.0 1e-06 
0.0 -0.3001 0 2.0 1e-06 
0.0 -0.3 0 2.0 1e-06 
0.0 -0.2999 0 2.0 1e-06 
0.0 -0.2998 0 2.0 1e-06 
0.0 -0.2997 0 2.0 1e-06 
0.0 -0.2996 0 2.0 1e-06 
0.0 -0.2995 0 2.0 1e-06 
0.0 -0.2994 0 2.0 1e-06 
0.0 -0.2993 0 2.0 1e-06 
0.0 -0.2992 0 2.0 1e-06 
0.0 -0.2991 0 2.0 1e-06 
0.0 -0.299 0 2.0 1e-06 
0.0 -0.2989 0 2.0 1e-06 
0.0 -0.2988 0 2.0 1e-06 
0.0 -0.2987 0 2.0 1e-06 
0.0 -0.2986 0 2.0 1e-06 
0.0 -0.2985 0 2.0 1e-06 
0.0 -0.2984 0 2.0 1e-06 
0.0 -0.2983 0 2.0 1e-06 
0.0 -0.2982 0 2.0 1e-06 
0.0 -0.2981 0 2.0 1e-06 
0.0 -0.298 0 2.0 1e-06 
0.0 -0.2979 0 2.0 1e-06 
0.0 -0.2978 0 2.0 1e-06 
0.0 -0.2977 0 2.0 1e-06 
0.0 -0.2976 0 2.0 1e-06 
0.0 -0.2975 0 2.0 1e-06 
0.0 -0.2974 0 2.0 1e-06 
0.0 -0.2973 0 2.0 1e-06 
0.0 -0.2972 0 2.0 1e-06 
0.0 -0.2971 0 2.0 1e-06 
0.0 -0.297 0 2.0 1e-06 
0.0 -0.2969 0 2.0 1e-06 
0.0 -0.2968 0 2.0 1e-06 
0.0 -0.2967 0 2.0 1e-06 
0.0 -0.2966 0 2.0 1e-06 
0.0 -0.2965 0 2.0 1e-06 
0.0 -0.2964 0 2.0 1e-06 
0.0 -0.2963 0 2.0 1e-06 
0.0 -0.2962 0 2.0 1e-06 
0.0 -0.2961 0 2.0 1e-06 
0.0 -0.296 0 2.0 1e-06 
0.0 -0.2959 0 2.0 1e-06 
0.0 -0.2958 0 2.0 1e-06 
0.0 -0.2957 0 2.0 1e-06 
0.0 -0.2956 0 2.0 1e-06 
0.0 -0.2955 0 2.0 1e-06 
0.0 -0.2954 0 2.0 1e-06 
0.0 -0.2953 0 2.0 1e-06 
0.0 -0.2952 0 2.0 1e-06 
0.0 -0.2951 0 2.0 1e-06 
0.0 -0.295 0 2.0 1e-06 
0.0 -0.2949 0 2.0 1e-06 
0.0 -0.2948 0 2.0 1e-06 
0.0 -0.2947 0 2.0 1e-06 
0.0 -0.2946 0 2.0 1e-06 
0.0 -0.2945 0 2.0 1e-06 
0.0 -0.2944 0 2.0 1e-06 
0.0 -0.2943 0 2.0 1e-06 
0.0 -0.2942 0 2.0 1e-06 
0.0 -0.2941 0 2.0 1e-06 
0.0 -0.294 0 2.0 1e-06 
0.0 -0.2939 0 2.0 1e-06 
0.0 -0.2938 0 2.0 1e-06 
0.0 -0.2937 0 2.0 1e-06 
0.0 -0.2936 0 2.0 1e-06 
0.0 -0.2935 0 2.0 1e-06 
0.0 -0.2934 0 2.0 1e-06 
0.0 -0.2933 0 2.0 1e-06 
0.0 -0.2932 0 2.0 1e-06 
0.0 -0.2931 0 2.0 1e-06 
0.0 -0.293 0 2.0 1e-06 
0.0 -0.2929 0 2.0 1e-06 
0.0 -0.2928 0 2.0 1e-06 
0.0 -0.2927 0 2.0 1e-06 
0.0 -0.2926 0 2.0 1e-06 
0.0 -0.2925 0 2.0 1e-06 
0.0 -0.2924 0 2.0 1e-06 
0.0 -0.2923 0 2.0 1e-06 
0.0 -0.2922 0 2.0 1e-06 
0.0 -0.2921 0 2.0 1e-06 
0.0 -0.292 0 2.0 1e-06 
0.0 -0.2919 0 2.0 1e-06 
0.0 -0.2918 0 2.0 1e-06 
0.0 -0.2917 0 2.0 1e-06 
0.0 -0.2916 0 2.0 1e-06 
0.0 -0.2915 0 2.0 1e-06 
0.0 -0.2914 0 2.0 1e-06 
0.0 -0.2913 0 2.0 1e-06 
0.0 -0.2912 0 2.0 1e-06 
0.0 -0.2911 0 2.0 1e-06 
0.0 -0.291 0 2.0 1e-06 
0.0 -0.2909 0 2.0 1e-06 
0.0 -0.2908 0 2.0 1e-06 
0.0 -0.2907 0 2.0 1e-06 
0.0 -0.2906 0 2.0 1e-06 
0.0 -0.2905 0 2.0 1e-06 
0.0 -0.2904 0 2.0 1e-06 
0.0 -0.2903 0 2.0 1e-06 
0.0 -0.2902 0 2.0 1e-06 
0.0 -0.2901 0 2.0 1e-06 
0.0 -0.29 0 2.0 1e-06 
0.0 -0.2899 0 2.0 1e-06 
0.0 -0.2898 0 2.0 1e-06 
0.0 -0.2897 0 2.0 1e-06 
0.0 -0.2896 0 2.0 1e-06 
0.0 -0.2895 0 2.0 1e-06 
0.0 -0.2894 0 2.0 1e-06 
0.0 -0.2893 0 2.0 1e-06 
0.0 -0.2892 0 2.0 1e-06 
0.0 -0.2891 0 2.0 1e-06 
0.0 -0.289 0 2.0 1e-06 
0.0 -0.2889 0 2.0 1e-06 
0.0 -0.2888 0 2.0 1e-06 
0.0 -0.2887 0 2.0 1e-06 
0.0 -0.2886 0 2.0 1e-06 
0.0 -0.2885 0 2.0 1e-06 
0.0 -0.2884 0 2.0 1e-06 
0.0 -0.2883 0 2.0 1e-06 
0.0 -0.2882 0 2.0 1e-06 
0.0 -0.2881 0 2.0 1e-06 
0.0 -0.288 0 2.0 1e-06 
0.0 -0.2879 0 2.0 1e-06 
0.0 -0.2878 0 2.0 1e-06 
0.0 -0.2877 0 2.0 1e-06 
0.0 -0.2876 0 2.0 1e-06 
0.0 -0.2875 0 2.0 1e-06 
0.0 -0.2874 0 2.0 1e-06 
0.0 -0.2873 0 2.0 1e-06 
0.0 -0.2872 0 2.0 1e-06 
0.0 -0.2871 0 2.0 1e-06 
0.0 -0.287 0 2.0 1e-06 
0.0 -0.2869 0 2.0 1e-06 
0.0 -0.2868 0 2.0 1e-06 
0.0 -0.2867 0 2.0 1e-06 
0.0 -0.2866 0 2.0 1e-06 
0.0 -0.2865 0 2.0 1e-06 
0.0 -0.2864 0 2.0 1e-06 
0.0 -0.2863 0 2.0 1e-06 
0.0 -0.2862 0 2.0 1e-06 
0.0 -0.2861 0 2.0 1e-06 
0.0 -0.286 0 2.0 1e-06 
0.0 -0.2859 0 2.0 1e-06 
0.0 -0.2858 0 2.0 1e-06 
0.0 -0.2857 0 2.0 1e-06 
0.0 -0.2856 0 2.0 1e-06 
0.0 -0.2855 0 2.0 1e-06 
0.0 -0.2854 0 2.0 1e-06 
0.0 -0.2853 0 2.0 1e-06 
0.0 -0.2852 0 2.0 1e-06 
0.0 -0.2851 0 2.0 1e-06 
0.0 -0.285 0 2.0 1e-06 
0.0 -0.2849 0 2.0 1e-06 
0.0 -0.2848 0 2.0 1e-06 
0.0 -0.2847 0 2.0 1e-06 
0.0 -0.2846 0 2.0 1e-06 
0.0 -0.2845 0 2.0 1e-06 
0.0 -0.2844 0 2.0 1e-06 
0.0 -0.2843 0 2.0 1e-06 
0.0 -0.2842 0 2.0 1e-06 
0.0 -0.2841 0 2.0 1e-06 
0.0 -0.284 0 2.0 1e-06 
0.0 -0.2839 0 2.0 1e-06 
0.0 -0.2838 0 2.0 1e-06 
0.0 -0.2837 0 2.0 1e-06 
0.0 -0.2836 0 2.0 1e-06 
0.0 -0.2835 0 2.0 1e-06 
0.0 -0.2834 0 2.0 1e-06 
0.0 -0.2833 0 2.0 1e-06 
0.0 -0.2832 0 2.0 1e-06 
0.0 -0.2831 0 2.0 1e-06 
0.0 -0.283 0 2.0 1e-06 
0.0 -0.2829 0 2.0 1e-06 
0.0 -0.2828 0 2.0 1e-06 
0.0 -0.2827 0 2.0 1e-06 
0.0 -0.2826 0 2.0 1e-06 
0.0 -0.2825 0 2.0 1e-06 
0.0 -0.2824 0 2.0 1e-06 
0.0 -0.2823 0 2.0 1e-06 
0.0 -0.2822 0 2.0 1e-06 
0.0 -0.2821 0 2.0 1e-06 
0.0 -0.282 0 2.0 1e-06 
0.0 -0.2819 0 2.0 1e-06 
0.0 -0.2818 0 2.0 1e-06 
0.0 -0.2817 0 2.0 1e-06 
0.0 -0.2816 0 2.0 1e-06 
0.0 -0.2815 0 2.0 1e-06 
0.0 -0.2814 0 2.0 1e-06 
0.0 -0.2813 0 2.0 1e-06 
0.0 -0.2812 0 2.0 1e-06 
0.0 -0.2811 0 2.0 1e-06 
0.0 -0.281 0 2.0 1e-06 
0.0 -0.2809 0 2.0 1e-06 
0.0 -0.2808 0 2.0 1e-06 
0.0 -0.2807 0 2.0 1e-06 
0.0 -0.2806 0 2.0 1e-06 
0.0 -0.2805 0 2.0 1e-06 
0.0 -0.2804 0 2.0 1e-06 
0.0 -0.2803 0 2.0 1e-06 
0.0 -0.2802 0 2.0 1e-06 
0.0 -0.2801 0 2.0 1e-06 
0.0 -0.28 0 2.0 1e-06 
0.0 -0.2799 0 2.0 1e-06 
0.0 -0.2798 0 2.0 1e-06 
0.0 -0.2797 0 2.0 1e-06 
0.0 -0.2796 0 2.0 1e-06 
0.0 -0.2795 0 2.0 1e-06 
0.0 -0.2794 0 2.0 1e-06 
0.0 -0.2793 0 2.0 1e-06 
0.0 -0.2792 0 2.0 1e-06 
0.0 -0.2791 0 2.0 1e-06 
0.0 -0.279 0 2.0 1e-06 
0.0 -0.2789 0 2.0 1e-06 
0.0 -0.2788 0 2.0 1e-06 
0.0 -0.2787 0 2.0 1e-06 
0.0 -0.2786 0 2.0 1e-06 
0.0 -0.2785 0 2.0 1e-06 
0.0 -0.2784 0 2.0 1e-06 
0.0 -0.2783 0 2.0 1e-06 
0.0 -0.2782 0 2.0 1e-06 
0.0 -0.2781 0 2.0 1e-06 
0.0 -0.278 0 2.0 1e-06 
0.0 -0.2779 0 2.0 1e-06 
0.0 -0.2778 0 2.0 1e-06 
0.0 -0.2777 0 2.0 1e-06 
0.0 -0.2776 0 2.0 1e-06 
0.0 -0.2775 0 2.0 1e-06 
0.0 -0.2774 0 2.0 1e-06 
0.0 -0.2773 0 2.0 1e-06 
0.0 -0.2772 0 2.0 1e-06 
0.0 -0.2771 0 2.0 1e-06 
0.0 -0.277 0 2.0 1e-06 
0.0 -0.2769 0 2.0 1e-06 
0.0 -0.2768 0 2.0 1e-06 
0.0 -0.2767 0 2.0 1e-06 
0.0 -0.2766 0 2.0 1e-06 
0.0 -0.2765 0 2.0 1e-06 
0.0 -0.2764 0 2.0 1e-06 
0.0 -0.2763 0 2.0 1e-06 
0.0 -0.2762 0 2.0 1e-06 
0.0 -0.2761 0 2.0 1e-06 
0.0 -0.276 0 2.0 1e-06 
0.0 -0.2759 0 2.0 1e-06 
0.0 -0.2758 0 2.0 1e-06 
0.0 -0.2757 0 2.0 1e-06 
0.0 -0.2756 0 2.0 1e-06 
0.0 -0.2755 0 2.0 1e-06 
0.0 -0.2754 0 2.0 1e-06 
0.0 -0.2753 0 2.0 1e-06 
0.0 -0.2752 0 2.0 1e-06 
0.0 -0.2751 0 2.0 1e-06 
0.0 -0.275 0 2.0 1e-06 
0.0 -0.2749 0 2.0 1e-06 
0.0 -0.2748 0 2.0 1e-06 
0.0 -0.2747 0 2.0 1e-06 
0.0 -0.2746 0 2.0 1e-06 
0.0 -0.2745 0 2.0 1e-06 
0.0 -0.2744 0 2.0 1e-06 
0.0 -0.2743 0 2.0 1e-06 
0.0 -0.2742 0 2.0 1e-06 
0.0 -0.2741 0 2.0 1e-06 
0.0 -0.274 0 2.0 1e-06 
0.0 -0.2739 0 2.0 1e-06 
0.0 -0.2738 0 2.0 1e-06 
0.0 -0.2737 0 2.0 1e-06 
0.0 -0.2736 0 2.0 1e-06 
0.0 -0.2735 0 2.0 1e-06 
0.0 -0.2734 0 2.0 1e-06 
0.0 -0.2733 0 2.0 1e-06 
0.0 -0.2732 0 2.0 1e-06 
0.0 -0.2731 0 2.0 1e-06 
0.0 -0.273 0 2.0 1e-06 
0.0 -0.2729 0 2.0 1e-06 
0.0 -0.2728 0 2.0 1e-06 
0.0 -0.2727 0 2.0 1e-06 
0.0 -0.2726 0 2.0 1e-06 
0.0 -0.2725 0 2.0 1e-06 
0.0 -0.2724 0 2.0 1e-06 
0.0 -0.2723 0 2.0 1e-06 
0.0 -0.2722 0 2.0 1e-06 
0.0 -0.2721 0 2.0 1e-06 
0.0 -0.272 0 2.0 1e-06 
0.0 -0.2719 0 2.0 1e-06 
0.0 -0.2718 0 2.0 1e-06 
0.0 -0.2717 0 2.0 1e-06 
0.0 -0.2716 0 2.0 1e-06 
0.0 -0.2715 0 2.0 1e-06 
0.0 -0.2714 0 2.0 1e-06 
0.0 -0.2713 0 2.0 1e-06 
0.0 -0.2712 0 2.0 1e-06 
0.0 -0.2711 0 2.0 1e-06 
0.0 -0.271 0 2.0 1e-06 
0.0 -0.2709 0 2.0 1e-06 
0.0 -0.2708 0 2.0 1e-06 
0.0 -0.2707 0 2.0 1e-06 
0.0 -0.2706 0 2.0 1e-06 
0.0 -0.2705 0 2.0 1e-06 
0.0 -0.2704 0 2.0 1e-06 
0.0 -0.2703 0 2.0 1e-06 
0.0 -0.2702 0 2.0 1e-06 
0.0 -0.2701 0 2.0 1e-06 
0.0 -0.27 0 2.0 1e-06 
0.0 -0.2699 0 2.0 1e-06 
0.0 -0.2698 0 2.0 1e-06 
0.0 -0.2697 0 2.0 1e-06 
0.0 -0.2696 0 2.0 1e-06 
0.0 -0.2695 0 2.0 1e-06 
0.0 -0.2694 0 2.0 1e-06 
0.0 -0.2693 0 2.0 1e-06 
0.0 -0.2692 0 2.0 1e-06 
0.0 -0.2691 0 2.0 1e-06 
0.0 -0.269 0 2.0 1e-06 
0.0 -0.2689 0 2.0 1e-06 
0.0 -0.2688 0 2.0 1e-06 
0.0 -0.2687 0 2.0 1e-06 
0.0 -0.2686 0 2.0 1e-06 
0.0 -0.2685 0 2.0 1e-06 
0.0 -0.2684 0 2.0 1e-06 
0.0 -0.2683 0 2.0 1e-06 
0.0 -0.2682 0 2.0 1e-06 
0.0 -0.2681 0 2.0 1e-06 
0.0 -0.268 0 2.0 1e-06 
0.0 -0.2679 0 2.0 1e-06 
0.0 -0.2678 0 2.0 1e-06 
0.0 -0.2677 0 2.0 1e-06 
0.0 -0.2676 0 2.0 1e-06 
0.0 -0.2675 0 2.0 1e-06 
0.0 -0.2674 0 2.0 1e-06 
0.0 -0.2673 0 2.0 1e-06 
0.0 -0.2672 0 2.0 1e-06 
0.0 -0.2671 0 2.0 1e-06 
0.0 -0.267 0 2.0 1e-06 
0.0 -0.2669 0 2.0 1e-06 
0.0 -0.2668 0 2.0 1e-06 
0.0 -0.2667 0 2.0 1e-06 
0.0 -0.2666 0 2.0 1e-06 
0.0 -0.2665 0 2.0 1e-06 
0.0 -0.2664 0 2.0 1e-06 
0.0 -0.2663 0 2.0 1e-06 
0.0 -0.2662 0 2.0 1e-06 
0.0 -0.2661 0 2.0 1e-06 
0.0 -0.266 0 2.0 1e-06 
0.0 -0.2659 0 2.0 1e-06 
0.0 -0.2658 0 2.0 1e-06 
0.0 -0.2657 0 2.0 1e-06 
0.0 -0.2656 0 2.0 1e-06 
0.0 -0.2655 0 2.0 1e-06 
0.0 -0.2654 0 2.0 1e-06 
0.0 -0.2653 0 2.0 1e-06 
0.0 -0.2652 0 2.0 1e-06 
0.0 -0.2651 0 2.0 1e-06 
0.0 -0.265 0 2.0 1e-06 
0.0 -0.2649 0 2.0 1e-06 
0.0 -0.2648 0 2.0 1e-06 
0.0 -0.2647 0 2.0 1e-06 
0.0 -0.2646 0 2.0 1e-06 
0.0 -0.2645 0 2.0 1e-06 
0.0 -0.2644 0 2.0 1e-06 
0.0 -0.2643 0 2.0 1e-06 
0.0 -0.2642 0 2.0 1e-06 
0.0 -0.2641 0 2.0 1e-06 
0.0 -0.264 0 2.0 1e-06 
0.0 -0.2639 0 2.0 1e-06 
0.0 -0.2638 0 2.0 1e-06 
0.0 -0.2637 0 2.0 1e-06 
0.0 -0.2636 0 2.0 1e-06 
0.0 -0.2635 0 2.0 1e-06 
0.0 -0.2634 0 2.0 1e-06 
0.0 -0.2633 0 2.0 1e-06 
0.0 -0.2632 0 2.0 1e-06 
0.0 -0.2631 0 2.0 1e-06 
0.0 -0.263 0 2.0 1e-06 
0.0 -0.2629 0 2.0 1e-06 
0.0 -0.2628 0 2.0 1e-06 
0.0 -0.2627 0 2.0 1e-06 
0.0 -0.2626 0 2.0 1e-06 
0.0 -0.2625 0 2.0 1e-06 
0.0 -0.2624 0 2.0 1e-06 
0.0 -0.2623 0 2.0 1e-06 
0.0 -0.2622 0 2.0 1e-06 
0.0 -0.2621 0 2.0 1e-06 
0.0 -0.262 0 2.0 1e-06 
0.0 -0.2619 0 2.0 1e-06 
0.0 -0.2618 0 2.0 1e-06 
0.0 -0.2617 0 2.0 1e-06 
0.0 -0.2616 0 2.0 1e-06 
0.0 -0.2615 0 2.0 1e-06 
0.0 -0.2614 0 2.0 1e-06 
0.0 -0.2613 0 2.0 1e-06 
0.0 -0.2612 0 2.0 1e-06 
0.0 -0.2611 0 2.0 1e-06 
0.0 -0.261 0 2.0 1e-06 
0.0 -0.2609 0 2.0 1e-06 
0.0 -0.2608 0 2.0 1e-06 
0.0 -0.2607 0 2.0 1e-06 
0.0 -0.2606 0 2.0 1e-06 
0.0 -0.2605 0 2.0 1e-06 
0.0 -0.2604 0 2.0 1e-06 
0.0 -0.2603 0 2.0 1e-06 
0.0 -0.2602 0 2.0 1e-06 
0.0 -0.2601 0 2.0 1e-06 
0.0 -0.26 0 2.0 1e-06 
0.0 -0.2599 0 2.0 1e-06 
0.0 -0.2598 0 2.0 1e-06 
0.0 -0.2597 0 2.0 1e-06 
0.0 -0.2596 0 2.0 1e-06 
0.0 -0.2595 0 2.0 1e-06 
0.0 -0.2594 0 2.0 1e-06 
0.0 -0.2593 0 2.0 1e-06 
0.0 -0.2592 0 2.0 1e-06 
0.0 -0.2591 0 2.0 1e-06 
0.0 -0.259 0 2.0 1e-06 
0.0 -0.2589 0 2.0 1e-06 
0.0 -0.2588 0 2.0 1e-06 
0.0 -0.2587 0 2.0 1e-06 
0.0 -0.2586 0 2.0 1e-06 
0.0 -0.2585 0 2.0 1e-06 
0.0 -0.2584 0 2.0 1e-06 
0.0 -0.2583 0 2.0 1e-06 
0.0 -0.2582 0 2.0 1e-06 
0.0 -0.2581 0 2.0 1e-06 
0.0 -0.258 0 2.0 1e-06 
0.0 -0.2579 0 2.0 1e-06 
0.0 -0.2578 0 2.0 1e-06 
0.0 -0.2577 0 2.0 1e-06 
0.0 -0.2576 0 2.0 1e-06 
0.0 -0.2575 0 2.0 1e-06 
0.0 -0.2574 0 2.0 1e-06 
0.0 -0.2573 0 2.0 1e-06 
0.0 -0.2572 0 2.0 1e-06 
0.0 -0.2571 0 2.0 1e-06 
0.0 -0.257 0 2.0 1e-06 
0.0 -0.2569 0 2.0 1e-06 
0.0 -0.2568 0 2.0 1e-06 
0.0 -0.2567 0 2.0 1e-06 
0.0 -0.2566 0 2.0 1e-06 
0.0 -0.2565 0 2.0 1e-06 
0.0 -0.2564 0 2.0 1e-06 
0.0 -0.2563 0 2.0 1e-06 
0.0 -0.2562 0 2.0 1e-06 
0.0 -0.2561 0 2.0 1e-06 
0.0 -0.256 0 2.0 1e-06 
0.0 -0.2559 0 2.0 1e-06 
0.0 -0.2558 0 2.0 1e-06 
0.0 -0.2557 0 2.0 1e-06 
0.0 -0.2556 0 2.0 1e-06 
0.0 -0.2555 0 2.0 1e-06 
0.0 -0.2554 0 2.0 1e-06 
0.0 -0.2553 0 2.0 1e-06 
0.0 -0.2552 0 2.0 1e-06 
0.0 -0.2551 0 2.0 1e-06 
0.0 -0.255 0 2.0 1e-06 
0.0 -0.2549 0 2.0 1e-06 
0.0 -0.2548 0 2.0 1e-06 
0.0 -0.2547 0 2.0 1e-06 
0.0 -0.2546 0 2.0 1e-06 
0.0 -0.2545 0 2.0 1e-06 
0.0 -0.2544 0 2.0 1e-06 
0.0 -0.2543 0 2.0 1e-06 
0.0 -0.2542 0 2.0 1e-06 
0.0 -0.2541 0 2.0 1e-06 
0.0 -0.254 0 2.0 1e-06 
0.0 -0.2539 0 2.0 1e-06 
0.0 -0.2538 0 2.0 1e-06 
0.0 -0.2537 0 2.0 1e-06 
0.0 -0.2536 0 2.0 1e-06 
0.0 -0.2535 0 2.0 1e-06 
0.0 -0.2534 0 2.0 1e-06 
0.0 -0.2533 0 2.0 1e-06 
0.0 -0.2532 0 2.0 1e-06 
0.0 -0.2531 0 2.0 1e-06 
0.0 -0.253 0 2.0 1e-06 
0.0 -0.2529 0 2.0 1e-06 
0.0 -0.2528 0 2.0 1e-06 
0.0 -0.2527 0 2.0 1e-06 
0.0 -0.2526 0 2.0 1e-06 
0.0 -0.2525 0 2.0 1e-06 
0.0 -0.2524 0 2.0 1e-06 
0.0 -0.2523 0 2.0 1e-06 
0.0 -0.2522 0 2.0 1e-06 
0.0 -0.2521 0 2.0 1e-06 
0.0 -0.252 0 2.0 1e-06 
0.0 -0.2519 0 2.0 1e-06 
0.0 -0.2518 0 2.0 1e-06 
0.0 -0.2517 0 2.0 1e-06 
0.0 -0.2516 0 2.0 1e-06 
0.0 -0.2515 0 2.0 1e-06 
0.0 -0.2514 0 2.0 1e-06 
0.0 -0.2513 0 2.0 1e-06 
0.0 -0.2512 0 2.0 1e-06 
0.0 -0.2511 0 2.0 1e-06 
0.0 -0.251 0 2.0 1e-06 
0.0 -0.2509 0 2.0 1e-06 
0.0 -0.2508 0 2.0 1e-06 
0.0 -0.2507 0 2.0 1e-06 
0.0 -0.2506 0 2.0 1e-06 
0.0 -0.2505 0 2.0 1e-06 
0.0 -0.2504 0 2.0 1e-06 
0.0 -0.2503 0 2.0 1e-06 
0.0 -0.2502 0 2.0 1e-06 
0.0 -0.2501 0 2.0 1e-06 
0.0 -0.25 0 2.0 1e-06 
0.0 -0.2499 0 2.0 1e-06 
0.0 -0.2498 0 2.0 1e-06 
0.0 -0.2497 0 2.0 1e-06 
0.0 -0.2496 0 2.0 1e-06 
0.0 -0.2495 0 2.0 1e-06 
0.0 -0.2494 0 2.0 1e-06 
0.0 -0.2493 0 2.0 1e-06 
0.0 -0.2492 0 2.0 1e-06 
0.0 -0.2491 0 2.0 1e-06 
0.0 -0.249 0 2.0 1e-06 
0.0 -0.2489 0 2.0 1e-06 
0.0 -0.2488 0 2.0 1e-06 
0.0 -0.2487 0 2.0 1e-06 
0.0 -0.2486 0 2.0 1e-06 
0.0 -0.2485 0 2.0 1e-06 
0.0 -0.2484 0 2.0 1e-06 
0.0 -0.2483 0 2.0 1e-06 
0.0 -0.2482 0 2.0 1e-06 
0.0 -0.2481 0 2.0 1e-06 
0.0 -0.248 0 2.0 1e-06 
0.0 -0.2479 0 2.0 1e-06 
0.0 -0.2478 0 2.0 1e-06 
0.0 -0.2477 0 2.0 1e-06 
0.0 -0.2476 0 2.0 1e-06 
0.0 -0.2475 0 2.0 1e-06 
0.0 -0.2474 0 2.0 1e-06 
0.0 -0.2473 0 2.0 1e-06 
0.0 -0.2472 0 2.0 1e-06 
0.0 -0.2471 0 2.0 1e-06 
0.0 -0.247 0 2.0 1e-06 
0.0 -0.2469 0 2.0 1e-06 
0.0 -0.2468 0 2.0 1e-06 
0.0 -0.2467 0 2.0 1e-06 
0.0 -0.2466 0 2.0 1e-06 
0.0 -0.2465 0 2.0 1e-06 
0.0 -0.2464 0 2.0 1e-06 
0.0 -0.2463 0 2.0 1e-06 
0.0 -0.2462 0 2.0 1e-06 
0.0 -0.2461 0 2.0 1e-06 
0.0 -0.246 0 2.0 1e-06 
0.0 -0.2459 0 2.0 1e-06 
0.0 -0.2458 0 2.0 1e-06 
0.0 -0.2457 0 2.0 1e-06 
0.0 -0.2456 0 2.0 1e-06 
0.0 -0.2455 0 2.0 1e-06 
0.0 -0.2454 0 2.0 1e-06 
0.0 -0.2453 0 2.0 1e-06 
0.0 -0.2452 0 2.0 1e-06 
0.0 -0.2451 0 2.0 1e-06 
0.0 -0.245 0 2.0 1e-06 
0.0 -0.2449 0 2.0 1e-06 
0.0 -0.2448 0 2.0 1e-06 
0.0 -0.2447 0 2.0 1e-06 
0.0 -0.2446 0 2.0 1e-06 
0.0 -0.2445 0 2.0 1e-06 
0.0 -0.2444 0 2.0 1e-06 
0.0 -0.2443 0 2.0 1e-06 
0.0 -0.2442 0 2.0 1e-06 
0.0 -0.2441 0 2.0 1e-06 
0.0 -0.244 0 2.0 1e-06 
0.0 -0.2439 0 2.0 1e-06 
0.0 -0.2438 0 2.0 1e-06 
0.0 -0.2437 0 2.0 1e-06 
0.0 -0.2436 0 2.0 1e-06 
0.0 -0.2435 0 2.0 1e-06 
0.0 -0.2434 0 2.0 1e-06 
0.0 -0.2433 0 2.0 1e-06 
0.0 -0.2432 0 2.0 1e-06 
0.0 -0.2431 0 2.0 1e-06 
0.0 -0.243 0 2.0 1e-06 
0.0 -0.2429 0 2.0 1e-06 
0.0 -0.2428 0 2.0 1e-06 
0.0 -0.2427 0 2.0 1e-06 
0.0 -0.2426 0 2.0 1e-06 
0.0 -0.2425 0 2.0 1e-06 
0.0 -0.2424 0 2.0 1e-06 
0.0 -0.2423 0 2.0 1e-06 
0.0 -0.2422 0 2.0 1e-06 
0.0 -0.2421 0 2.0 1e-06 
0.0 -0.242 0 2.0 1e-06 
0.0 -0.2419 0 2.0 1e-06 
0.0 -0.2418 0 2.0 1e-06 
0.0 -0.2417 0 2.0 1e-06 
0.0 -0.2416 0 2.0 1e-06 
0.0 -0.2415 0 2.0 1e-06 
0.0 -0.2414 0 2.0 1e-06 
0.0 -0.2413 0 2.0 1e-06 
0.0 -0.2412 0 2.0 1e-06 
0.0 -0.2411 0 2.0 1e-06 
0.0 -0.241 0 2.0 1e-06 
0.0 -0.2409 0 2.0 1e-06 
0.0 -0.2408 0 2.0 1e-06 
0.0 -0.2407 0 2.0 1e-06 
0.0 -0.2406 0 2.0 1e-06 
0.0 -0.2405 0 2.0 1e-06 
0.0 -0.2404 0 2.0 1e-06 
0.0 -0.2403 0 2.0 1e-06 
0.0 -0.2402 0 2.0 1e-06 
0.0 -0.2401 0 2.0 1e-06 
0.0 -0.24 0 2.0 1e-06 
0.0 -0.2399 0 2.0 1e-06 
0.0 -0.2398 0 2.0 1e-06 
0.0 -0.2397 0 2.0 1e-06 
0.0 -0.2396 0 2.0 1e-06 
0.0 -0.2395 0 2.0 1e-06 
0.0 -0.2394 0 2.0 1e-06 
0.0 -0.2393 0 2.0 1e-06 
0.0 -0.2392 0 2.0 1e-06 
0.0 -0.2391 0 2.0 1e-06 
0.0 -0.239 0 2.0 1e-06 
0.0 -0.2389 0 2.0 1e-06 
0.0 -0.2388 0 2.0 1e-06 
0.0 -0.2387 0 2.0 1e-06 
0.0 -0.2386 0 2.0 1e-06 
0.0 -0.2385 0 2.0 1e-06 
0.0 -0.2384 0 2.0 1e-06 
0.0 -0.2383 0 2.0 1e-06 
0.0 -0.2382 0 2.0 1e-06 
0.0 -0.2381 0 2.0 1e-06 
0.0 -0.238 0 2.0 1e-06 
0.0 -0.2379 0 2.0 1e-06 
0.0 -0.2378 0 2.0 1e-06 
0.0 -0.2377 0 2.0 1e-06 
0.0 -0.2376 0 2.0 1e-06 
0.0 -0.2375 0 2.0 1e-06 
0.0 -0.2374 0 2.0 1e-06 
0.0 -0.2373 0 2.0 1e-06 
0.0 -0.2372 0 2.0 1e-06 
0.0 -0.2371 0 2.0 1e-06 
0.0 -0.237 0 2.0 1e-06 
0.0 -0.2369 0 2.0 1e-06 
0.0 -0.2368 0 2.0 1e-06 
0.0 -0.2367 0 2.0 1e-06 
0.0 -0.2366 0 2.0 1e-06 
0.0 -0.2365 0 2.0 1e-06 
0.0 -0.2364 0 2.0 1e-06 
0.0 -0.2363 0 2.0 1e-06 
0.0 -0.2362 0 2.0 1e-06 
0.0 -0.2361 0 2.0 1e-06 
0.0 -0.236 0 2.0 1e-06 
0.0 -0.2359 0 2.0 1e-06 
0.0 -0.2358 0 2.0 1e-06 
0.0 -0.2357 0 2.0 1e-06 
0.0 -0.2356 0 2.0 1e-06 
0.0 -0.2355 0 2.0 1e-06 
0.0 -0.2354 0 2.0 1e-06 
0.0 -0.2353 0 2.0 1e-06 
0.0 -0.2352 0 2.0 1e-06 
0.0 -0.2351 0 2.0 1e-06 
0.0 -0.235 0 2.0 1e-06 
0.0 -0.2349 0 2.0 1e-06 
0.0 -0.2348 0 2.0 1e-06 
0.0 -0.2347 0 2.0 1e-06 
0.0 -0.2346 0 2.0 1e-06 
0.0 -0.2345 0 2.0 1e-06 
0.0 -0.2344 0 2.0 1e-06 
0.0 -0.2343 0 2.0 1e-06 
0.0 -0.2342 0 2.0 1e-06 
0.0 -0.2341 0 2.0 1e-06 
0.0 -0.234 0 2.0 1e-06 
0.0 -0.2339 0 2.0 1e-06 
0.0 -0.2338 0 2.0 1e-06 
0.0 -0.2337 0 2.0 1e-06 
0.0 -0.2336 0 2.0 1e-06 
0.0 -0.2335 0 2.0 1e-06 
0.0 -0.2334 0 2.0 1e-06 
0.0 -0.2333 0 2.0 1e-06 
0.0 -0.2332 0 2.0 1e-06 
0.0 -0.2331 0 2.0 1e-06 
0.0 -0.233 0 2.0 1e-06 
0.0 -0.2329 0 2.0 1e-06 
0.0 -0.2328 0 2.0 1e-06 
0.0 -0.2327 0 2.0 1e-06 
0.0 -0.2326 0 2.0 1e-06 
0.0 -0.2325 0 2.0 1e-06 
0.0 -0.2324 0 2.0 1e-06 
0.0 -0.2323 0 2.0 1e-06 
0.0 -0.2322 0 2.0 1e-06 
0.0 -0.2321 0 2.0 1e-06 
0.0 -0.232 0 2.0 1e-06 
0.0 -0.2319 0 2.0 1e-06 
0.0 -0.2318 0 2.0 1e-06 
0.0 -0.2317 0 2.0 1e-06 
0.0 -0.2316 0 2.0 1e-06 
0.0 -0.2315 0 2.0 1e-06 
0.0 -0.2314 0 2.0 1e-06 
0.0 -0.2313 0 2.0 1e-06 
0.0 -0.2312 0 2.0 1e-06 
0.0 -0.2311 0 2.0 1e-06 
0.0 -0.231 0 2.0 1e-06 
0.0 -0.2309 0 2.0 1e-06 
0.0 -0.2308 0 2.0 1e-06 
0.0 -0.2307 0 2.0 1e-06 
0.0 -0.2306 0 2.0 1e-06 
0.0 -0.2305 0 2.0 1e-06 
0.0 -0.2304 0 2.0 1e-06 
0.0 -0.2303 0 2.0 1e-06 
0.0 -0.2302 0 2.0 1e-06 
0.0 -0.2301 0 2.0 1e-06 
0.0 -0.23 0 2.0 1e-06 
0.0 -0.2299 0 2.0 1e-06 
0.0 -0.2298 0 2.0 1e-06 
0.0 -0.2297 0 2.0 1e-06 
0.0 -0.2296 0 2.0 1e-06 
0.0 -0.2295 0 2.0 1e-06 
0.0 -0.2294 0 2.0 1e-06 
0.0 -0.2293 0 2.0 1e-06 
0.0 -0.2292 0 2.0 1e-06 
0.0 -0.2291 0 2.0 1e-06 
0.0 -0.229 0 2.0 1e-06 
0.0 -0.2289 0 2.0 1e-06 
0.0 -0.2288 0 2.0 1e-06 
0.0 -0.2287 0 2.0 1e-06 
0.0 -0.2286 0 2.0 1e-06 
0.0 -0.2285 0 2.0 1e-06 
0.0 -0.2284 0 2.0 1e-06 
0.0 -0.2283 0 2.0 1e-06 
0.0 -0.2282 0 2.0 1e-06 
0.0 -0.2281 0 2.0 1e-06 
0.0 -0.228 0 2.0 1e-06 
0.0 -0.2279 0 2.0 1e-06 
0.0 -0.2278 0 2.0 1e-06 
0.0 -0.2277 0 2.0 1e-06 
0.0 -0.2276 0 2.0 1e-06 
0.0 -0.2275 0 2.0 1e-06 
0.0 -0.2274 0 2.0 1e-06 
0.0 -0.2273 0 2.0 1e-06 
0.0 -0.2272 0 2.0 1e-06 
0.0 -0.2271 0 2.0 1e-06 
0.0 -0.227 0 2.0 1e-06 
0.0 -0.2269 0 2.0 1e-06 
0.0 -0.2268 0 2.0 1e-06 
0.0 -0.2267 0 2.0 1e-06 
0.0 -0.2266 0 2.0 1e-06 
0.0 -0.2265 0 2.0 1e-06 
0.0 -0.2264 0 2.0 1e-06 
0.0 -0.2263 0 2.0 1e-06 
0.0 -0.2262 0 2.0 1e-06 
0.0 -0.2261 0 2.0 1e-06 
0.0 -0.226 0 2.0 1e-06 
0.0 -0.2259 0 2.0 1e-06 
0.0 -0.2258 0 2.0 1e-06 
0.0 -0.2257 0 2.0 1e-06 
0.0 -0.2256 0 2.0 1e-06 
0.0 -0.2255 0 2.0 1e-06 
0.0 -0.2254 0 2.0 1e-06 
0.0 -0.2253 0 2.0 1e-06 
0.0 -0.2252 0 2.0 1e-06 
0.0 -0.2251 0 2.0 1e-06 
0.0 -0.225 0 2.0 1e-06 
0.0 -0.2249 0 2.0 1e-06 
0.0 -0.2248 0 2.0 1e-06 
0.0 -0.2247 0 2.0 1e-06 
0.0 -0.2246 0 2.0 1e-06 
0.0 -0.2245 0 2.0 1e-06 
0.0 -0.2244 0 2.0 1e-06 
0.0 -0.2243 0 2.0 1e-06 
0.0 -0.2242 0 2.0 1e-06 
0.0 -0.2241 0 2.0 1e-06 
0.0 -0.224 0 2.0 1e-06 
0.0 -0.2239 0 2.0 1e-06 
0.0 -0.2238 0 2.0 1e-06 
0.0 -0.2237 0 2.0 1e-06 
0.0 -0.2236 0 2.0 1e-06 
0.0 -0.2235 0 2.0 1e-06 
0.0 -0.2234 0 2.0 1e-06 
0.0 -0.2233 0 2.0 1e-06 
0.0 -0.2232 0 2.0 1e-06 
0.0 -0.2231 0 2.0 1e-06 
0.0 -0.223 0 2.0 1e-06 
0.0 -0.2229 0 2.0 1e-06 
0.0 -0.2228 0 2.0 1e-06 
0.0 -0.2227 0 2.0 1e-06 
0.0 -0.2226 0 2.0 1e-06 
0.0 -0.2225 0 2.0 1e-06 
0.0 -0.2224 0 2.0 1e-06 
0.0 -0.2223 0 2.0 1e-06 
0.0 -0.2222 0 2.0 1e-06 
0.0 -0.2221 0 2.0 1e-06 
0.0 -0.222 0 2.0 1e-06 
0.0 -0.2219 0 2.0 1e-06 
0.0 -0.2218 0 2.0 1e-06 
0.0 -0.2217 0 2.0 1e-06 
0.0 -0.2216 0 2.0 1e-06 
0.0 -0.2215 0 2.0 1e-06 
0.0 -0.2214 0 2.0 1e-06 
0.0 -0.2213 0 2.0 1e-06 
0.0 -0.2212 0 2.0 1e-06 
0.0 -0.2211 0 2.0 1e-06 
0.0 -0.221 0 2.0 1e-06 
0.0 -0.2209 0 2.0 1e-06 
0.0 -0.2208 0 2.0 1e-06 
0.0 -0.2207 0 2.0 1e-06 
0.0 -0.2206 0 2.0 1e-06 
0.0 -0.2205 0 2.0 1e-06 
0.0 -0.2204 0 2.0 1e-06 
0.0 -0.2203 0 2.0 1e-06 
0.0 -0.2202 0 2.0 1e-06 
0.0 -0.2201 0 2.0 1e-06 
0.0 -0.22 0 2.0 1e-06 
0.0 -0.2199 0 2.0 1e-06 
0.0 -0.2198 0 2.0 1e-06 
0.0 -0.2197 0 2.0 1e-06 
0.0 -0.2196 0 2.0 1e-06 
0.0 -0.2195 0 2.0 1e-06 
0.0 -0.2194 0 2.0 1e-06 
0.0 -0.2193 0 2.0 1e-06 
0.0 -0.2192 0 2.0 1e-06 
0.0 -0.2191 0 2.0 1e-06 
0.0 -0.219 0 2.0 1e-06 
0.0 -0.2189 0 2.0 1e-06 
0.0 -0.2188 0 2.0 1e-06 
0.0 -0.2187 0 2.0 1e-06 
0.0 -0.2186 0 2.0 1e-06 
0.0 -0.2185 0 2.0 1e-06 
0.0 -0.2184 0 2.0 1e-06 
0.0 -0.2183 0 2.0 1e-06 
0.0 -0.2182 0 2.0 1e-06 
0.0 -0.2181 0 2.0 1e-06 
0.0 -0.218 0 2.0 1e-06 
0.0 -0.2179 0 2.0 1e-06 
0.0 -0.2178 0 2.0 1e-06 
0.0 -0.2177 0 2.0 1e-06 
0.0 -0.2176 0 2.0 1e-06 
0.0 -0.2175 0 2.0 1e-06 
0.0 -0.2174 0 2.0 1e-06 
0.0 -0.2173 0 2.0 1e-06 
0.0 -0.2172 0 2.0 1e-06 
0.0 -0.2171 0 2.0 1e-06 
0.0 -0.217 0 2.0 1e-06 
0.0 -0.2169 0 2.0 1e-06 
0.0 -0.2168 0 2.0 1e-06 
0.0 -0.2167 0 2.0 1e-06 
0.0 -0.2166 0 2.0 1e-06 
0.0 -0.2165 0 2.0 1e-06 
0.0 -0.2164 0 2.0 1e-06 
0.0 -0.2163 0 2.0 1e-06 
0.0 -0.2162 0 2.0 1e-06 
0.0 -0.2161 0 2.0 1e-06 
0.0 -0.216 0 2.0 1e-06 
0.0 -0.2159 0 2.0 1e-06 
0.0 -0.2158 0 2.0 1e-06 
0.0 -0.2157 0 2.0 1e-06 
0.0 -0.2156 0 2.0 1e-06 
0.0 -0.2155 0 2.0 1e-06 
0.0 -0.2154 0 2.0 1e-06 
0.0 -0.2153 0 2.0 1e-06 
0.0 -0.2152 0 2.0 1e-06 
0.0 -0.2151 0 2.0 1e-06 
0.0 -0.215 0 2.0 1e-06 
0.0 -0.2149 0 2.0 1e-06 
0.0 -0.2148 0 2.0 1e-06 
0.0 -0.2147 0 2.0 1e-06 
0.0 -0.2146 0 2.0 1e-06 
0.0 -0.2145 0 2.0 1e-06 
0.0 -0.2144 0 2.0 1e-06 
0.0 -0.2143 0 2.0 1e-06 
0.0 -0.2142 0 2.0 1e-06 
0.0 -0.2141 0 2.0 1e-06 
0.0 -0.214 0 2.0 1e-06 
0.0 -0.2139 0 2.0 1e-06 
0.0 -0.2138 0 2.0 1e-06 
0.0 -0.2137 0 2.0 1e-06 
0.0 -0.2136 0 2.0 1e-06 
0.0 -0.2135 0 2.0 1e-06 
0.0 -0.2134 0 2.0 1e-06 
0.0 -0.2133 0 2.0 1e-06 
0.0 -0.2132 0 2.0 1e-06 
0.0 -0.2131 0 2.0 1e-06 
0.0 -0.213 0 2.0 1e-06 
0.0 -0.2129 0 2.0 1e-06 
0.0 -0.2128 0 2.0 1e-06 
0.0 -0.2127 0 2.0 1e-06 
0.0 -0.2126 0 2.0 1e-06 
0.0 -0.2125 0 2.0 1e-06 
0.0 -0.2124 0 2.0 1e-06 
0.0 -0.2123 0 2.0 1e-06 
0.0 -0.2122 0 2.0 1e-06 
0.0 -0.2121 0 2.0 1e-06 
0.0 -0.212 0 2.0 1e-06 
0.0 -0.2119 0 2.0 1e-06 
0.0 -0.2118 0 2.0 1e-06 
0.0 -0.2117 0 2.0 1e-06 
0.0 -0.2116 0 2.0 1e-06 
0.0 -0.2115 0 2.0 1e-06 
0.0 -0.2114 0 2.0 1e-06 
0.0 -0.2113 0 2.0 1e-06 
0.0 -0.2112 0 2.0 1e-06 
0.0 -0.2111 0 2.0 1e-06 
0.0 -0.211 0 2.0 1e-06 
0.0 -0.2109 0 2.0 1e-06 
0.0 -0.2108 0 2.0 1e-06 
0.0 -0.2107 0 2.0 1e-06 
0.0 -0.2106 0 2.0 1e-06 
0.0 -0.2105 0 2.0 1e-06 
0.0 -0.2104 0 2.0 1e-06 
0.0 -0.2103 0 2.0 1e-06 
0.0 -0.2102 0 2.0 1e-06 
0.0 -0.2101 0 2.0 1e-06 
0.0 -0.21 0 2.0 1e-06 
0.0 -0.2099 0 2.0 1e-06 
0.0 -0.2098 0 2.0 1e-06 
0.0 -0.2097 0 2.0 1e-06 
0.0 -0.2096 0 2.0 1e-06 
0.0 -0.2095 0 2.0 1e-06 
0.0 -0.2094 0 2.0 1e-06 
0.0 -0.2093 0 2.0 1e-06 
0.0 -0.2092 0 2.0 1e-06 
0.0 -0.2091 0 2.0 1e-06 
0.0 -0.209 0 2.0 1e-06 
0.0 -0.2089 0 2.0 1e-06 
0.0 -0.2088 0 2.0 1e-06 
0.0 -0.2087 0 2.0 1e-06 
0.0 -0.2086 0 2.0 1e-06 
0.0 -0.2085 0 2.0 1e-06 
0.0 -0.2084 0 2.0 1e-06 
0.0 -0.2083 0 2.0 1e-06 
0.0 -0.2082 0 2.0 1e-06 
0.0 -0.2081 0 2.0 1e-06 
0.0 -0.208 0 2.0 1e-06 
0.0 -0.2079 0 2.0 1e-06 
0.0 -0.2078 0 2.0 1e-06 
0.0 -0.2077 0 2.0 1e-06 
0.0 -0.2076 0 2.0 1e-06 
0.0 -0.2075 0 2.0 1e-06 
0.0 -0.2074 0 2.0 1e-06 
0.0 -0.2073 0 2.0 1e-06 
0.0 -0.2072 0 2.0 1e-06 
0.0 -0.2071 0 2.0 1e-06 
0.0 -0.207 0 2.0 1e-06 
0.0 -0.2069 0 2.0 1e-06 
0.0 -0.2068 0 2.0 1e-06 
0.0 -0.2067 0 2.0 1e-06 
0.0 -0.2066 0 2.0 1e-06 
0.0 -0.2065 0 2.0 1e-06 
0.0 -0.2064 0 2.0 1e-06 
0.0 -0.2063 0 2.0 1e-06 
0.0 -0.2062 0 2.0 1e-06 
0.0 -0.2061 0 2.0 1e-06 
0.0 -0.206 0 2.0 1e-06 
0.0 -0.2059 0 2.0 1e-06 
0.0 -0.2058 0 2.0 1e-06 
0.0 -0.2057 0 2.0 1e-06 
0.0 -0.2056 0 2.0 1e-06 
0.0 -0.2055 0 2.0 1e-06 
0.0 -0.2054 0 2.0 1e-06 
0.0 -0.2053 0 2.0 1e-06 
0.0 -0.2052 0 2.0 1e-06 
0.0 -0.2051 0 2.0 1e-06 
0.0 -0.205 0 2.0 1e-06 
0.0 -0.2049 0 2.0 1e-06 
0.0 -0.2048 0 2.0 1e-06 
0.0 -0.2047 0 2.0 1e-06 
0.0 -0.2046 0 2.0 1e-06 
0.0 -0.2045 0 2.0 1e-06 
0.0 -0.2044 0 2.0 1e-06 
0.0 -0.2043 0 2.0 1e-06 
0.0 -0.2042 0 2.0 1e-06 
0.0 -0.2041 0 2.0 1e-06 
0.0 -0.204 0 2.0 1e-06 
0.0 -0.2039 0 2.0 1e-06 
0.0 -0.2038 0 2.0 1e-06 
0.0 -0.2037 0 2.0 1e-06 
0.0 -0.2036 0 2.0 1e-06 
0.0 -0.2035 0 2.0 1e-06 
0.0 -0.2034 0 2.0 1e-06 
0.0 -0.2033 0 2.0 1e-06 
0.0 -0.2032 0 2.0 1e-06 
0.0 -0.2031 0 2.0 1e-06 
0.0 -0.203 0 2.0 1e-06 
0.0 -0.2029 0 2.0 1e-06 
0.0 -0.2028 0 2.0 1e-06 
0.0 -0.2027 0 2.0 1e-06 
0.0 -0.2026 0 2.0 1e-06 
0.0 -0.2025 0 2.0 1e-06 
0.0 -0.2024 0 2.0 1e-06 
0.0 -0.2023 0 2.0 1e-06 
0.0 -0.2022 0 2.0 1e-06 
0.0 -0.2021 0 2.0 1e-06 
0.0 -0.202 0 2.0 1e-06 
0.0 -0.2019 0 2.0 1e-06 
0.0 -0.2018 0 2.0 1e-06 
0.0 -0.2017 0 2.0 1e-06 
0.0 -0.2016 0 2.0 1e-06 
0.0 -0.2015 0 2.0 1e-06 
0.0 -0.2014 0 2.0 1e-06 
0.0 -0.2013 0 2.0 1e-06 
0.0 -0.2012 0 2.0 1e-06 
0.0 -0.2011 0 2.0 1e-06 
0.0 -0.201 0 2.0 1e-06 
0.0 -0.2009 0 2.0 1e-06 
0.0 -0.2008 0 2.0 1e-06 
0.0 -0.2007 0 2.0 1e-06 
0.0 -0.2006 0 2.0 1e-06 
0.0 -0.2005 0 2.0 1e-06 
0.0 -0.2004 0 2.0 1e-06 
0.0 -0.2003 0 2.0 1e-06 
0.0 -0.2002 0 2.0 1e-06 
0.0 -0.2001 0 2.0 1e-06 
0.0 -0.2 0 2.0 1e-06 
0.0 -0.1999 0 2.0 1e-06 
0.0 -0.1998 0 2.0 1e-06 
0.0 -0.1997 0 2.0 1e-06 
0.0 -0.1996 0 2.0 1e-06 
0.0 -0.1995 0 2.0 1e-06 
0.0 -0.1994 0 2.0 1e-06 
0.0 -0.1993 0 2.0 1e-06 
0.0 -0.1992 0 2.0 1e-06 
0.0 -0.1991 0 2.0 1e-06 
0.0 -0.199 0 2.0 1e-06 
0.0 -0.1989 0 2.0 1e-06 
0.0 -0.1988 0 2.0 1e-06 
0.0 -0.1987 0 2.0 1e-06 
0.0 -0.1986 0 2.0 1e-06 
0.0 -0.1985 0 2.0 1e-06 
0.0 -0.1984 0 2.0 1e-06 
0.0 -0.1983 0 2.0 1e-06 
0.0 -0.1982 0 2.0 1e-06 
0.0 -0.1981 0 2.0 1e-06 
0.0 -0.198 0 2.0 1e-06 
0.0 -0.1979 0 2.0 1e-06 
0.0 -0.1978 0 2.0 1e-06 
0.0 -0.1977 0 2.0 1e-06 
0.0 -0.1976 0 2.0 1e-06 
0.0 -0.1975 0 2.0 1e-06 
0.0 -0.1974 0 2.0 1e-06 
0.0 -0.1973 0 2.0 1e-06 
0.0 -0.1972 0 2.0 1e-06 
0.0 -0.1971 0 2.0 1e-06 
0.0 -0.197 0 2.0 1e-06 
0.0 -0.1969 0 2.0 1e-06 
0.0 -0.1968 0 2.0 1e-06 
0.0 -0.1967 0 2.0 1e-06 
0.0 -0.1966 0 2.0 1e-06 
0.0 -0.1965 0 2.0 1e-06 
0.0 -0.1964 0 2.0 1e-06 
0.0 -0.1963 0 2.0 1e-06 
0.0 -0.1962 0 2.0 1e-06 
0.0 -0.1961 0 2.0 1e-06 
0.0 -0.196 0 2.0 1e-06 
0.0 -0.1959 0 2.0 1e-06 
0.0 -0.1958 0 2.0 1e-06 
0.0 -0.1957 0 2.0 1e-06 
0.0 -0.1956 0 2.0 1e-06 
0.0 -0.1955 0 2.0 1e-06 
0.0 -0.1954 0 2.0 1e-06 
0.0 -0.1953 0 2.0 1e-06 
0.0 -0.1952 0 2.0 1e-06 
0.0 -0.1951 0 2.0 1e-06 
0.0 -0.195 0 2.0 1e-06 
0.0 -0.1949 0 2.0 1e-06 
0.0 -0.1948 0 2.0 1e-06 
0.0 -0.1947 0 2.0 1e-06 
0.0 -0.1946 0 2.0 1e-06 
0.0 -0.1945 0 2.0 1e-06 
0.0 -0.1944 0 2.0 1e-06 
0.0 -0.1943 0 2.0 1e-06 
0.0 -0.1942 0 2.0 1e-06 
0.0 -0.1941 0 2.0 1e-06 
0.0 -0.194 0 2.0 1e-06 
0.0 -0.1939 0 2.0 1e-06 
0.0 -0.1938 0 2.0 1e-06 
0.0 -0.1937 0 2.0 1e-06 
0.0 -0.1936 0 2.0 1e-06 
0.0 -0.1935 0 2.0 1e-06 
0.0 -0.1934 0 2.0 1e-06 
0.0 -0.1933 0 2.0 1e-06 
0.0 -0.1932 0 2.0 1e-06 
0.0 -0.1931 0 2.0 1e-06 
0.0 -0.193 0 2.0 1e-06 
0.0 -0.1929 0 2.0 1e-06 
0.0 -0.1928 0 2.0 1e-06 
0.0 -0.1927 0 2.0 1e-06 
0.0 -0.1926 0 2.0 1e-06 
0.0 -0.1925 0 2.0 1e-06 
0.0 -0.1924 0 2.0 1e-06 
0.0 -0.1923 0 2.0 1e-06 
0.0 -0.1922 0 2.0 1e-06 
0.0 -0.1921 0 2.0 1e-06 
0.0 -0.192 0 2.0 1e-06 
0.0 -0.1919 0 2.0 1e-06 
0.0 -0.1918 0 2.0 1e-06 
0.0 -0.1917 0 2.0 1e-06 
0.0 -0.1916 0 2.0 1e-06 
0.0 -0.1915 0 2.0 1e-06 
0.0 -0.1914 0 2.0 1e-06 
0.0 -0.1913 0 2.0 1e-06 
0.0 -0.1912 0 2.0 1e-06 
0.0 -0.1911 0 2.0 1e-06 
0.0 -0.191 0 2.0 1e-06 
0.0 -0.1909 0 2.0 1e-06 
0.0 -0.1908 0 2.0 1e-06 
0.0 -0.1907 0 2.0 1e-06 
0.0 -0.1906 0 2.0 1e-06 
0.0 -0.1905 0 2.0 1e-06 
0.0 -0.1904 0 2.0 1e-06 
0.0 -0.1903 0 2.0 1e-06 
0.0 -0.1902 0 2.0 1e-06 
0.0 -0.1901 0 2.0 1e-06 
0.0 -0.19 0 2.0 1e-06 
0.0 -0.1899 0 2.0 1e-06 
0.0 -0.1898 0 2.0 1e-06 
0.0 -0.1897 0 2.0 1e-06 
0.0 -0.1896 0 2.0 1e-06 
0.0 -0.1895 0 2.0 1e-06 
0.0 -0.1894 0 2.0 1e-06 
0.0 -0.1893 0 2.0 1e-06 
0.0 -0.1892 0 2.0 1e-06 
0.0 -0.1891 0 2.0 1e-06 
0.0 -0.189 0 2.0 1e-06 
0.0 -0.1889 0 2.0 1e-06 
0.0 -0.1888 0 2.0 1e-06 
0.0 -0.1887 0 2.0 1e-06 
0.0 -0.1886 0 2.0 1e-06 
0.0 -0.1885 0 2.0 1e-06 
0.0 -0.1884 0 2.0 1e-06 
0.0 -0.1883 0 2.0 1e-06 
0.0 -0.1882 0 2.0 1e-06 
0.0 -0.1881 0 2.0 1e-06 
0.0 -0.188 0 2.0 1e-06 
0.0 -0.1879 0 2.0 1e-06 
0.0 -0.1878 0 2.0 1e-06 
0.0 -0.1877 0 2.0 1e-06 
0.0 -0.1876 0 2.0 1e-06 
0.0 -0.1875 0 2.0 1e-06 
0.0 -0.1874 0 2.0 1e-06 
0.0 -0.1873 0 2.0 1e-06 
0.0 -0.1872 0 2.0 1e-06 
0.0 -0.1871 0 2.0 1e-06 
0.0 -0.187 0 2.0 1e-06 
0.0 -0.1869 0 2.0 1e-06 
0.0 -0.1868 0 2.0 1e-06 
0.0 -0.1867 0 2.0 1e-06 
0.0 -0.1866 0 2.0 1e-06 
0.0 -0.1865 0 2.0 1e-06 
0.0 -0.1864 0 2.0 1e-06 
0.0 -0.1863 0 2.0 1e-06 
0.0 -0.1862 0 2.0 1e-06 
0.0 -0.1861 0 2.0 1e-06 
0.0 -0.186 0 2.0 1e-06 
0.0 -0.1859 0 2.0 1e-06 
0.0 -0.1858 0 2.0 1e-06 
0.0 -0.1857 0 2.0 1e-06 
0.0 -0.1856 0 2.0 1e-06 
0.0 -0.1855 0 2.0 1e-06 
0.0 -0.1854 0 2.0 1e-06 
0.0 -0.1853 0 2.0 1e-06 
0.0 -0.1852 0 2.0 1e-06 
0.0 -0.1851 0 2.0 1e-06 
0.0 -0.185 0 2.0 1e-06 
0.0 -0.1849 0 2.0 1e-06 
0.0 -0.1848 0 2.0 1e-06 
0.0 -0.1847 0 2.0 1e-06 
0.0 -0.1846 0 2.0 1e-06 
0.0 -0.1845 0 2.0 1e-06 
0.0 -0.1844 0 2.0 1e-06 
0.0 -0.1843 0 2.0 1e-06 
0.0 -0.1842 0 2.0 1e-06 
0.0 -0.1841 0 2.0 1e-06 
0.0 -0.184 0 2.0 1e-06 
0.0 -0.1839 0 2.0 1e-06 
0.0 -0.1838 0 2.0 1e-06 
0.0 -0.1837 0 2.0 1e-06 
0.0 -0.1836 0 2.0 1e-06 
0.0 -0.1835 0 2.0 1e-06 
0.0 -0.1834 0 2.0 1e-06 
0.0 -0.1833 0 2.0 1e-06 
0.0 -0.1832 0 2.0 1e-06 
0.0 -0.1831 0 2.0 1e-06 
0.0 -0.183 0 2.0 1e-06 
0.0 -0.1829 0 2.0 1e-06 
0.0 -0.1828 0 2.0 1e-06 
0.0 -0.1827 0 2.0 1e-06 
0.0 -0.1826 0 2.0 1e-06 
0.0 -0.1825 0 2.0 1e-06 
0.0 -0.1824 0 2.0 1e-06 
0.0 -0.1823 0 2.0 1e-06 
0.0 -0.1822 0 2.0 1e-06 
0.0 -0.1821 0 2.0 1e-06 
0.0 -0.182 0 2.0 1e-06 
0.0 -0.1819 0 2.0 1e-06 
0.0 -0.1818 0 2.0 1e-06 
0.0 -0.1817 0 2.0 1e-06 
0.0 -0.1816 0 2.0 1e-06 
0.0 -0.1815 0 2.0 1e-06 
0.0 -0.1814 0 2.0 1e-06 
0.0 -0.1813 0 2.0 1e-06 
0.0 -0.1812 0 2.0 1e-06 
0.0 -0.1811 0 2.0 1e-06 
0.0 -0.181 0 2.0 1e-06 
0.0 -0.1809 0 2.0 1e-06 
0.0 -0.1808 0 2.0 1e-06 
0.0 -0.1807 0 2.0 1e-06 
0.0 -0.1806 0 2.0 1e-06 
0.0 -0.1805 0 2.0 1e-06 
0.0 -0.1804 0 2.0 1e-06 
0.0 -0.1803 0 2.0 1e-06 
0.0 -0.1802 0 2.0 1e-06 
0.0 -0.1801 0 2.0 1e-06 
0.0 -0.18 0 2.0 1e-06 
0.0 -0.1799 0 2.0 1e-06 
0.0 -0.1798 0 2.0 1e-06 
0.0 -0.1797 0 2.0 1e-06 
0.0 -0.1796 0 2.0 1e-06 
0.0 -0.1795 0 2.0 1e-06 
0.0 -0.1794 0 2.0 1e-06 
0.0 -0.1793 0 2.0 1e-06 
0.0 -0.1792 0 2.0 1e-06 
0.0 -0.1791 0 2.0 1e-06 
0.0 -0.179 0 2.0 1e-06 
0.0 -0.1789 0 2.0 1e-06 
0.0 -0.1788 0 2.0 1e-06 
0.0 -0.1787 0 2.0 1e-06 
0.0 -0.1786 0 2.0 1e-06 
0.0 -0.1785 0 2.0 1e-06 
0.0 -0.1784 0 2.0 1e-06 
0.0 -0.1783 0 2.0 1e-06 
0.0 -0.1782 0 2.0 1e-06 
0.0 -0.1781 0 2.0 1e-06 
0.0 -0.178 0 2.0 1e-06 
0.0 -0.1779 0 2.0 1e-06 
0.0 -0.1778 0 2.0 1e-06 
0.0 -0.1777 0 2.0 1e-06 
0.0 -0.1776 0 2.0 1e-06 
0.0 -0.1775 0 2.0 1e-06 
0.0 -0.1774 0 2.0 1e-06 
0.0 -0.1773 0 2.0 1e-06 
0.0 -0.1772 0 2.0 1e-06 
0.0 -0.1771 0 2.0 1e-06 
0.0 -0.177 0 2.0 1e-06 
0.0 -0.1769 0 2.0 1e-06 
0.0 -0.1768 0 2.0 1e-06 
0.0 -0.1767 0 2.0 1e-06 
0.0 -0.1766 0 2.0 1e-06 
0.0 -0.1765 0 2.0 1e-06 
0.0 -0.1764 0 2.0 1e-06 
0.0 -0.1763 0 2.0 1e-06 
0.0 -0.1762 0 2.0 1e-06 
0.0 -0.1761 0 2.0 1e-06 
0.0 -0.176 0 2.0 1e-06 
0.0 -0.1759 0 2.0 1e-06 
0.0 -0.1758 0 2.0 1e-06 
0.0 -0.1757 0 2.0 1e-06 
0.0 -0.1756 0 2.0 1e-06 
0.0 -0.1755 0 2.0 1e-06 
0.0 -0.1754 0 2.0 1e-06 
0.0 -0.1753 0 2.0 1e-06 
0.0 -0.1752 0 2.0 1e-06 
0.0 -0.1751 0 2.0 1e-06 
0.0 -0.175 0 2.0 1e-06 
0.0 -0.1749 0 2.0 1e-06 
0.0 -0.1748 0 2.0 1e-06 
0.0 -0.1747 0 2.0 1e-06 
0.0 -0.1746 0 2.0 1e-06 
0.0 -0.1745 0 2.0 1e-06 
0.0 -0.1744 0 2.0 1e-06 
0.0 -0.1743 0 2.0 1e-06 
0.0 -0.1742 0 2.0 1e-06 
0.0 -0.1741 0 2.0 1e-06 
0.0 -0.174 0 2.0 1e-06 
0.0 -0.1739 0 2.0 1e-06 
0.0 -0.1738 0 2.0 1e-06 
0.0 -0.1737 0 2.0 1e-06 
0.0 -0.1736 0 2.0 1e-06 
0.0 -0.1735 0 2.0 1e-06 
0.0 -0.1734 0 2.0 1e-06 
0.0 -0.1733 0 2.0 1e-06 
0.0 -0.1732 0 2.0 1e-06 
0.0 -0.1731 0 2.0 1e-06 
0.0 -0.173 0 2.0 1e-06 
0.0 -0.1729 0 2.0 1e-06 
0.0 -0.1728 0 2.0 1e-06 
0.0 -0.1727 0 2.0 1e-06 
0.0 -0.1726 0 2.0 1e-06 
0.0 -0.1725 0 2.0 1e-06 
0.0 -0.1724 0 2.0 1e-06 
0.0 -0.1723 0 2.0 1e-06 
0.0 -0.1722 0 2.0 1e-06 
0.0 -0.1721 0 2.0 1e-06 
0.0 -0.172 0 2.0 1e-06 
0.0 -0.1719 0 2.0 1e-06 
0.0 -0.1718 0 2.0 1e-06 
0.0 -0.1717 0 2.0 1e-06 
0.0 -0.1716 0 2.0 1e-06 
0.0 -0.1715 0 2.0 1e-06 
0.0 -0.1714 0 2.0 1e-06 
0.0 -0.1713 0 2.0 1e-06 
0.0 -0.1712 0 2.0 1e-06 
0.0 -0.1711 0 2.0 1e-06 
0.0 -0.171 0 2.0 1e-06 
0.0 -0.1709 0 2.0 1e-06 
0.0 -0.1708 0 2.0 1e-06 
0.0 -0.1707 0 2.0 1e-06 
0.0 -0.1706 0 2.0 1e-06 
0.0 -0.1705 0 2.0 1e-06 
0.0 -0.1704 0 2.0 1e-06 
0.0 -0.1703 0 2.0 1e-06 
0.0 -0.1702 0 2.0 1e-06 
0.0 -0.1701 0 2.0 1e-06 
0.0 -0.17 0 2.0 1e-06 
0.0 -0.1699 0 2.0 1e-06 
0.0 -0.1698 0 2.0 1e-06 
0.0 -0.1697 0 2.0 1e-06 
0.0 -0.1696 0 2.0 1e-06 
0.0 -0.1695 0 2.0 1e-06 
0.0 -0.1694 0 2.0 1e-06 
0.0 -0.1693 0 2.0 1e-06 
0.0 -0.1692 0 2.0 1e-06 
0.0 -0.1691 0 2.0 1e-06 
0.0 -0.169 0 2.0 1e-06 
0.0 -0.1689 0 2.0 1e-06 
0.0 -0.1688 0 2.0 1e-06 
0.0 -0.1687 0 2.0 1e-06 
0.0 -0.1686 0 2.0 1e-06 
0.0 -0.1685 0 2.0 1e-06 
0.0 -0.1684 0 2.0 1e-06 
0.0 -0.1683 0 2.0 1e-06 
0.0 -0.1682 0 2.0 1e-06 
0.0 -0.1681 0 2.0 1e-06 
0.0 -0.168 0 2.0 1e-06 
0.0 -0.1679 0 2.0 1e-06 
0.0 -0.1678 0 2.0 1e-06 
0.0 -0.1677 0 2.0 1e-06 
0.0 -0.1676 0 2.0 1e-06 
0.0 -0.1675 0 2.0 1e-06 
0.0 -0.1674 0 2.0 1e-06 
0.0 -0.1673 0 2.0 1e-06 
0.0 -0.1672 0 2.0 1e-06 
0.0 -0.1671 0 2.0 1e-06 
0.0 -0.167 0 2.0 1e-06 
0.0 -0.1669 0 2.0 1e-06 
0.0 -0.1668 0 2.0 1e-06 
0.0 -0.1667 0 2.0 1e-06 
0.0 -0.1666 0 2.0 1e-06 
0.0 -0.1665 0 2.0 1e-06 
0.0 -0.1664 0 2.0 1e-06 
0.0 -0.1663 0 2.0 1e-06 
0.0 -0.1662 0 2.0 1e-06 
0.0 -0.1661 0 2.0 1e-06 
0.0 -0.166 0 2.0 1e-06 
0.0 -0.1659 0 2.0 1e-06 
0.0 -0.1658 0 2.0 1e-06 
0.0 -0.1657 0 2.0 1e-06 
0.0 -0.1656 0 2.0 1e-06 
0.0 -0.1655 0 2.0 1e-06 
0.0 -0.1654 0 2.0 1e-06 
0.0 -0.1653 0 2.0 1e-06 
0.0 -0.1652 0 2.0 1e-06 
0.0 -0.1651 0 2.0 1e-06 
0.0 -0.165 0 2.0 1e-06 
0.0 -0.1649 0 2.0 1e-06 
0.0 -0.1648 0 2.0 1e-06 
0.0 -0.1647 0 2.0 1e-06 
0.0 -0.1646 0 2.0 1e-06 
0.0 -0.1645 0 2.0 1e-06 
0.0 -0.1644 0 2.0 1e-06 
0.0 -0.1643 0 2.0 1e-06 
0.0 -0.1642 0 2.0 1e-06 
0.0 -0.1641 0 2.0 1e-06 
0.0 -0.164 0 2.0 1e-06 
0.0 -0.1639 0 2.0 1e-06 
0.0 -0.1638 0 2.0 1e-06 
0.0 -0.1637 0 2.0 1e-06 
0.0 -0.1636 0 2.0 1e-06 
0.0 -0.1635 0 2.0 1e-06 
0.0 -0.1634 0 2.0 1e-06 
0.0 -0.1633 0 2.0 1e-06 
0.0 -0.1632 0 2.0 1e-06 
0.0 -0.1631 0 2.0 1e-06 
0.0 -0.163 0 2.0 1e-06 
0.0 -0.1629 0 2.0 1e-06 
0.0 -0.1628 0 2.0 1e-06 
0.0 -0.1627 0 2.0 1e-06 
0.0 -0.1626 0 2.0 1e-06 
0.0 -0.1625 0 2.0 1e-06 
0.0 -0.1624 0 2.0 1e-06 
0.0 -0.1623 0 2.0 1e-06 
0.0 -0.1622 0 2.0 1e-06 
0.0 -0.1621 0 2.0 1e-06 
0.0 -0.162 0 2.0 1e-06 
0.0 -0.1619 0 2.0 1e-06 
0.0 -0.1618 0 2.0 1e-06 
0.0 -0.1617 0 2.0 1e-06 
0.0 -0.1616 0 2.0 1e-06 
0.0 -0.1615 0 2.0 1e-06 
0.0 -0.1614 0 2.0 1e-06 
0.0 -0.1613 0 2.0 1e-06 
0.0 -0.1612 0 2.0 1e-06 
0.0 -0.1611 0 2.0 1e-06 
0.0 -0.161 0 2.0 1e-06 
0.0 -0.1609 0 2.0 1e-06 
0.0 -0.1608 0 2.0 1e-06 
0.0 -0.1607 0 2.0 1e-06 
0.0 -0.1606 0 2.0 1e-06 
0.0 -0.1605 0 2.0 1e-06 
0.0 -0.1604 0 2.0 1e-06 
0.0 -0.1603 0 2.0 1e-06 
0.0 -0.1602 0 2.0 1e-06 
0.0 -0.1601 0 2.0 1e-06 
0.0 -0.16 0 2.0 1e-06 
0.0 -0.1599 0 2.0 1e-06 
0.0 -0.1598 0 2.0 1e-06 
0.0 -0.1597 0 2.0 1e-06 
0.0 -0.1596 0 2.0 1e-06 
0.0 -0.1595 0 2.0 1e-06 
0.0 -0.1594 0 2.0 1e-06 
0.0 -0.1593 0 2.0 1e-06 
0.0 -0.1592 0 2.0 1e-06 
0.0 -0.1591 0 2.0 1e-06 
0.0 -0.159 0 2.0 1e-06 
0.0 -0.1589 0 2.0 1e-06 
0.0 -0.1588 0 2.0 1e-06 
0.0 -0.1587 0 2.0 1e-06 
0.0 -0.1586 0 2.0 1e-06 
0.0 -0.1585 0 2.0 1e-06 
0.0 -0.1584 0 2.0 1e-06 
0.0 -0.1583 0 2.0 1e-06 
0.0 -0.1582 0 2.0 1e-06 
0.0 -0.1581 0 2.0 1e-06 
0.0 -0.158 0 2.0 1e-06 
0.0 -0.1579 0 2.0 1e-06 
0.0 -0.1578 0 2.0 1e-06 
0.0 -0.1577 0 2.0 1e-06 
0.0 -0.1576 0 2.0 1e-06 
0.0 -0.1575 0 2.0 1e-06 
0.0 -0.1574 0 2.0 1e-06 
0.0 -0.1573 0 2.0 1e-06 
0.0 -0.1572 0 2.0 1e-06 
0.0 -0.1571 0 2.0 1e-06 
0.0 -0.157 0 2.0 1e-06 
0.0 -0.1569 0 2.0 1e-06 
0.0 -0.1568 0 2.0 1e-06 
0.0 -0.1567 0 2.0 1e-06 
0.0 -0.1566 0 2.0 1e-06 
0.0 -0.1565 0 2.0 1e-06 
0.0 -0.1564 0 2.0 1e-06 
0.0 -0.1563 0 2.0 1e-06 
0.0 -0.1562 0 2.0 1e-06 
0.0 -0.1561 0 2.0 1e-06 
0.0 -0.156 0 2.0 1e-06 
0.0 -0.1559 0 2.0 1e-06 
0.0 -0.1558 0 2.0 1e-06 
0.0 -0.1557 0 2.0 1e-06 
0.0 -0.1556 0 2.0 1e-06 
0.0 -0.1555 0 2.0 1e-06 
0.0 -0.1554 0 2.0 1e-06 
0.0 -0.1553 0 2.0 1e-06 
0.0 -0.1552 0 2.0 1e-06 
0.0 -0.1551 0 2.0 1e-06 
0.0 -0.155 0 2.0 1e-06 
0.0 -0.1549 0 2.0 1e-06 
0.0 -0.1548 0 2.0 1e-06 
0.0 -0.1547 0 2.0 1e-06 
0.0 -0.1546 0 2.0 1e-06 
0.0 -0.1545 0 2.0 1e-06 
0.0 -0.1544 0 2.0 1e-06 
0.0 -0.1543 0 2.0 1e-06 
0.0 -0.1542 0 2.0 1e-06 
0.0 -0.1541 0 2.0 1e-06 
0.0 -0.154 0 2.0 1e-06 
0.0 -0.1539 0 2.0 1e-06 
0.0 -0.1538 0 2.0 1e-06 
0.0 -0.1537 0 2.0 1e-06 
0.0 -0.1536 0 2.0 1e-06 
0.0 -0.1535 0 2.0 1e-06 
0.0 -0.1534 0 2.0 1e-06 
0.0 -0.1533 0 2.0 1e-06 
0.0 -0.1532 0 2.0 1e-06 
0.0 -0.1531 0 2.0 1e-06 
0.0 -0.153 0 2.0 1e-06 
0.0 -0.1529 0 2.0 1e-06 
0.0 -0.1528 0 2.0 1e-06 
0.0 -0.1527 0 2.0 1e-06 
0.0 -0.1526 0 2.0 1e-06 
0.0 -0.1525 0 2.0 1e-06 
0.0 -0.1524 0 2.0 1e-06 
0.0 -0.1523 0 2.0 1e-06 
0.0 -0.1522 0 2.0 1e-06 
0.0 -0.1521 0 2.0 1e-06 
0.0 -0.152 0 2.0 1e-06 
0.0 -0.1519 0 2.0 1e-06 
0.0 -0.1518 0 2.0 1e-06 
0.0 -0.1517 0 2.0 1e-06 
0.0 -0.1516 0 2.0 1e-06 
0.0 -0.1515 0 2.0 1e-06 
0.0 -0.1514 0 2.0 1e-06 
0.0 -0.1513 0 2.0 1e-06 
0.0 -0.1512 0 2.0 1e-06 
0.0 -0.1511 0 2.0 1e-06 
0.0 -0.151 0 2.0 1e-06 
0.0 -0.1509 0 2.0 1e-06 
0.0 -0.1508 0 2.0 1e-06 
0.0 -0.1507 0 2.0 1e-06 
0.0 -0.1506 0 2.0 1e-06 
0.0 -0.1505 0 2.0 1e-06 
0.0 -0.1504 0 2.0 1e-06 
0.0 -0.1503 0 2.0 1e-06 
0.0 -0.1502 0 2.0 1e-06 
0.0 -0.1501 0 2.0 1e-06 
0.0 -0.15 0 2.0 1e-06 
0.0 -0.1499 0 2.0 1e-06 
0.0 -0.1498 0 2.0 1e-06 
0.0 -0.1497 0 2.0 1e-06 
0.0 -0.1496 0 2.0 1e-06 
0.0 -0.1495 0 2.0 1e-06 
0.0 -0.1494 0 2.0 1e-06 
0.0 -0.1493 0 2.0 1e-06 
0.0 -0.1492 0 2.0 1e-06 
0.0 -0.1491 0 2.0 1e-06 
0.0 -0.149 0 2.0 1e-06 
0.0 -0.1489 0 2.0 1e-06 
0.0 -0.1488 0 2.0 1e-06 
0.0 -0.1487 0 2.0 1e-06 
0.0 -0.1486 0 2.0 1e-06 
0.0 -0.1485 0 2.0 1e-06 
0.0 -0.1484 0 2.0 1e-06 
0.0 -0.1483 0 2.0 1e-06 
0.0 -0.1482 0 2.0 1e-06 
0.0 -0.1481 0 2.0 1e-06 
0.0 -0.148 0 2.0 1e-06 
0.0 -0.1479 0 2.0 1e-06 
0.0 -0.1478 0 2.0 1e-06 
0.0 -0.1477 0 2.0 1e-06 
0.0 -0.1476 0 2.0 1e-06 
0.0 -0.1475 0 2.0 1e-06 
0.0 -0.1474 0 2.0 1e-06 
0.0 -0.1473 0 2.0 1e-06 
0.0 -0.1472 0 2.0 1e-06 
0.0 -0.1471 0 2.0 1e-06 
0.0 -0.147 0 2.0 1e-06 
0.0 -0.1469 0 2.0 1e-06 
0.0 -0.1468 0 2.0 1e-06 
0.0 -0.1467 0 2.0 1e-06 
0.0 -0.1466 0 2.0 1e-06 
0.0 -0.1465 0 2.0 1e-06 
0.0 -0.1464 0 2.0 1e-06 
0.0 -0.1463 0 2.0 1e-06 
0.0 -0.1462 0 2.0 1e-06 
0.0 -0.1461 0 2.0 1e-06 
0.0 -0.146 0 2.0 1e-06 
0.0 -0.1459 0 2.0 1e-06 
0.0 -0.1458 0 2.0 1e-06 
0.0 -0.1457 0 2.0 1e-06 
0.0 -0.1456 0 2.0 1e-06 
0.0 -0.1455 0 2.0 1e-06 
0.0 -0.1454 0 2.0 1e-06 
0.0 -0.1453 0 2.0 1e-06 
0.0 -0.1452 0 2.0 1e-06 
0.0 -0.1451 0 2.0 1e-06 
0.0 -0.145 0 2.0 1e-06 
0.0 -0.1449 0 2.0 1e-06 
0.0 -0.1448 0 2.0 1e-06 
0.0 -0.1447 0 2.0 1e-06 
0.0 -0.1446 0 2.0 1e-06 
0.0 -0.1445 0 2.0 1e-06 
0.0 -0.1444 0 2.0 1e-06 
0.0 -0.1443 0 2.0 1e-06 
0.0 -0.1442 0 2.0 1e-06 
0.0 -0.1441 0 2.0 1e-06 
0.0 -0.144 0 2.0 1e-06 
0.0 -0.1439 0 2.0 1e-06 
0.0 -0.1438 0 2.0 1e-06 
0.0 -0.1437 0 2.0 1e-06 
0.0 -0.1436 0 2.0 1e-06 
0.0 -0.1435 0 2.0 1e-06 
0.0 -0.1434 0 2.0 1e-06 
0.0 -0.1433 0 2.0 1e-06 
0.0 -0.1432 0 2.0 1e-06 
0.0 -0.1431 0 2.0 1e-06 
0.0 -0.143 0 2.0 1e-06 
0.0 -0.1429 0 2.0 1e-06 
0.0 -0.1428 0 2.0 1e-06 
0.0 -0.1427 0 2.0 1e-06 
0.0 -0.1426 0 2.0 1e-06 
0.0 -0.1425 0 2.0 1e-06 
0.0 -0.1424 0 2.0 1e-06 
0.0 -0.1423 0 2.0 1e-06 
0.0 -0.1422 0 2.0 1e-06 
0.0 -0.1421 0 2.0 1e-06 
0.0 -0.142 0 2.0 1e-06 
0.0 -0.1419 0 2.0 1e-06 
0.0 -0.1418 0 2.0 1e-06 
0.0 -0.1417 0 2.0 1e-06 
0.0 -0.1416 0 2.0 1e-06 
0.0 -0.1415 0 2.0 1e-06 
0.0 -0.1414 0 2.0 1e-06 
0.0 -0.1413 0 2.0 1e-06 
0.0 -0.1412 0 2.0 1e-06 
0.0 -0.1411 0 2.0 1e-06 
0.0 -0.141 0 2.0 1e-06 
0.0 -0.1409 0 2.0 1e-06 
0.0 -0.1408 0 2.0 1e-06 
0.0 -0.1407 0 2.0 1e-06 
0.0 -0.1406 0 2.0 1e-06 
0.0 -0.1405 0 2.0 1e-06 
0.0 -0.1404 0 2.0 1e-06 
0.0 -0.1403 0 2.0 1e-06 
0.0 -0.1402 0 2.0 1e-06 
0.0 -0.1401 0 2.0 1e-06 
0.0 -0.14 0 2.0 1e-06 
0.0 -0.1399 0 2.0 1e-06 
0.0 -0.1398 0 2.0 1e-06 
0.0 -0.1397 0 2.0 1e-06 
0.0 -0.1396 0 2.0 1e-06 
0.0 -0.1395 0 2.0 1e-06 
0.0 -0.1394 0 2.0 1e-06 
0.0 -0.1393 0 2.0 1e-06 
0.0 -0.1392 0 2.0 1e-06 
0.0 -0.1391 0 2.0 1e-06 
0.0 -0.139 0 2.0 1e-06 
0.0 -0.1389 0 2.0 1e-06 
0.0 -0.1388 0 2.0 1e-06 
0.0 -0.1387 0 2.0 1e-06 
0.0 -0.1386 0 2.0 1e-06 
0.0 -0.1385 0 2.0 1e-06 
0.0 -0.1384 0 2.0 1e-06 
0.0 -0.1383 0 2.0 1e-06 
0.0 -0.1382 0 2.0 1e-06 
0.0 -0.1381 0 2.0 1e-06 
0.0 -0.138 0 2.0 1e-06 
0.0 -0.1379 0 2.0 1e-06 
0.0 -0.1378 0 2.0 1e-06 
0.0 -0.1377 0 2.0 1e-06 
0.0 -0.1376 0 2.0 1e-06 
0.0 -0.1375 0 2.0 1e-06 
0.0 -0.1374 0 2.0 1e-06 
0.0 -0.1373 0 2.0 1e-06 
0.0 -0.1372 0 2.0 1e-06 
0.0 -0.1371 0 2.0 1e-06 
0.0 -0.137 0 2.0 1e-06 
0.0 -0.1369 0 2.0 1e-06 
0.0 -0.1368 0 2.0 1e-06 
0.0 -0.1367 0 2.0 1e-06 
0.0 -0.1366 0 2.0 1e-06 
0.0 -0.1365 0 2.0 1e-06 
0.0 -0.1364 0 2.0 1e-06 
0.0 -0.1363 0 2.0 1e-06 
0.0 -0.1362 0 2.0 1e-06 
0.0 -0.1361 0 2.0 1e-06 
0.0 -0.136 0 2.0 1e-06 
0.0 -0.1359 0 2.0 1e-06 
0.0 -0.1358 0 2.0 1e-06 
0.0 -0.1357 0 2.0 1e-06 
0.0 -0.1356 0 2.0 1e-06 
0.0 -0.1355 0 2.0 1e-06 
0.0 -0.1354 0 2.0 1e-06 
0.0 -0.1353 0 2.0 1e-06 
0.0 -0.1352 0 2.0 1e-06 
0.0 -0.1351 0 2.0 1e-06 
0.0 -0.135 0 2.0 1e-06 
0.0 -0.1349 0 2.0 1e-06 
0.0 -0.1348 0 2.0 1e-06 
0.0 -0.1347 0 2.0 1e-06 
0.0 -0.1346 0 2.0 1e-06 
0.0 -0.1345 0 2.0 1e-06 
0.0 -0.1344 0 2.0 1e-06 
0.0 -0.1343 0 2.0 1e-06 
0.0 -0.1342 0 2.0 1e-06 
0.0 -0.1341 0 2.0 1e-06 
0.0 -0.134 0 2.0 1e-06 
0.0 -0.1339 0 2.0 1e-06 
0.0 -0.1338 0 2.0 1e-06 
0.0 -0.1337 0 2.0 1e-06 
0.0 -0.1336 0 2.0 1e-06 
0.0 -0.1335 0 2.0 1e-06 
0.0 -0.1334 0 2.0 1e-06 
0.0 -0.1333 0 2.0 1e-06 
0.0 -0.1332 0 2.0 1e-06 
0.0 -0.1331 0 2.0 1e-06 
0.0 -0.133 0 2.0 1e-06 
0.0 -0.1329 0 2.0 1e-06 
0.0 -0.1328 0 2.0 1e-06 
0.0 -0.1327 0 2.0 1e-06 
0.0 -0.1326 0 2.0 1e-06 
0.0 -0.1325 0 2.0 1e-06 
0.0 -0.1324 0 2.0 1e-06 
0.0 -0.1323 0 2.0 1e-06 
0.0 -0.1322 0 2.0 1e-06 
0.0 -0.1321 0 2.0 1e-06 
0.0 -0.132 0 2.0 1e-06 
0.0 -0.1319 0 2.0 1e-06 
0.0 -0.1318 0 2.0 1e-06 
0.0 -0.1317 0 2.0 1e-06 
0.0 -0.1316 0 2.0 1e-06 
0.0 -0.1315 0 2.0 1e-06 
0.0 -0.1314 0 2.0 1e-06 
0.0 -0.1313 0 2.0 1e-06 
0.0 -0.1312 0 2.0 1e-06 
0.0 -0.1311 0 2.0 1e-06 
0.0 -0.131 0 2.0 1e-06 
0.0 -0.1309 0 2.0 1e-06 
0.0 -0.1308 0 2.0 1e-06 
0.0 -0.1307 0 2.0 1e-06 
0.0 -0.1306 0 2.0 1e-06 
0.0 -0.1305 0 2.0 1e-06 
0.0 -0.1304 0 2.0 1e-06 
0.0 -0.1303 0 2.0 1e-06 
0.0 -0.1302 0 2.0 1e-06 
0.0 -0.1301 0 2.0 1e-06 
0.0 -0.13 0 2.0 1e-06 
0.0 -0.1299 0 2.0 1e-06 
0.0 -0.1298 0 2.0 1e-06 
0.0 -0.1297 0 2.0 1e-06 
0.0 -0.1296 0 2.0 1e-06 
0.0 -0.1295 0 2.0 1e-06 
0.0 -0.1294 0 2.0 1e-06 
0.0 -0.1293 0 2.0 1e-06 
0.0 -0.1292 0 2.0 1e-06 
0.0 -0.1291 0 2.0 1e-06 
0.0 -0.129 0 2.0 1e-06 
0.0 -0.1289 0 2.0 1e-06 
0.0 -0.1288 0 2.0 1e-06 
0.0 -0.1287 0 2.0 1e-06 
0.0 -0.1286 0 2.0 1e-06 
0.0 -0.1285 0 2.0 1e-06 
0.0 -0.1284 0 2.0 1e-06 
0.0 -0.1283 0 2.0 1e-06 
0.0 -0.1282 0 2.0 1e-06 
0.0 -0.1281 0 2.0 1e-06 
0.0 -0.128 0 2.0 1e-06 
0.0 -0.1279 0 2.0 1e-06 
0.0 -0.1278 0 2.0 1e-06 
0.0 -0.1277 0 2.0 1e-06 
0.0 -0.1276 0 2.0 1e-06 
0.0 -0.1275 0 2.0 1e-06 
0.0 -0.1274 0 2.0 1e-06 
0.0 -0.1273 0 2.0 1e-06 
0.0 -0.1272 0 2.0 1e-06 
0.0 -0.1271 0 2.0 1e-06 
0.0 -0.127 0 2.0 1e-06 
0.0 -0.1269 0 2.0 1e-06 
0.0 -0.1268 0 2.0 1e-06 
0.0 -0.1267 0 2.0 1e-06 
0.0 -0.1266 0 2.0 1e-06 
0.0 -0.1265 0 2.0 1e-06 
0.0 -0.1264 0 2.0 1e-06 
0.0 -0.1263 0 2.0 1e-06 
0.0 -0.1262 0 2.0 1e-06 
0.0 -0.1261 0 2.0 1e-06 
0.0 -0.126 0 2.0 1e-06 
0.0 -0.1259 0 2.0 1e-06 
0.0 -0.1258 0 2.0 1e-06 
0.0 -0.1257 0 2.0 1e-06 
0.0 -0.1256 0 2.0 1e-06 
0.0 -0.1255 0 2.0 1e-06 
0.0 -0.1254 0 2.0 1e-06 
0.0 -0.1253 0 2.0 1e-06 
0.0 -0.1252 0 2.0 1e-06 
0.0 -0.1251 0 2.0 1e-06 
0.0 -0.125 0 2.0 1e-06 
0.0 -0.1249 0 2.0 1e-06 
0.0 -0.1248 0 2.0 1e-06 
0.0 -0.1247 0 2.0 1e-06 
0.0 -0.1246 0 2.0 1e-06 
0.0 -0.1245 0 2.0 1e-06 
0.0 -0.1244 0 2.0 1e-06 
0.0 -0.1243 0 2.0 1e-06 
0.0 -0.1242 0 2.0 1e-06 
0.0 -0.1241 0 2.0 1e-06 
0.0 -0.124 0 2.0 1e-06 
0.0 -0.1239 0 2.0 1e-06 
0.0 -0.1238 0 2.0 1e-06 
0.0 -0.1237 0 2.0 1e-06 
0.0 -0.1236 0 2.0 1e-06 
0.0 -0.1235 0 2.0 1e-06 
0.0 -0.1234 0 2.0 1e-06 
0.0 -0.1233 0 2.0 1e-06 
0.0 -0.1232 0 2.0 1e-06 
0.0 -0.1231 0 2.0 1e-06 
0.0 -0.123 0 2.0 1e-06 
0.0 -0.1229 0 2.0 1e-06 
0.0 -0.1228 0 2.0 1e-06 
0.0 -0.1227 0 2.0 1e-06 
0.0 -0.1226 0 2.0 1e-06 
0.0 -0.1225 0 2.0 1e-06 
0.0 -0.1224 0 2.0 1e-06 
0.0 -0.1223 0 2.0 1e-06 
0.0 -0.1222 0 2.0 1e-06 
0.0 -0.1221 0 2.0 1e-06 
0.0 -0.122 0 2.0 1e-06 
0.0 -0.1219 0 2.0 1e-06 
0.0 -0.1218 0 2.0 1e-06 
0.0 -0.1217 0 2.0 1e-06 
0.0 -0.1216 0 2.0 1e-06 
0.0 -0.1215 0 2.0 1e-06 
0.0 -0.1214 0 2.0 1e-06 
0.0 -0.1213 0 2.0 1e-06 
0.0 -0.1212 0 2.0 1e-06 
0.0 -0.1211 0 2.0 1e-06 
0.0 -0.121 0 2.0 1e-06 
0.0 -0.1209 0 2.0 1e-06 
0.0 -0.1208 0 2.0 1e-06 
0.0 -0.1207 0 2.0 1e-06 
0.0 -0.1206 0 2.0 1e-06 
0.0 -0.1205 0 2.0 1e-06 
0.0 -0.1204 0 2.0 1e-06 
0.0 -0.1203 0 2.0 1e-06 
0.0 -0.1202 0 2.0 1e-06 
0.0 -0.1201 0 2.0 1e-06 
0.0 -0.12 0 2.0 1e-06 
0.0 -0.1199 0 2.0 1e-06 
0.0 -0.1198 0 2.0 1e-06 
0.0 -0.1197 0 2.0 1e-06 
0.0 -0.1196 0 2.0 1e-06 
0.0 -0.1195 0 2.0 1e-06 
0.0 -0.1194 0 2.0 1e-06 
0.0 -0.1193 0 2.0 1e-06 
0.0 -0.1192 0 2.0 1e-06 
0.0 -0.1191 0 2.0 1e-06 
0.0 -0.119 0 2.0 1e-06 
0.0 -0.1189 0 2.0 1e-06 
0.0 -0.1188 0 2.0 1e-06 
0.0 -0.1187 0 2.0 1e-06 
0.0 -0.1186 0 2.0 1e-06 
0.0 -0.1185 0 2.0 1e-06 
0.0 -0.1184 0 2.0 1e-06 
0.0 -0.1183 0 2.0 1e-06 
0.0 -0.1182 0 2.0 1e-06 
0.0 -0.1181 0 2.0 1e-06 
0.0 -0.118 0 2.0 1e-06 
0.0 -0.1179 0 2.0 1e-06 
0.0 -0.1178 0 2.0 1e-06 
0.0 -0.1177 0 2.0 1e-06 
0.0 -0.1176 0 2.0 1e-06 
0.0 -0.1175 0 2.0 1e-06 
0.0 -0.1174 0 2.0 1e-06 
0.0 -0.1173 0 2.0 1e-06 
0.0 -0.1172 0 2.0 1e-06 
0.0 -0.1171 0 2.0 1e-06 
0.0 -0.117 0 2.0 1e-06 
0.0 -0.1169 0 2.0 1e-06 
0.0 -0.1168 0 2.0 1e-06 
0.0 -0.1167 0 2.0 1e-06 
0.0 -0.1166 0 2.0 1e-06 
0.0 -0.1165 0 2.0 1e-06 
0.0 -0.1164 0 2.0 1e-06 
0.0 -0.1163 0 2.0 1e-06 
0.0 -0.1162 0 2.0 1e-06 
0.0 -0.1161 0 2.0 1e-06 
0.0 -0.116 0 2.0 1e-06 
0.0 -0.1159 0 2.0 1e-06 
0.0 -0.1158 0 2.0 1e-06 
0.0 -0.1157 0 2.0 1e-06 
0.0 -0.1156 0 2.0 1e-06 
0.0 -0.1155 0 2.0 1e-06 
0.0 -0.1154 0 2.0 1e-06 
0.0 -0.1153 0 2.0 1e-06 
0.0 -0.1152 0 2.0 1e-06 
0.0 -0.1151 0 2.0 1e-06 
0.0 -0.115 0 2.0 1e-06 
0.0 -0.1149 0 2.0 1e-06 
0.0 -0.1148 0 2.0 1e-06 
0.0 -0.1147 0 2.0 1e-06 
0.0 -0.1146 0 2.0 1e-06 
0.0 -0.1145 0 2.0 1e-06 
0.0 -0.1144 0 2.0 1e-06 
0.0 -0.1143 0 2.0 1e-06 
0.0 -0.1142 0 2.0 1e-06 
0.0 -0.1141 0 2.0 1e-06 
0.0 -0.114 0 2.0 1e-06 
0.0 -0.1139 0 2.0 1e-06 
0.0 -0.1138 0 2.0 1e-06 
0.0 -0.1137 0 2.0 1e-06 
0.0 -0.1136 0 2.0 1e-06 
0.0 -0.1135 0 2.0 1e-06 
0.0 -0.1134 0 2.0 1e-06 
0.0 -0.1133 0 2.0 1e-06 
0.0 -0.1132 0 2.0 1e-06 
0.0 -0.1131 0 2.0 1e-06 
0.0 -0.113 0 2.0 1e-06 
0.0 -0.1129 0 2.0 1e-06 
0.0 -0.1128 0 2.0 1e-06 
0.0 -0.1127 0 2.0 1e-06 
0.0 -0.1126 0 2.0 1e-06 
0.0 -0.1125 0 2.0 1e-06 
0.0 -0.1124 0 2.0 1e-06 
0.0 -0.1123 0 2.0 1e-06 
0.0 -0.1122 0 2.0 1e-06 
0.0 -0.1121 0 2.0 1e-06 
0.0 -0.112 0 2.0 1e-06 
0.0 -0.1119 0 2.0 1e-06 
0.0 -0.1118 0 2.0 1e-06 
0.0 -0.1117 0 2.0 1e-06 
0.0 -0.1116 0 2.0 1e-06 
0.0 -0.1115 0 2.0 1e-06 
0.0 -0.1114 0 2.0 1e-06 
0.0 -0.1113 0 2.0 1e-06 
0.0 -0.1112 0 2.0 1e-06 
0.0 -0.1111 0 2.0 1e-06 
0.0 -0.111 0 2.0 1e-06 
0.0 -0.1109 0 2.0 1e-06 
0.0 -0.1108 0 2.0 1e-06 
0.0 -0.1107 0 2.0 1e-06 
0.0 -0.1106 0 2.0 1e-06 
0.0 -0.1105 0 2.0 1e-06 
0.0 -0.1104 0 2.0 1e-06 
0.0 -0.1103 0 2.0 1e-06 
0.0 -0.1102 0 2.0 1e-06 
0.0 -0.1101 0 2.0 1e-06 
0.0 -0.11 0 2.0 1e-06 
0.0 -0.1099 0 2.0 1e-06 
0.0 -0.1098 0 2.0 1e-06 
0.0 -0.1097 0 2.0 1e-06 
0.0 -0.1096 0 2.0 1e-06 
0.0 -0.1095 0 2.0 1e-06 
0.0 -0.1094 0 2.0 1e-06 
0.0 -0.1093 0 2.0 1e-06 
0.0 -0.1092 0 2.0 1e-06 
0.0 -0.1091 0 2.0 1e-06 
0.0 -0.109 0 2.0 1e-06 
0.0 -0.1089 0 2.0 1e-06 
0.0 -0.1088 0 2.0 1e-06 
0.0 -0.1087 0 2.0 1e-06 
0.0 -0.1086 0 2.0 1e-06 
0.0 -0.1085 0 2.0 1e-06 
0.0 -0.1084 0 2.0 1e-06 
0.0 -0.1083 0 2.0 1e-06 
0.0 -0.1082 0 2.0 1e-06 
0.0 -0.1081 0 2.0 1e-06 
0.0 -0.108 0 2.0 1e-06 
0.0 -0.1079 0 2.0 1e-06 
0.0 -0.1078 0 2.0 1e-06 
0.0 -0.1077 0 2.0 1e-06 
0.0 -0.1076 0 2.0 1e-06 
0.0 -0.1075 0 2.0 1e-06 
0.0 -0.1074 0 2.0 1e-06 
0.0 -0.1073 0 2.0 1e-06 
0.0 -0.1072 0 2.0 1e-06 
0.0 -0.1071 0 2.0 1e-06 
0.0 -0.107 0 2.0 1e-06 
0.0 -0.1069 0 2.0 1e-06 
0.0 -0.1068 0 2.0 1e-06 
0.0 -0.1067 0 2.0 1e-06 
0.0 -0.1066 0 2.0 1e-06 
0.0 -0.1065 0 2.0 1e-06 
0.0 -0.1064 0 2.0 1e-06 
0.0 -0.1063 0 2.0 1e-06 
0.0 -0.1062 0 2.0 1e-06 
0.0 -0.1061 0 2.0 1e-06 
0.0 -0.106 0 2.0 1e-06 
0.0 -0.1059 0 2.0 1e-06 
0.0 -0.1058 0 2.0 1e-06 
0.0 -0.1057 0 2.0 1e-06 
0.0 -0.1056 0 2.0 1e-06 
0.0 -0.1055 0 2.0 1e-06 
0.0 -0.1054 0 2.0 1e-06 
0.0 -0.1053 0 2.0 1e-06 
0.0 -0.1052 0 2.0 1e-06 
0.0 -0.1051 0 2.0 1e-06 
0.0 -0.105 0 2.0 1e-06 
0.0 -0.1049 0 2.0 1e-06 
0.0 -0.1048 0 2.0 1e-06 
0.0 -0.1047 0 2.0 1e-06 
0.0 -0.1046 0 2.0 1e-06 
0.0 -0.1045 0 2.0 1e-06 
0.0 -0.1044 0 2.0 1e-06 
0.0 -0.1043 0 2.0 1e-06 
0.0 -0.1042 0 2.0 1e-06 
0.0 -0.1041 0 2.0 1e-06 
0.0 -0.104 0 2.0 1e-06 
0.0 -0.1039 0 2.0 1e-06 
0.0 -0.1038 0 2.0 1e-06 
0.0 -0.1037 0 2.0 1e-06 
0.0 -0.1036 0 2.0 1e-06 
0.0 -0.1035 0 2.0 1e-06 
0.0 -0.1034 0 2.0 1e-06 
0.0 -0.1033 0 2.0 1e-06 
0.0 -0.1032 0 2.0 1e-06 
0.0 -0.1031 0 2.0 1e-06 
0.0 -0.103 0 2.0 1e-06 
0.0 -0.1029 0 2.0 1e-06 
0.0 -0.1028 0 2.0 1e-06 
0.0 -0.1027 0 2.0 1e-06 
0.0 -0.1026 0 2.0 1e-06 
0.0 -0.1025 0 2.0 1e-06 
0.0 -0.1024 0 2.0 1e-06 
0.0 -0.1023 0 2.0 1e-06 
0.0 -0.1022 0 2.0 1e-06 
0.0 -0.1021 0 2.0 1e-06 
0.0 -0.102 0 2.0 1e-06 
0.0 -0.1019 0 2.0 1e-06 
0.0 -0.1018 0 2.0 1e-06 
0.0 -0.1017 0 2.0 1e-06 
0.0 -0.1016 0 2.0 1e-06 
0.0 -0.1015 0 2.0 1e-06 
0.0 -0.1014 0 2.0 1e-06 
0.0 -0.1013 0 2.0 1e-06 
0.0 -0.1012 0 2.0 1e-06 
0.0 -0.1011 0 2.0 1e-06 
0.0 -0.101 0 2.0 1e-06 
0.0 -0.1009 0 2.0 1e-06 
0.0 -0.1008 0 2.0 1e-06 
0.0 -0.1007 0 2.0 1e-06 
0.0 -0.1006 0 2.0 1e-06 
0.0 -0.1005 0 2.0 1e-06 
0.0 -0.1004 0 2.0 1e-06 
0.0 -0.1003 0 2.0 1e-06 
0.0 -0.1002 0 2.0 1e-06 
0.0 -0.1001 0 2.0 1e-06 
0.0 -0.1 0 2.0 1e-06 
0.0 -0.0999000000002 0 2.0 1e-06 
0.0 -0.0998000000002 0 2.0 1e-06 
0.0 -0.0997000000002 0 2.0 1e-06 
0.0 -0.0996000000002 0 2.0 1e-06 
0.0 -0.0995000000002 0 2.0 1e-06 
0.0 -0.0994000000002 0 2.0 1e-06 
0.0 -0.0993000000002 0 2.0 1e-06 
0.0 -0.0992000000002 0 2.0 1e-06 
0.0 -0.0991000000002 0 2.0 1e-06 
0.0 -0.0990000000002 0 2.0 1e-06 
0.0 -0.0989000000002 0 2.0 1e-06 
0.0 -0.0988000000002 0 2.0 1e-06 
0.0 -0.0987000000002 0 2.0 1e-06 
0.0 -0.0986000000002 0 2.0 1e-06 
0.0 -0.0985000000002 0 2.0 1e-06 
0.0 -0.0984000000002 0 2.0 1e-06 
0.0 -0.0983000000002 0 2.0 1e-06 
0.0 -0.0982000000002 0 2.0 1e-06 
0.0 -0.0981000000002 0 2.0 1e-06 
0.0 -0.0980000000002 0 2.0 1e-06 
0.0 -0.0979000000002 0 2.0 1e-06 
0.0 -0.0978000000002 0 2.0 1e-06 
0.0 -0.0977000000002 0 2.0 1e-06 
0.0 -0.0976000000002 0 2.0 1e-06 
0.0 -0.0975000000002 0 2.0 1e-06 
0.0 -0.0974000000002 0 2.0 1e-06 
0.0 -0.0973000000002 0 2.0 1e-06 
0.0 -0.0972000000002 0 2.0 1e-06 
0.0 -0.0971000000002 0 2.0 1e-06 
0.0 -0.0970000000002 0 2.0 1e-06 
0.0 -0.0969000000002 0 2.0 1e-06 
0.0 -0.0968000000002 0 2.0 1e-06 
0.0 -0.0967000000002 0 2.0 1e-06 
0.0 -0.0966000000002 0 2.0 1e-06 
0.0 -0.0965000000002 0 2.0 1e-06 
0.0 -0.0964000000002 0 2.0 1e-06 
0.0 -0.0963000000002 0 2.0 1e-06 
0.0 -0.0962000000002 0 2.0 1e-06 
0.0 -0.0961000000002 0 2.0 1e-06 
0.0 -0.0960000000002 0 2.0 1e-06 
0.0 -0.0959000000002 0 2.0 1e-06 
0.0 -0.0958000000002 0 2.0 1e-06 
0.0 -0.0957000000002 0 2.0 1e-06 
0.0 -0.0956000000002 0 2.0 1e-06 
0.0 -0.0955000000002 0 2.0 1e-06 
0.0 -0.0954000000002 0 2.0 1e-06 
0.0 -0.0953000000002 0 2.0 1e-06 
0.0 -0.0952000000002 0 2.0 1e-06 
0.0 -0.0951000000002 0 2.0 1e-06 
0.0 -0.0950000000002 0 2.0 1e-06 
0.0 -0.0949000000002 0 2.0 1e-06 
0.0 -0.0948000000002 0 2.0 1e-06 
0.0 -0.0947000000002 0 2.0 1e-06 
0.0 -0.0946000000002 0 2.0 1e-06 
0.0 -0.0945000000002 0 2.0 1e-06 
0.0 -0.0944000000002 0 2.0 1e-06 
0.0 -0.0943000000002 0 2.0 1e-06 
0.0 -0.0942000000002 0 2.0 1e-06 
0.0 -0.0941000000002 0 2.0 1e-06 
0.0 -0.0940000000002 0 2.0 1e-06 
0.0 -0.0939000000002 0 2.0 1e-06 
0.0 -0.0938000000002 0 2.0 1e-06 
0.0 -0.0937000000002 0 2.0 1e-06 
0.0 -0.0936000000002 0 2.0 1e-06 
0.0 -0.0935000000002 0 2.0 1e-06 
0.0 -0.0934000000002 0 2.0 1e-06 
0.0 -0.0933000000002 0 2.0 1e-06 
0.0 -0.0932000000002 0 2.0 1e-06 
0.0 -0.0931000000002 0 2.0 1e-06 
0.0 -0.0930000000002 0 2.0 1e-06 
0.0 -0.0929000000002 0 2.0 1e-06 
0.0 -0.0928000000002 0 2.0 1e-06 
0.0 -0.0927000000002 0 2.0 1e-06 
0.0 -0.0926000000002 0 2.0 1e-06 
0.0 -0.0925000000002 0 2.0 1e-06 
0.0 -0.0924000000002 0 2.0 1e-06 
0.0 -0.0923000000002 0 2.0 1e-06 
0.0 -0.0922000000002 0 2.0 1e-06 
0.0 -0.0921000000002 0 2.0 1e-06 
0.0 -0.0920000000002 0 2.0 1e-06 
0.0 -0.0919000000002 0 2.0 1e-06 
0.0 -0.0918000000002 0 2.0 1e-06 
0.0 -0.0917000000002 0 2.0 1e-06 
0.0 -0.0916000000002 0 2.0 1e-06 
0.0 -0.0915000000002 0 2.0 1e-06 
0.0 -0.0914000000002 0 2.0 1e-06 
0.0 -0.0913000000002 0 2.0 1e-06 
0.0 -0.0912000000002 0 2.0 1e-06 
0.0 -0.0911000000002 0 2.0 1e-06 
0.0 -0.0910000000002 0 2.0 1e-06 
0.0 -0.0909000000002 0 2.0 1e-06 
0.0 -0.0908000000002 0 2.0 1e-06 
0.0 -0.0907000000002 0 2.0 1e-06 
0.0 -0.0906000000002 0 2.0 1e-06 
0.0 -0.0905000000002 0 2.0 1e-06 
0.0 -0.0904000000002 0 2.0 1e-06 
0.0 -0.0903000000002 0 2.0 1e-06 
0.0 -0.0902000000002 0 2.0 1e-06 
0.0 -0.0901000000002 0 2.0 1e-06 
0.0 -0.0900000000002 0 2.0 1e-06 
0.0 -0.0899000000002 0 2.0 1e-06 
0.0 -0.0898000000002 0 2.0 1e-06 
0.0 -0.0897000000002 0 2.0 1e-06 
0.0 -0.0896000000002 0 2.0 1e-06 
0.0 -0.0895000000002 0 2.0 1e-06 
0.0 -0.0894000000002 0 2.0 1e-06 
0.0 -0.0893000000002 0 2.0 1e-06 
0.0 -0.0892000000002 0 2.0 1e-06 
0.0 -0.0891000000002 0 2.0 1e-06 
0.0 -0.0890000000002 0 2.0 1e-06 
0.0 -0.0889000000002 0 2.0 1e-06 
0.0 -0.0888000000002 0 2.0 1e-06 
0.0 -0.0887000000002 0 2.0 1e-06 
0.0 -0.0886000000002 0 2.0 1e-06 
0.0 -0.0885000000002 0 2.0 1e-06 
0.0 -0.0884000000002 0 2.0 1e-06 
0.0 -0.0883000000002 0 2.0 1e-06 
0.0 -0.0882000000002 0 2.0 1e-06 
0.0 -0.0881000000002 0 2.0 1e-06 
0.0 -0.0880000000002 0 2.0 1e-06 
0.0 -0.0879000000002 0 2.0 1e-06 
0.0 -0.0878000000002 0 2.0 1e-06 
0.0 -0.0877000000002 0 2.0 1e-06 
0.0 -0.0876000000002 0 2.0 1e-06 
0.0 -0.0875000000002 0 2.0 1e-06 
0.0 -0.0874000000002 0 2.0 1e-06 
0.0 -0.0873000000002 0 2.0 1e-06 
0.0 -0.0872000000002 0 2.0 1e-06 
0.0 -0.0871000000002 0 2.0 1e-06 
0.0 -0.0870000000002 0 2.0 1e-06 
0.0 -0.0869000000002 0 2.0 1e-06 
0.0 -0.0868000000002 0 2.0 1e-06 
0.0 -0.0867000000002 0 2.0 1e-06 
0.0 -0.0866000000002 0 2.0 1e-06 
0.0 -0.0865000000002 0 2.0 1e-06 
0.0 -0.0864000000002 0 2.0 1e-06 
0.0 -0.0863000000002 0 2.0 1e-06 
0.0 -0.0862000000002 0 2.0 1e-06 
0.0 -0.0861000000002 0 2.0 1e-06 
0.0 -0.0860000000002 0 2.0 1e-06 
0.0 -0.0859000000002 0 2.0 1e-06 
0.0 -0.0858000000002 0 2.0 1e-06 
0.0 -0.0857000000002 0 2.0 1e-06 
0.0 -0.0856000000002 0 2.0 1e-06 
0.0 -0.0855000000002 0 2.0 1e-06 
0.0 -0.0854000000002 0 2.0 1e-06 
0.0 -0.0853000000002 0 2.0 1e-06 
0.0 -0.0852000000002 0 2.0 1e-06 
0.0 -0.0851000000002 0 2.0 1e-06 
0.0 -0.0850000000002 0 2.0 1e-06 
0.0 -0.0849000000002 0 2.0 1e-06 
0.0 -0.0848000000002 0 2.0 1e-06 
0.0 -0.0847000000002 0 2.0 1e-06 
0.0 -0.0846000000002 0 2.0 1e-06 
0.0 -0.0845000000002 0 2.0 1e-06 
0.0 -0.0844000000002 0 2.0 1e-06 
0.0 -0.0843000000002 0 2.0 1e-06 
0.0 -0.0842000000002 0 2.0 1e-06 
0.0 -0.0841000000002 0 2.0 1e-06 
0.0 -0.0840000000002 0 2.0 1e-06 
0.0 -0.0839000000002 0 2.0 1e-06 
0.0 -0.0838000000002 0 2.0 1e-06 
0.0 -0.0837000000002 0 2.0 1e-06 
0.0 -0.0836000000002 0 2.0 1e-06 
0.0 -0.0835000000002 0 2.0 1e-06 
0.0 -0.0834000000002 0 2.0 1e-06 
0.0 -0.0833000000002 0 2.0 1e-06 
0.0 -0.0832000000002 0 2.0 1e-06 
0.0 -0.0831000000002 0 2.0 1e-06 
0.0 -0.0830000000002 0 2.0 1e-06 
0.0 -0.0829000000002 0 2.0 1e-06 
0.0 -0.0828000000002 0 2.0 1e-06 
0.0 -0.0827000000002 0 2.0 1e-06 
0.0 -0.0826000000002 0 2.0 1e-06 
0.0 -0.0825000000002 0 2.0 1e-06 
0.0 -0.0824000000002 0 2.0 1e-06 
0.0 -0.0823000000002 0 2.0 1e-06 
0.0 -0.0822000000002 0 2.0 1e-06 
0.0 -0.0821000000002 0 2.0 1e-06 
0.0 -0.0820000000002 0 2.0 1e-06 
0.0 -0.0819000000002 0 2.0 1e-06 
0.0 -0.0818000000002 0 2.0 1e-06 
0.0 -0.0817000000002 0 2.0 1e-06 
0.0 -0.0816000000002 0 2.0 1e-06 
0.0 -0.0815000000002 0 2.0 1e-06 
0.0 -0.0814000000002 0 2.0 1e-06 
0.0 -0.0813000000002 0 2.0 1e-06 
0.0 -0.0812000000002 0 2.0 1e-06 
0.0 -0.0811000000002 0 2.0 1e-06 
0.0 -0.0810000000002 0 2.0 1e-06 
0.0 -0.0809000000002 0 2.0 1e-06 
0.0 -0.0808000000002 0 2.0 1e-06 
0.0 -0.0807000000002 0 2.0 1e-06 
0.0 -0.0806000000002 0 2.0 1e-06 
0.0 -0.0805000000002 0 2.0 1e-06 
0.0 -0.0804000000002 0 2.0 1e-06 
0.0 -0.0803000000002 0 2.0 1e-06 
0.0 -0.0802000000002 0 2.0 1e-06 
0.0 -0.0801000000002 0 2.0 1e-06 
0.0 -0.0800000000002 0 2.0 1e-06 
0.0 -0.0799000000002 0 2.0 1e-06 
0.0 -0.0798000000002 0 2.0 1e-06 
0.0 -0.0797000000002 0 2.0 1e-06 
0.0 -0.0796000000002 0 2.0 1e-06 
0.0 -0.0795000000002 0 2.0 1e-06 
0.0 -0.0794000000002 0 2.0 1e-06 
0.0 -0.0793000000002 0 2.0 1e-06 
0.0 -0.0792000000002 0 2.0 1e-06 
0.0 -0.0791000000002 0 2.0 1e-06 
0.0 -0.0790000000002 0 2.0 1e-06 
0.0 -0.0789000000002 0 2.0 1e-06 
0.0 -0.0788000000002 0 2.0 1e-06 
0.0 -0.0787000000002 0 2.0 1e-06 
0.0 -0.0786000000002 0 2.0 1e-06 
0.0 -0.0785000000002 0 2.0 1e-06 
0.0 -0.0784000000002 0 2.0 1e-06 
0.0 -0.0783000000002 0 2.0 1e-06 
0.0 -0.0782000000002 0 2.0 1e-06 
0.0 -0.0781000000002 0 2.0 1e-06 
0.0 -0.0780000000002 0 2.0 1e-06 
0.0 -0.0779000000002 0 2.0 1e-06 
0.0 -0.0778000000002 0 2.0 1e-06 
0.0 -0.0777000000002 0 2.0 1e-06 
0.0 -0.0776000000002 0 2.0 1e-06 
0.0 -0.0775000000002 0 2.0 1e-06 
0.0 -0.0774000000002 0 2.0 1e-06 
0.0 -0.0773000000002 0 2.0 1e-06 
0.0 -0.0772000000002 0 2.0 1e-06 
0.0 -0.0771000000002 0 2.0 1e-06 
0.0 -0.0770000000002 0 2.0 1e-06 
0.0 -0.0769000000002 0 2.0 1e-06 
0.0 -0.0768000000002 0 2.0 1e-06 
0.0 -0.0767000000002 0 2.0 1e-06 
0.0 -0.0766000000002 0 2.0 1e-06 
0.0 -0.0765000000002 0 2.0 1e-06 
0.0 -0.0764000000002 0 2.0 1e-06 
0.0 -0.0763000000002 0 2.0 1e-06 
0.0 -0.0762000000002 0 2.0 1e-06 
0.0 -0.0761000000002 0 2.0 1e-06 
0.0 -0.0760000000002 0 2.0 1e-06 
0.0 -0.0759000000002 0 2.0 1e-06 
0.0 -0.0758000000002 0 2.0 1e-06 
0.0 -0.0757000000002 0 2.0 1e-06 
0.0 -0.0756000000002 0 2.0 1e-06 
0.0 -0.0755000000002 0 2.0 1e-06 
0.0 -0.0754000000002 0 2.0 1e-06 
0.0 -0.0753000000002 0 2.0 1e-06 
0.0 -0.0752000000002 0 2.0 1e-06 
0.0 -0.0751000000002 0 2.0 1e-06 
0.0 -0.0750000000002 0 2.0 1e-06 
0.0 -0.0749000000002 0 2.0 1e-06 
0.0 -0.0748000000002 0 2.0 1e-06 
0.0 -0.0747000000002 0 2.0 1e-06 
0.0 -0.0746000000002 0 2.0 1e-06 
0.0 -0.0745000000002 0 2.0 1e-06 
0.0 -0.0744000000002 0 2.0 1e-06 
0.0 -0.0743000000002 0 2.0 1e-06 
0.0 -0.0742000000002 0 2.0 1e-06 
0.0 -0.0741000000002 0 2.0 1e-06 
0.0 -0.0740000000002 0 2.0 1e-06 
0.0 -0.0739000000002 0 2.0 1e-06 
0.0 -0.0738000000002 0 2.0 1e-06 
0.0 -0.0737000000002 0 2.0 1e-06 
0.0 -0.0736000000002 0 2.0 1e-06 
0.0 -0.0735000000002 0 2.0 1e-06 
0.0 -0.0734000000002 0 2.0 1e-06 
0.0 -0.0733000000002 0 2.0 1e-06 
0.0 -0.0732000000002 0 2.0 1e-06 
0.0 -0.0731000000002 0 2.0 1e-06 
0.0 -0.0730000000002 0 2.0 1e-06 
0.0 -0.0729000000002 0 2.0 1e-06 
0.0 -0.0728000000002 0 2.0 1e-06 
0.0 -0.0727000000002 0 2.0 1e-06 
0.0 -0.0726000000002 0 2.0 1e-06 
0.0 -0.0725000000002 0 2.0 1e-06 
0.0 -0.0724000000002 0 2.0 1e-06 
0.0 -0.0723000000002 0 2.0 1e-06 
0.0 -0.0722000000002 0 2.0 1e-06 
0.0 -0.0721000000002 0 2.0 1e-06 
0.0 -0.0720000000002 0 2.0 1e-06 
0.0 -0.0719000000002 0 2.0 1e-06 
0.0 -0.0718000000002 0 2.0 1e-06 
0.0 -0.0717000000002 0 2.0 1e-06 
0.0 -0.0716000000002 0 2.0 1e-06 
0.0 -0.0715000000002 0 2.0 1e-06 
0.0 -0.0714000000002 0 2.0 1e-06 
0.0 -0.0713000000002 0 2.0 1e-06 
0.0 -0.0712000000002 0 2.0 1e-06 
0.0 -0.0711000000002 0 2.0 1e-06 
0.0 -0.0710000000002 0 2.0 1e-06 
0.0 -0.0709000000002 0 2.0 1e-06 
0.0 -0.0708000000002 0 2.0 1e-06 
0.0 -0.0707000000002 0 2.0 1e-06 
0.0 -0.0706000000002 0 2.0 1e-06 
0.0 -0.0705000000002 0 2.0 1e-06 
0.0 -0.0704000000002 0 2.0 1e-06 
0.0 -0.0703000000002 0 2.0 1e-06 
0.0 -0.0702000000002 0 2.0 1e-06 
0.0 -0.0701000000002 0 2.0 1e-06 
0.0 -0.0700000000002 0 2.0 1e-06 
0.0 -0.0699000000002 0 2.0 1e-06 
0.0 -0.0698000000002 0 2.0 1e-06 
0.0 -0.0697000000002 0 2.0 1e-06 
0.0 -0.0696000000002 0 2.0 1e-06 
0.0 -0.0695000000002 0 2.0 1e-06 
0.0 -0.0694000000002 0 2.0 1e-06 
0.0 -0.0693000000002 0 2.0 1e-06 
0.0 -0.0692000000002 0 2.0 1e-06 
0.0 -0.0691000000002 0 2.0 1e-06 
0.0 -0.0690000000002 0 2.0 1e-06 
0.0 -0.0689000000002 0 2.0 1e-06 
0.0 -0.0688000000002 0 2.0 1e-06 
0.0 -0.0687000000002 0 2.0 1e-06 
0.0 -0.0686000000002 0 2.0 1e-06 
0.0 -0.0685000000002 0 2.0 1e-06 
0.0 -0.0684000000002 0 2.0 1e-06 
0.0 -0.0683000000002 0 2.0 1e-06 
0.0 -0.0682000000002 0 2.0 1e-06 
0.0 -0.0681000000002 0 2.0 1e-06 
0.0 -0.0680000000002 0 2.0 1e-06 
0.0 -0.0679000000002 0 2.0 1e-06 
0.0 -0.0678000000002 0 2.0 1e-06 
0.0 -0.0677000000002 0 2.0 1e-06 
0.0 -0.0676000000002 0 2.0 1e-06 
0.0 -0.0675000000002 0 2.0 1e-06 
0.0 -0.0674000000002 0 2.0 1e-06 
0.0 -0.0673000000002 0 2.0 1e-06 
0.0 -0.0672000000002 0 2.0 1e-06 
0.0 -0.0671000000002 0 2.0 1e-06 
0.0 -0.0670000000002 0 2.0 1e-06 
0.0 -0.0669000000002 0 2.0 1e-06 
0.0 -0.0668000000002 0 2.0 1e-06 
0.0 -0.0667000000002 0 2.0 1e-06 
0.0 -0.0666000000002 0 2.0 1e-06 
0.0 -0.0665000000002 0 2.0 1e-06 
0.0 -0.0664000000002 0 2.0 1e-06 
0.0 -0.0663000000002 0 2.0 1e-06 
0.0 -0.0662000000002 0 2.0 1e-06 
0.0 -0.0661000000002 0 2.0 1e-06 
0.0 -0.0660000000002 0 2.0 1e-06 
0.0 -0.0659000000002 0 2.0 1e-06 
0.0 -0.0658000000002 0 2.0 1e-06 
0.0 -0.0657000000002 0 2.0 1e-06 
0.0 -0.0656000000002 0 2.0 1e-06 
0.0 -0.0655000000002 0 2.0 1e-06 
0.0 -0.0654000000002 0 2.0 1e-06 
0.0 -0.0653000000002 0 2.0 1e-06 
0.0 -0.0652000000002 0 2.0 1e-06 
0.0 -0.0651000000002 0 2.0 1e-06 
0.0 -0.0650000000002 0 2.0 1e-06 
0.0 -0.0649000000002 0 2.0 1e-06 
0.0 -0.0648000000002 0 2.0 1e-06 
0.0 -0.0647000000002 0 2.0 1e-06 
0.0 -0.0646000000002 0 2.0 1e-06 
0.0 -0.0645000000002 0 2.0 1e-06 
0.0 -0.0644000000002 0 2.0 1e-06 
0.0 -0.0643000000002 0 2.0 1e-06 
0.0 -0.0642000000002 0 2.0 1e-06 
0.0 -0.0641000000002 0 2.0 1e-06 
0.0 -0.0640000000002 0 2.0 1e-06 
0.0 -0.0639000000002 0 2.0 1e-06 
0.0 -0.0638000000002 0 2.0 1e-06 
0.0 -0.0637000000002 0 2.0 1e-06 
0.0 -0.0636000000002 0 2.0 1e-06 
0.0 -0.0635000000002 0 2.0 1e-06 
0.0 -0.0634000000002 0 2.0 1e-06 
0.0 -0.0633000000002 0 2.0 1e-06 
0.0 -0.0632000000002 0 2.0 1e-06 
0.0 -0.0631000000002 0 2.0 1e-06 
0.0 -0.0630000000002 0 2.0 1e-06 
0.0 -0.0629000000002 0 2.0 1e-06 
0.0 -0.0628000000002 0 2.0 1e-06 
0.0 -0.0627000000002 0 2.0 1e-06 
0.0 -0.0626000000002 0 2.0 1e-06 
0.0 -0.0625000000002 0 2.0 1e-06 
0.0 -0.0624000000002 0 2.0 1e-06 
0.0 -0.0623000000002 0 2.0 1e-06 
0.0 -0.0622000000002 0 2.0 1e-06 
0.0 -0.0621000000002 0 2.0 1e-06 
0.0 -0.0620000000002 0 2.0 1e-06 
0.0 -0.0619000000002 0 2.0 1e-06 
0.0 -0.0618000000002 0 2.0 1e-06 
0.0 -0.0617000000002 0 2.0 1e-06 
0.0 -0.0616000000002 0 2.0 1e-06 
0.0 -0.0615000000002 0 2.0 1e-06 
0.0 -0.0614000000002 0 2.0 1e-06 
0.0 -0.0613000000002 0 2.0 1e-06 
0.0 -0.0612000000002 0 2.0 1e-06 
0.0 -0.0611000000002 0 2.0 1e-06 
0.0 -0.0610000000002 0 2.0 1e-06 
0.0 -0.0609000000002 0 2.0 1e-06 
0.0 -0.0608000000002 0 2.0 1e-06 
0.0 -0.0607000000002 0 2.0 1e-06 
0.0 -0.0606000000002 0 2.0 1e-06 
0.0 -0.0605000000002 0 2.0 1e-06 
0.0 -0.0604000000002 0 2.0 1e-06 
0.0 -0.0603000000002 0 2.0 1e-06 
0.0 -0.0602000000002 0 2.0 1e-06 
0.0 -0.0601000000002 0 2.0 1e-06 
0.0 -0.0600000000002 0 2.0 1e-06 
0.0 -0.0599000000002 0 2.0 1e-06 
0.0 -0.0598000000002 0 2.0 1e-06 
0.0 -0.0597000000002 0 2.0 1e-06 
0.0 -0.0596000000002 0 2.0 1e-06 
0.0 -0.0595000000002 0 2.0 1e-06 
0.0 -0.0594000000002 0 2.0 1e-06 
0.0 -0.0593000000002 0 2.0 1e-06 
0.0 -0.0592000000002 0 2.0 1e-06 
0.0 -0.0591000000002 0 2.0 1e-06 
0.0 -0.0590000000002 0 2.0 1e-06 
0.0 -0.0589000000002 0 2.0 1e-06 
0.0 -0.0588000000002 0 2.0 1e-06 
0.0 -0.0587000000002 0 2.0 1e-06 
0.0 -0.0586000000002 0 2.0 1e-06 
0.0 -0.0585000000002 0 2.0 1e-06 
0.0 -0.0584000000002 0 2.0 1e-06 
0.0 -0.0583000000002 0 2.0 1e-06 
0.0 -0.0582000000002 0 2.0 1e-06 
0.0 -0.0581000000002 0 2.0 1e-06 
0.0 -0.0580000000002 0 2.0 1e-06 
0.0 -0.0579000000002 0 2.0 1e-06 
0.0 -0.0578000000002 0 2.0 1e-06 
0.0 -0.0577000000002 0 2.0 1e-06 
0.0 -0.0576000000002 0 2.0 1e-06 
0.0 -0.0575000000002 0 2.0 1e-06 
0.0 -0.0574000000002 0 2.0 1e-06 
0.0 -0.0573000000002 0 2.0 1e-06 
0.0 -0.0572000000002 0 2.0 1e-06 
0.0 -0.0571000000002 0 2.0 1e-06 
0.0 -0.0570000000002 0 2.0 1e-06 
0.0 -0.0569000000002 0 2.0 1e-06 
0.0 -0.0568000000002 0 2.0 1e-06 
0.0 -0.0567000000002 0 2.0 1e-06 
0.0 -0.0566000000002 0 2.0 1e-06 
0.0 -0.0565000000002 0 2.0 1e-06 
0.0 -0.0564000000002 0 2.0 1e-06 
0.0 -0.0563000000002 0 2.0 1e-06 
0.0 -0.0562000000002 0 2.0 1e-06 
0.0 -0.0561000000002 0 2.0 1e-06 
0.0 -0.0560000000002 0 2.0 1e-06 
0.0 -0.0559000000002 0 2.0 1e-06 
0.0 -0.0558000000002 0 2.0 1e-06 
0.0 -0.0557000000002 0 2.0 1e-06 
0.0 -0.0556000000002 0 2.0 1e-06 
0.0 -0.0555000000002 0 2.0 1e-06 
0.0 -0.0554000000002 0 2.0 1e-06 
0.0 -0.0553000000002 0 2.0 1e-06 
0.0 -0.0552000000002 0 2.0 1e-06 
0.0 -0.0551000000002 0 2.0 1e-06 
0.0 -0.0550000000002 0 2.0 1e-06 
0.0 -0.0549000000002 0 2.0 1e-06 
0.0 -0.0548000000002 0 2.0 1e-06 
0.0 -0.0547000000002 0 2.0 1e-06 
0.0 -0.0546000000002 0 2.0 1e-06 
0.0 -0.0545000000002 0 2.0 1e-06 
0.0 -0.0544000000002 0 2.0 1e-06 
0.0 -0.0543000000002 0 2.0 1e-06 
0.0 -0.0542000000002 0 2.0 1e-06 
0.0 -0.0541000000002 0 2.0 1e-06 
0.0 -0.0540000000002 0 2.0 1e-06 
0.0 -0.0539000000002 0 2.0 1e-06 
0.0 -0.0538000000002 0 2.0 1e-06 
0.0 -0.0537000000002 0 2.0 1e-06 
0.0 -0.0536000000002 0 2.0 1e-06 
0.0 -0.0535000000002 0 2.0 1e-06 
0.0 -0.0534000000002 0 2.0 1e-06 
0.0 -0.0533000000002 0 2.0 1e-06 
0.0 -0.0532000000002 0 2.0 1e-06 
0.0 -0.0531000000002 0 2.0 1e-06 
0.0 -0.0530000000002 0 2.0 1e-06 
0.0 -0.0529000000002 0 2.0 1e-06 
0.0 -0.0528000000002 0 2.0 1e-06 
0.0 -0.0527000000002 0 2.0 1e-06 
0.0 -0.0526000000002 0 2.0 1e-06 
0.0 -0.0525000000002 0 2.0 1e-06 
0.0 -0.0524000000002 0 2.0 1e-06 
0.0 -0.0523000000002 0 2.0 1e-06 
0.0 -0.0522000000002 0 2.0 1e-06 
0.0 -0.0521000000002 0 2.0 1e-06 
0.0 -0.0520000000002 0 2.0 1e-06 
0.0 -0.0519000000002 0 2.0 1e-06 
0.0 -0.0518000000002 0 2.0 1e-06 
0.0 -0.0517000000002 0 2.0 1e-06 
0.0 -0.0516000000002 0 2.0 1e-06 
0.0 -0.0515000000002 0 2.0 1e-06 
0.0 -0.0514000000002 0 2.0 1e-06 
0.0 -0.0513000000002 0 2.0 1e-06 
0.0 -0.0512000000002 0 2.0 1e-06 
0.0 -0.0511000000002 0 2.0 1e-06 
0.0 -0.0510000000002 0 2.0 1e-06 
0.0 -0.0509000000002 0 2.0 1e-06 
0.0 -0.0508000000002 0 2.0 1e-06 
0.0 -0.0507000000002 0 2.0 1e-06 
0.0 -0.0506000000002 0 2.0 1e-06 
0.0 -0.0505000000002 0 2.0 1e-06 
0.0 -0.0504000000002 0 2.0 1e-06 
0.0 -0.0503000000002 0 2.0 1e-06 
0.0 -0.0502000000002 0 2.0 1e-06 
0.0 -0.0501000000002 0 2.0 1e-06 
0.0 -0.0500000000002 0 2.0 1e-06 
0.0 -0.0499000000002 0 2.0 1e-06 
0.0 -0.0498000000002 0 2.0 1e-06 
0.0 -0.0497000000002 0 2.0 1e-06 
0.0 -0.0496000000002 0 2.0 1e-06 
0.0 -0.0495000000002 0 2.0 1e-06 
0.0 -0.0494000000002 0 2.0 1e-06 
0.0 -0.0493000000002 0 2.0 1e-06 
0.0 -0.0492000000002 0 2.0 1e-06 
0.0 -0.0491000000002 0 2.0 1e-06 
0.0 -0.0490000000002 0 2.0 1e-06 
0.0 -0.0489000000002 0 2.0 1e-06 
0.0 -0.0488000000002 0 2.0 1e-06 
0.0 -0.0487000000002 0 2.0 1e-06 
0.0 -0.0486000000002 0 2.0 1e-06 
0.0 -0.0485000000002 0 2.0 1e-06 
0.0 -0.0484000000002 0 2.0 1e-06 
0.0 -0.0483000000002 0 2.0 1e-06 
0.0 -0.0482000000002 0 2.0 1e-06 
0.0 -0.0481000000002 0 2.0 1e-06 
0.0 -0.0480000000002 0 2.0 1e-06 
0.0 -0.0479000000002 0 2.0 1e-06 
0.0 -0.0478000000002 0 2.0 1e-06 
0.0 -0.0477000000002 0 2.0 1e-06 
0.0 -0.0476000000002 0 2.0 1e-06 
0.0 -0.0475000000002 0 2.0 1e-06 
0.0 -0.0474000000002 0 2.0 1e-06 
0.0 -0.0473000000002 0 2.0 1e-06 
0.0 -0.0472000000002 0 2.0 1e-06 
0.0 -0.0471000000002 0 2.0 1e-06 
0.0 -0.0470000000002 0 2.0 1e-06 
0.0 -0.0469000000002 0 2.0 1e-06 
0.0 -0.0468000000002 0 2.0 1e-06 
0.0 -0.0467000000002 0 2.0 1e-06 
0.0 -0.0466000000002 0 2.0 1e-06 
0.0 -0.0465000000002 0 2.0 1e-06 
0.0 -0.0464000000002 0 2.0 1e-06 
0.0 -0.0463000000002 0 2.0 1e-06 
0.0 -0.0462000000002 0 2.0 1e-06 
0.0 -0.0461000000002 0 2.0 1e-06 
0.0 -0.0460000000002 0 2.0 1e-06 
0.0 -0.0459000000002 0 2.0 1e-06 
0.0 -0.0458000000002 0 2.0 1e-06 
0.0 -0.0457000000002 0 2.0 1e-06 
0.0 -0.0456000000002 0 2.0 1e-06 
0.0 -0.0455000000002 0 2.0 1e-06 
0.0 -0.0454000000002 0 2.0 1e-06 
0.0 -0.0453000000002 0 2.0 1e-06 
0.0 -0.0452000000002 0 2.0 1e-06 
0.0 -0.0451000000002 0 2.0 1e-06 
0.0 -0.0450000000002 0 2.0 1e-06 
0.0 -0.0449000000002 0 2.0 1e-06 
0.0 -0.0448000000002 0 2.0 1e-06 
0.0 -0.0447000000002 0 2.0 1e-06 
0.0 -0.0446000000002 0 2.0 1e-06 
0.0 -0.0445000000002 0 2.0 1e-06 
0.0 -0.0444000000002 0 2.0 1e-06 
0.0 -0.0443000000002 0 2.0 1e-06 
0.0 -0.0442000000002 0 2.0 1e-06 
0.0 -0.0441000000002 0 2.0 1e-06 
0.0 -0.0440000000002 0 2.0 1e-06 
0.0 -0.0439000000002 0 2.0 1e-06 
0.0 -0.0438000000002 0 2.0 1e-06 
0.0 -0.0437000000002 0 2.0 1e-06 
0.0 -0.0436000000002 0 2.0 1e-06 
0.0 -0.0435000000002 0 2.0 1e-06 
0.0 -0.0434000000002 0 2.0 1e-06 
0.0 -0.0433000000002 0 2.0 1e-06 
0.0 -0.0432000000002 0 2.0 1e-06 
0.0 -0.0431000000002 0 2.0 1e-06 
0.0 -0.0430000000002 0 2.0 1e-06 
0.0 -0.0429000000002 0 2.0 1e-06 
0.0 -0.0428000000002 0 2.0 1e-06 
0.0 -0.0427000000002 0 2.0 1e-06 
0.0 -0.0426000000002 0 2.0 1e-06 
0.0 -0.0425000000002 0 2.0 1e-06 
0.0 -0.0424000000002 0 2.0 1e-06 
0.0 -0.0423000000002 0 2.0 1e-06 
0.0 -0.0422000000002 0 2.0 1e-06 
0.0 -0.0421000000002 0 2.0 1e-06 
0.0 -0.0420000000002 0 2.0 1e-06 
0.0 -0.0419000000002 0 2.0 1e-06 
0.0 -0.0418000000002 0 2.0 1e-06 
0.0 -0.0417000000002 0 2.0 1e-06 
0.0 -0.0416000000002 0 2.0 1e-06 
0.0 -0.0415000000002 0 2.0 1e-06 
0.0 -0.0414000000002 0 2.0 1e-06 
0.0 -0.0413000000002 0 2.0 1e-06 
0.0 -0.0412000000002 0 2.0 1e-06 
0.0 -0.0411000000002 0 2.0 1e-06 
0.0 -0.0410000000002 0 2.0 1e-06 
0.0 -0.0409000000002 0 2.0 1e-06 
0.0 -0.0408000000002 0 2.0 1e-06 
0.0 -0.0407000000002 0 2.0 1e-06 
0.0 -0.0406000000002 0 2.0 1e-06 
0.0 -0.0405000000002 0 2.0 1e-06 
0.0 -0.0404000000002 0 2.0 1e-06 
0.0 -0.0403000000002 0 2.0 1e-06 
0.0 -0.0402000000002 0 2.0 1e-06 
0.0 -0.0401000000002 0 2.0 1e-06 
0.0 -0.0400000000002 0 2.0 1e-06 
0.0 -0.0399000000002 0 2.0 1e-06 
0.0 -0.0398000000002 0 2.0 1e-06 
0.0 -0.0397000000002 0 2.0 1e-06 
0.0 -0.0396000000002 0 2.0 1e-06 
0.0 -0.0395000000002 0 2.0 1e-06 
0.0 -0.0394000000002 0 2.0 1e-06 
0.0 -0.0393000000002 0 2.0 1e-06 
0.0 -0.0392000000002 0 2.0 1e-06 
0.0 -0.0391000000002 0 2.0 1e-06 
0.0 -0.0390000000002 0 2.0 1e-06 
0.0 -0.0389000000002 0 2.0 1e-06 
0.0 -0.0388000000002 0 2.0 1e-06 
0.0 -0.0387000000002 0 2.0 1e-06 
0.0 -0.0386000000002 0 2.0 1e-06 
0.0 -0.0385000000002 0 2.0 1e-06 
0.0 -0.0384000000002 0 2.0 1e-06 
0.0 -0.0383000000002 0 2.0 1e-06 
0.0 -0.0382000000002 0 2.0 1e-06 
0.0 -0.0381000000002 0 2.0 1e-06 
0.0 -0.0380000000002 0 2.0 1e-06 
0.0 -0.0379000000002 0 2.0 1e-06 
0.0 -0.0378000000002 0 2.0 1e-06 
0.0 -0.0377000000002 0 2.0 1e-06 
0.0 -0.0376000000002 0 2.0 1e-06 
0.0 -0.0375000000002 0 2.0 1e-06 
0.0 -0.0374000000002 0 2.0 1e-06 
0.0 -0.0373000000002 0 2.0 1e-06 
0.0 -0.0372000000002 0 2.0 1e-06 
0.0 -0.0371000000002 0 2.0 1e-06 
0.0 -0.0370000000002 0 2.0 1e-06 
0.0 -0.0369000000002 0 2.0 1e-06 
0.0 -0.0368000000002 0 2.0 1e-06 
0.0 -0.0367000000002 0 2.0 1e-06 
0.0 -0.0366000000002 0 2.0 1e-06 
0.0 -0.0365000000002 0 2.0 1e-06 
0.0 -0.0364000000002 0 2.0 1e-06 
0.0 -0.0363000000002 0 2.0 1e-06 
0.0 -0.0362000000002 0 2.0 1e-06 
0.0 -0.0361000000002 0 2.0 1e-06 
0.0 -0.0360000000002 0 2.0 1e-06 
0.0 -0.0359000000002 0 2.0 1e-06 
0.0 -0.0358000000002 0 2.0 1e-06 
0.0 -0.0357000000002 0 2.0 1e-06 
0.0 -0.0356000000002 0 2.0 1e-06 
0.0 -0.0355000000002 0 2.0 1e-06 
0.0 -0.0354000000002 0 2.0 1e-06 
0.0 -0.0353000000002 0 2.0 1e-06 
0.0 -0.0352000000002 0 2.0 1e-06 
0.0 -0.0351000000002 0 2.0 1e-06 
0.0 -0.0350000000002 0 2.0 1e-06 
0.0 -0.0349000000002 0 2.0 1e-06 
0.0 -0.0348000000002 0 2.0 1e-06 
0.0 -0.0347000000002 0 2.0 1e-06 
0.0 -0.0346000000002 0 2.0 1e-06 
0.0 -0.0345000000002 0 2.0 1e-06 
0.0 -0.0344000000002 0 2.0 1e-06 
0.0 -0.0343000000002 0 2.0 1e-06 
0.0 -0.0342000000002 0 2.0 1e-06 
0.0 -0.0341000000002 0 2.0 1e-06 
0.0 -0.0340000000002 0 2.0 1e-06 
0.0 -0.0339000000002 0 2.0 1e-06 
0.0 -0.0338000000002 0 2.0 1e-06 
0.0 -0.0337000000002 0 2.0 1e-06 
0.0 -0.0336000000002 0 2.0 1e-06 
0.0 -0.0335000000002 0 2.0 1e-06 
0.0 -0.0334000000002 0 2.0 1e-06 
0.0 -0.0333000000002 0 2.0 1e-06 
0.0 -0.0332000000002 0 2.0 1e-06 
0.0 -0.0331000000002 0 2.0 1e-06 
0.0 -0.0330000000002 0 2.0 1e-06 
0.0 -0.0329000000002 0 2.0 1e-06 
0.0 -0.0328000000002 0 2.0 1e-06 
0.0 -0.0327000000002 0 2.0 1e-06 
0.0 -0.0326000000002 0 2.0 1e-06 
0.0 -0.0325000000002 0 2.0 1e-06 
0.0 -0.0324000000002 0 2.0 1e-06 
0.0 -0.0323000000002 0 2.0 1e-06 
0.0 -0.0322000000002 0 2.0 1e-06 
0.0 -0.0321000000002 0 2.0 1e-06 
0.0 -0.0320000000002 0 2.0 1e-06 
0.0 -0.0319000000002 0 2.0 1e-06 
0.0 -0.0318000000002 0 2.0 1e-06 
0.0 -0.0317000000002 0 2.0 1e-06 
0.0 -0.0316000000002 0 2.0 1e-06 
0.0 -0.0315000000002 0 2.0 1e-06 
0.0 -0.0314000000002 0 2.0 1e-06 
0.0 -0.0313000000002 0 2.0 1e-06 
0.0 -0.0312000000002 0 2.0 1e-06 
0.0 -0.0311000000002 0 2.0 1e-06 
0.0 -0.0310000000002 0 2.0 1e-06 
0.0 -0.0309000000002 0 2.0 1e-06 
0.0 -0.0308000000002 0 2.0 1e-06 
0.0 -0.0307000000002 0 2.0 1e-06 
0.0 -0.0306000000002 0 2.0 1e-06 
0.0 -0.0305000000002 0 2.0 1e-06 
0.0 -0.0304000000002 0 2.0 1e-06 
0.0 -0.0303000000002 0 2.0 1e-06 
0.0 -0.0302000000002 0 2.0 1e-06 
0.0 -0.0301000000002 0 2.0 1e-06 
0.0 -0.0300000000002 0 2.0 1e-06 
0.0 -0.0299000000002 0 2.0 1e-06 
0.0 -0.0298000000002 0 2.0 1e-06 
0.0 -0.0297000000002 0 2.0 1e-06 
0.0 -0.0296000000002 0 2.0 1e-06 
0.0 -0.0295000000002 0 2.0 1e-06 
0.0 -0.0294000000002 0 2.0 1e-06 
0.0 -0.0293000000002 0 2.0 1e-06 
0.0 -0.0292000000002 0 2.0 1e-06 
0.0 -0.0291000000002 0 2.0 1e-06 
0.0 -0.0290000000002 0 2.0 1e-06 
0.0 -0.0289000000002 0 2.0 1e-06 
0.0 -0.0288000000002 0 2.0 1e-06 
0.0 -0.0287000000002 0 2.0 1e-06 
0.0 -0.0286000000002 0 2.0 1e-06 
0.0 -0.0285000000002 0 2.0 1e-06 
0.0 -0.0284000000002 0 2.0 1e-06 
0.0 -0.0283000000002 0 2.0 1e-06 
0.0 -0.0282000000002 0 2.0 1e-06 
0.0 -0.0281000000002 0 2.0 1e-06 
0.0 -0.0280000000002 0 2.0 1e-06 
0.0 -0.0279000000002 0 2.0 1e-06 
0.0 -0.0278000000002 0 2.0 1e-06 
0.0 -0.0277000000002 0 2.0 1e-06 
0.0 -0.0276000000002 0 2.0 1e-06 
0.0 -0.0275000000002 0 2.0 1e-06 
0.0 -0.0274000000002 0 2.0 1e-06 
0.0 -0.0273000000002 0 2.0 1e-06 
0.0 -0.0272000000002 0 2.0 1e-06 
0.0 -0.0271000000002 0 2.0 1e-06 
0.0 -0.0270000000002 0 2.0 1e-06 
0.0 -0.0269000000002 0 2.0 1e-06 
0.0 -0.0268000000002 0 2.0 1e-06 
0.0 -0.0267000000002 0 2.0 1e-06 
0.0 -0.0266000000002 0 2.0 1e-06 
0.0 -0.0265000000002 0 2.0 1e-06 
0.0 -0.0264000000002 0 2.0 1e-06 
0.0 -0.0263000000002 0 2.0 1e-06 
0.0 -0.0262000000002 0 2.0 1e-06 
0.0 -0.0261000000002 0 2.0 1e-06 
0.0 -0.0260000000002 0 2.0 1e-06 
0.0 -0.0259000000002 0 2.0 1e-06 
0.0 -0.0258000000002 0 2.0 1e-06 
0.0 -0.0257000000002 0 2.0 1e-06 
0.0 -0.0256000000002 0 2.0 1e-06 
0.0 -0.0255000000002 0 2.0 1e-06 
0.0 -0.0254000000002 0 2.0 1e-06 
0.0 -0.0253000000002 0 2.0 1e-06 
0.0 -0.0252000000002 0 2.0 1e-06 
0.0 -0.0251000000002 0 2.0 1e-06 
0.0 -0.0250000000002 0 2.0 1e-06 
0.0 -0.0249000000002 0 2.0 1e-06 
0.0 -0.0248000000002 0 2.0 1e-06 
0.0 -0.0247000000002 0 2.0 1e-06 
0.0 -0.0246000000002 0 2.0 1e-06 
0.0 -0.0245000000002 0 2.0 1e-06 
0.0 -0.0244000000002 0 2.0 1e-06 
0.0 -0.0243000000002 0 2.0 1e-06 
0.0 -0.0242000000002 0 2.0 1e-06 
0.0 -0.0241000000002 0 2.0 1e-06 
0.0 -0.0240000000002 0 2.0 1e-06 
0.0 -0.0239000000002 0 2.0 1e-06 
0.0 -0.0238000000002 0 2.0 1e-06 
0.0 -0.0237000000002 0 2.0 1e-06 
0.0 -0.0236000000002 0 2.0 1e-06 
0.0 -0.0235000000002 0 2.0 1e-06 
0.0 -0.0234000000002 0 2.0 1e-06 
0.0 -0.0233000000002 0 2.0 1e-06 
0.0 -0.0232000000002 0 2.0 1e-06 
0.0 -0.0231000000002 0 2.0 1e-06 
0.0 -0.0230000000002 0 2.0 1e-06 
0.0 -0.0229000000002 0 2.0 1e-06 
0.0 -0.0228000000002 0 2.0 1e-06 
0.0 -0.0227000000002 0 2.0 1e-06 
0.0 -0.0226000000002 0 2.0 1e-06 
0.0 -0.0225000000002 0 2.0 1e-06 
0.0 -0.0224000000002 0 2.0 1e-06 
0.0 -0.0223000000002 0 2.0 1e-06 
0.0 -0.0222000000002 0 2.0 1e-06 
0.0 -0.0221000000002 0 2.0 1e-06 
0.0 -0.0220000000002 0 2.0 1e-06 
0.0 -0.0219000000002 0 2.0 1e-06 
0.0 -0.0218000000002 0 2.0 1e-06 
0.0 -0.0217000000002 0 2.0 1e-06 
0.0 -0.0216000000002 0 2.0 1e-06 
0.0 -0.0215000000002 0 2.0 1e-06 
0.0 -0.0214000000002 0 2.0 1e-06 
0.0 -0.0213000000002 0 2.0 1e-06 
0.0 -0.0212000000002 0 2.0 1e-06 
0.0 -0.0211000000002 0 2.0 1e-06 
0.0 -0.0210000000002 0 2.0 1e-06 
0.0 -0.0209000000002 0 2.0 1e-06 
0.0 -0.0208000000002 0 2.0 1e-06 
0.0 -0.0207000000002 0 2.0 1e-06 
0.0 -0.0206000000002 0 2.0 1e-06 
0.0 -0.0205000000002 0 2.0 1e-06 
0.0 -0.0204000000002 0 2.0 1e-06 
0.0 -0.0203000000002 0 2.0 1e-06 
0.0 -0.0202000000002 0 2.0 1e-06 
0.0 -0.0201000000002 0 2.0 1e-06 
0.0 -0.0200000000002 0 2.0 1e-06 
0.0 -0.0199000000002 0 2.0 1e-06 
0.0 -0.0198000000002 0 2.0 1e-06 
0.0 -0.0197000000002 0 2.0 1e-06 
0.0 -0.0196000000002 0 2.0 1e-06 
0.0 -0.0195000000002 0 2.0 1e-06 
0.0 -0.0194000000002 0 2.0 1e-06 
0.0 -0.0193000000002 0 2.0 1e-06 
0.0 -0.0192000000002 0 2.0 1e-06 
0.0 -0.0191000000002 0 2.0 1e-06 
0.0 -0.0190000000002 0 2.0 1e-06 
0.0 -0.0189000000002 0 2.0 1e-06 
0.0 -0.0188000000002 0 2.0 1e-06 
0.0 -0.0187000000002 0 2.0 1e-06 
0.0 -0.0186000000002 0 2.0 1e-06 
0.0 -0.0185000000002 0 2.0 1e-06 
0.0 -0.0184000000002 0 2.0 1e-06 
0.0 -0.0183000000002 0 2.0 1e-06 
0.0 -0.0182000000002 0 2.0 1e-06 
0.0 -0.0181000000002 0 2.0 1e-06 
0.0 -0.0180000000002 0 2.0 1e-06 
0.0 -0.0179000000002 0 2.0 1e-06 
0.0 -0.0178000000002 0 2.0 1e-06 
0.0 -0.0177000000002 0 2.0 1e-06 
0.0 -0.0176000000002 0 2.0 1e-06 
0.0 -0.0175000000002 0 2.0 1e-06 
0.0 -0.0174000000002 0 2.0 1e-06 
0.0 -0.0173000000002 0 2.0 1e-06 
0.0 -0.0172000000002 0 2.0 1e-06 
0.0 -0.0171000000002 0 2.0 1e-06 
0.0 -0.0170000000002 0 2.0 1e-06 
0.0 -0.0169000000002 0 2.0 1e-06 
0.0 -0.0168000000002 0 2.0 1e-06 
0.0 -0.0167000000002 0 2.0 1e-06 
0.0 -0.0166000000002 0 2.0 1e-06 
0.0 -0.0165000000002 0 2.0 1e-06 
0.0 -0.0164000000002 0 2.0 1e-06 
0.0 -0.0163000000002 0 2.0 1e-06 
0.0 -0.0162000000002 0 2.0 1e-06 
0.0 -0.0161000000002 0 2.0 1e-06 
0.0 -0.0160000000002 0 2.0 1e-06 
0.0 -0.0159000000002 0 2.0 1e-06 
0.0 -0.0158000000002 0 2.0 1e-06 
0.0 -0.0157000000002 0 2.0 1e-06 
0.0 -0.0156000000002 0 2.0 1e-06 
0.0 -0.0155000000002 0 2.0 1e-06 
0.0 -0.0154000000002 0 2.0 1e-06 
0.0 -0.0153000000002 0 2.0 1e-06 
0.0 -0.0152000000002 0 2.0 1e-06 
0.0 -0.0151000000002 0 2.0 1e-06 
0.0 -0.0150000000002 0 2.0 1e-06 
0.0 -0.0149000000002 0 2.0 1e-06 
0.0 -0.0148000000002 0 2.0 1e-06 
0.0 -0.0147000000002 0 2.0 1e-06 
0.0 -0.0146000000002 0 2.0 1e-06 
0.0 -0.0145000000002 0 2.0 1e-06 
0.0 -0.0144000000002 0 2.0 1e-06 
0.0 -0.0143000000002 0 2.0 1e-06 
0.0 -0.0142000000002 0 2.0 1e-06 
0.0 -0.0141000000002 0 2.0 1e-06 
0.0 -0.0140000000002 0 2.0 1e-06 
0.0 -0.0139000000002 0 2.0 1e-06 
0.0 -0.0138000000002 0 2.0 1e-06 
0.0 -0.0137000000002 0 2.0 1e-06 
0.0 -0.0136000000002 0 2.0 1e-06 
0.0 -0.0135000000002 0 2.0 1e-06 
0.0 -0.0134000000002 0 2.0 1e-06 
0.0 -0.0133000000002 0 2.0 1e-06 
0.0 -0.0132000000002 0 2.0 1e-06 
0.0 -0.0131000000002 0 2.0 1e-06 
0.0 -0.0130000000002 0 2.0 1e-06 
0.0 -0.0129000000002 0 2.0 1e-06 
0.0 -0.0128000000002 0 2.0 1e-06 
0.0 -0.0127000000002 0 2.0 1e-06 
0.0 -0.0126000000002 0 2.0 1e-06 
0.0 -0.0125000000002 0 2.0 1e-06 
0.0 -0.0124000000002 0 2.0 1e-06 
0.0 -0.0123000000002 0 2.0 1e-06 
0.0 -0.0122000000002 0 2.0 1e-06 
0.0 -0.0121000000002 0 2.0 1e-06 
0.0 -0.0120000000002 0 2.0 1e-06 
0.0 -0.0119000000002 0 2.0 1e-06 
0.0 -0.0118000000002 0 2.0 1e-06 
0.0 -0.0117000000002 0 2.0 1e-06 
0.0 -0.0116000000002 0 2.0 1e-06 
0.0 -0.0115000000002 0 2.0 1e-06 
0.0 -0.0114000000002 0 2.0 1e-06 
0.0 -0.0113000000002 0 2.0 1e-06 
0.0 -0.0112000000002 0 2.0 1e-06 
0.0 -0.0111000000002 0 2.0 1e-06 
0.0 -0.0110000000002 0 2.0 1e-06 
0.0 -0.0109000000002 0 2.0 1e-06 
0.0 -0.0108000000002 0 2.0 1e-06 
0.0 -0.0107000000002 0 2.0 1e-06 
0.0 -0.0106000000002 0 2.0 1e-06 
0.0 -0.0105000000002 0 2.0 1e-06 
0.0 -0.0104000000002 0 2.0 1e-06 
0.0 -0.0103000000002 0 2.0 1e-06 
0.0 -0.0102000000002 0 2.0 1e-06 
0.0 -0.0101000000002 0 2.0 1e-06 
0.0 -0.0100000000002 0 2.0 1e-06 
0.0 -0.00990000000016 0 2.0 1e-06 
0.0 -0.00980000000016 0 2.0 1e-06 
0.0 -0.00970000000016 0 2.0 1e-06 
0.0 -0.00960000000016 0 2.0 1e-06 
0.0 -0.00950000000016 0 2.0 1e-06 
0.0 -0.00940000000016 0 2.0 1e-06 
0.0 -0.00930000000016 0 2.0 1e-06 
0.0 -0.00920000000016 0 2.0 1e-06 
0.0 -0.00910000000016 0 2.0 1e-06 
0.0 -0.00900000000016 0 2.0 1e-06 
0.0 -0.00890000000016 0 2.0 1e-06 
0.0 -0.00880000000016 0 2.0 1e-06 
0.0 -0.00870000000016 0 2.0 1e-06 
0.0 -0.00860000000016 0 2.0 1e-06 
0.0 -0.00850000000016 0 2.0 1e-06 
0.0 -0.00840000000016 0 2.0 1e-06 
0.0 -0.00830000000016 0 2.0 1e-06 
0.0 -0.00820000000016 0 2.0 1e-06 
0.0 -0.00810000000016 0 2.0 1e-06 
0.0 -0.00800000000016 0 2.0 1e-06 
0.0 -0.00790000000016 0 2.0 1e-06 
0.0 -0.00780000000016 0 2.0 1e-06 
0.0 -0.00770000000016 0 2.0 1e-06 
0.0 -0.00760000000016 0 2.0 1e-06 
0.0 -0.00750000000016 0 2.0 1e-06 
0.0 -0.00740000000016 0 2.0 1e-06 
0.0 -0.00730000000016 0 2.0 1e-06 
0.0 -0.00720000000016 0 2.0 1e-06 
0.0 -0.00710000000016 0 2.0 1e-06 
0.0 -0.00700000000016 0 2.0 1e-06 
0.0 -0.00690000000016 0 2.0 1e-06 
0.0 -0.00680000000016 0 2.0 1e-06 
0.0 -0.00670000000016 0 2.0 1e-06 
0.0 -0.00660000000016 0 2.0 1e-06 
0.0 -0.00650000000016 0 2.0 1e-06 
0.0 -0.00640000000016 0 2.0 1e-06 
0.0 -0.00630000000016 0 2.0 1e-06 
0.0 -0.00620000000016 0 2.0 1e-06 
0.0 -0.00610000000016 0 2.0 1e-06 
0.0 -0.00600000000016 0 2.0 1e-06 
0.0 -0.00590000000016 0 2.0 1e-06 
0.0 -0.00580000000016 0 2.0 1e-06 
0.0 -0.00570000000016 0 2.0 1e-06 
0.0 -0.00560000000016 0 2.0 1e-06 
0.0 -0.00550000000016 0 2.0 1e-06 
0.0 -0.00540000000016 0 2.0 1e-06 
0.0 -0.00530000000016 0 2.0 1e-06 
0.0 -0.00520000000016 0 2.0 1e-06 
0.0 -0.00510000000016 0 2.0 1e-06 
0.0 -0.00500000000016 0 2.0 1e-06 
0.0 -0.00490000000016 0 2.0 1e-06 
0.0 -0.00480000000016 0 2.0 1e-06 
0.0 -0.00470000000016 0 2.0 1e-06 
0.0 -0.00460000000016 0 2.0 1e-06 
0.0 -0.00450000000016 0 2.0 1e-06 
0.0 -0.00440000000016 0 2.0 1e-06 
0.0 -0.00430000000016 0 2.0 1e-06 
0.0 -0.00420000000016 0 2.0 1e-06 
0.0 -0.00410000000016 0 2.0 1e-06 
0.0 -0.00400000000016 0 2.0 1e-06 
0.0 -0.00390000000016 0 2.0 1e-06 
0.0 -0.00380000000016 0 2.0 1e-06 
0.0 -0.00370000000016 0 2.0 1e-06 
0.0 -0.00360000000016 0 2.0 1e-06 
0.0 -0.00350000000016 0 2.0 1e-06 
0.0 -0.00340000000016 0 2.0 1e-06 
0.0 -0.00330000000016 0 2.0 1e-06 
0.0 -0.00320000000016 0 2.0 1e-06 
0.0 -0.00310000000016 0 2.0 1e-06 
0.0 -0.00300000000016 0 2.0 1e-06 
0.0 -0.00290000000016 0 2.0 1e-06 
0.0 -0.00280000000016 0 2.0 1e-06 
0.0 -0.00270000000016 0 2.0 1e-06 
0.0 -0.00260000000016 0 2.0 1e-06 
0.0 -0.00250000000016 0 2.0 1e-06 
0.0 -0.00240000000016 0 2.0 1e-06 
0.0 -0.00230000000016 0 2.0 1e-06 
0.0 -0.00220000000016 0 2.0 1e-06 
0.0 -0.00210000000016 0 2.0 1e-06 
0.0 -0.00200000000016 0 2.0 1e-06 
0.0 -0.00190000000016 0 2.0 1e-06 
0.0 -0.00180000000017 0 2.0 1e-06 
0.0 -0.00170000000017 0 2.0 1e-06 
0.0 -0.00160000000017 0 2.0 1e-06 
0.0 -0.00150000000017 0 2.0 1e-06 
0.0 -0.00140000000017 0 2.0 1e-06 
0.0 -0.00130000000017 0 2.0 1e-06 
0.0 -0.00120000000017 0 2.0 1e-06 
0.0 -0.00110000000017 0 2.0 1e-06 
0.0 -0.00100000000017 0 2.0 1e-06 
0.0 -0.000900000000165 0 2.0 1e-06 
0.0 -0.000800000000165 0 2.0 1e-06 
0.0 -0.000700000000165 0 2.0 1e-06 
0.0 -0.000600000000165 0 2.0 1e-06 
0.0 -0.000500000000165 0 2.0 1e-06 
0.0 -0.000400000000165 0 2.0 1e-06 
0.0 -0.000300000000165 0 2.0 1e-06 
0.0 -0.000200000000165 0 2.0 1e-06 
0.0 -0.000100000000165 0 2.0 1e-06 
0.0 -1.65201186064e-13 0 2.0 1e-06 
0.0 9.99999998348e-05 0 2.0 1e-06 
0.0 0.000199999999835 0 2.0 1e-06 
0.0 0.000299999999835 0 2.0 1e-06 
0.0 0.000399999999835 0 2.0 1e-06 
0.0 0.000499999999835 0 2.0 1e-06 
0.0 0.000599999999835 0 2.0 1e-06 
0.0 0.000699999999835 0 2.0 1e-06 
0.0 0.000799999999835 0 2.0 1e-06 
0.0 0.000899999999835 0 2.0 1e-06 
0.0 0.000999999999835 0 2.0 1e-06 
0.0 0.00109999999983 0 2.0 1e-06 
0.0 0.00119999999983 0 2.0 1e-06 
0.0 0.00129999999983 0 2.0 1e-06 
0.0 0.00139999999983 0 2.0 1e-06 
0.0 0.00149999999983 0 2.0 1e-06 
0.0 0.00159999999983 0 2.0 1e-06 
0.0 0.00169999999983 0 2.0 1e-06 
0.0 0.00179999999983 0 2.0 1e-06 
0.0 0.00189999999983 0 2.0 1e-06 
0.0 0.00199999999983 0 2.0 1e-06 
0.0 0.00209999999983 0 2.0 1e-06 
0.0 0.00219999999983 0 2.0 1e-06 
0.0 0.00229999999983 0 2.0 1e-06 
0.0 0.00239999999983 0 2.0 1e-06 
0.0 0.00249999999983 0 2.0 1e-06 
0.0 0.00259999999983 0 2.0 1e-06 
0.0 0.00269999999983 0 2.0 1e-06 
0.0 0.00279999999983 0 2.0 1e-06 
0.0 0.00289999999983 0 2.0 1e-06 
0.0 0.00299999999983 0 2.0 1e-06 
0.0 0.00309999999983 0 2.0 1e-06 
0.0 0.00319999999983 0 2.0 1e-06 
0.0 0.00329999999983 0 2.0 1e-06 
0.0 0.00339999999983 0 2.0 1e-06 
0.0 0.00349999999983 0 2.0 1e-06 
0.0 0.00359999999983 0 2.0 1e-06 
0.0 0.00369999999983 0 2.0 1e-06 
0.0 0.00379999999983 0 2.0 1e-06 
0.0 0.00389999999983 0 2.0 1e-06 
0.0 0.00399999999983 0 2.0 1e-06 
0.0 0.00409999999983 0 2.0 1e-06 
0.0 0.00419999999983 0 2.0 1e-06 
0.0 0.00429999999983 0 2.0 1e-06 
0.0 0.00439999999983 0 2.0 1e-06 
0.0 0.00449999999983 0 2.0 1e-06 
0.0 0.00459999999983 0 2.0 1e-06 
0.0 0.00469999999983 0 2.0 1e-06 
0.0 0.00479999999983 0 2.0 1e-06 
0.0 0.00489999999983 0 2.0 1e-06 
0.0 0.00499999999983 0 2.0 1e-06 
0.0 0.00509999999983 0 2.0 1e-06 
0.0 0.00519999999983 0 2.0 1e-06 
0.0 0.00529999999983 0 2.0 1e-06 
0.0 0.00539999999983 0 2.0 1e-06 
0.0 0.00549999999983 0 2.0 1e-06 
0.0 0.00559999999983 0 2.0 1e-06 
0.0 0.00569999999983 0 2.0 1e-06 
0.0 0.00579999999983 0 2.0 1e-06 
0.0 0.00589999999983 0 2.0 1e-06 
0.0 0.00599999999983 0 2.0 1e-06 
0.0 0.00609999999983 0 2.0 1e-06 
0.0 0.00619999999983 0 2.0 1e-06 
0.0 0.00629999999983 0 2.0 1e-06 
0.0 0.00639999999983 0 2.0 1e-06 
0.0 0.00649999999983 0 2.0 1e-06 
0.0 0.00659999999983 0 2.0 1e-06 
0.0 0.00669999999983 0 2.0 1e-06 
0.0 0.00679999999983 0 2.0 1e-06 
0.0 0.00689999999983 0 2.0 1e-06 
0.0 0.00699999999983 0 2.0 1e-06 
0.0 0.00709999999983 0 2.0 1e-06 
0.0 0.00719999999983 0 2.0 1e-06 
0.0 0.00729999999983 0 2.0 1e-06 
0.0 0.00739999999983 0 2.0 1e-06 
0.0 0.00749999999983 0 2.0 1e-06 
0.0 0.00759999999983 0 2.0 1e-06 
0.0 0.00769999999983 0 2.0 1e-06 
0.0 0.00779999999983 0 2.0 1e-06 
0.0 0.00789999999983 0 2.0 1e-06 
0.0 0.00799999999983 0 2.0 1e-06 
0.0 0.00809999999983 0 2.0 1e-06 
0.0 0.00819999999983 0 2.0 1e-06 
0.0 0.00829999999983 0 2.0 1e-06 
0.0 0.00839999999983 0 2.0 1e-06 
0.0 0.00849999999983 0 2.0 1e-06 
0.0 0.00859999999983 0 2.0 1e-06 
0.0 0.00869999999983 0 2.0 1e-06 
0.0 0.00879999999983 0 2.0 1e-06 
0.0 0.00889999999983 0 2.0 1e-06 
0.0 0.00899999999983 0 2.0 1e-06 
0.0 0.00909999999983 0 2.0 1e-06 
0.0 0.00919999999983 0 2.0 1e-06 
0.0 0.00929999999983 0 2.0 1e-06 
0.0 0.00939999999983 0 2.0 1e-06 
0.0 0.00949999999983 0 2.0 1e-06 
0.0 0.00959999999983 0 2.0 1e-06 
0.0 0.00969999999983 0 2.0 1e-06 
0.0 0.00979999999983 0 2.0 1e-06 
0.0 0.00989999999983 0 2.0 1e-06 
0.0 0.00999999999983 0 2.0 1e-06 
0.0 0.0100999999998 0 2.0 1e-06 
0.0 0.0101999999998 0 2.0 1e-06 
0.0 0.0102999999998 0 2.0 1e-06 
0.0 0.0103999999998 0 2.0 1e-06 
0.0 0.0104999999998 0 2.0 1e-06 
0.0 0.0105999999998 0 2.0 1e-06 
0.0 0.0106999999998 0 2.0 1e-06 
0.0 0.0107999999998 0 2.0 1e-06 
0.0 0.0108999999998 0 2.0 1e-06 
0.0 0.0109999999998 0 2.0 1e-06 
0.0 0.0110999999998 0 2.0 1e-06 
0.0 0.0111999999998 0 2.0 1e-06 
0.0 0.0112999999998 0 2.0 1e-06 
0.0 0.0113999999998 0 2.0 1e-06 
0.0 0.0114999999998 0 2.0 1e-06 
0.0 0.0115999999998 0 2.0 1e-06 
0.0 0.0116999999998 0 2.0 1e-06 
0.0 0.0117999999998 0 2.0 1e-06 
0.0 0.0118999999998 0 2.0 1e-06 
0.0 0.0119999999998 0 2.0 1e-06 
0.0 0.0120999999998 0 2.0 1e-06 
0.0 0.0121999999998 0 2.0 1e-06 
0.0 0.0122999999998 0 2.0 1e-06 
0.0 0.0123999999998 0 2.0 1e-06 
0.0 0.0124999999998 0 2.0 1e-06 
0.0 0.0125999999998 0 2.0 1e-06 
0.0 0.0126999999998 0 2.0 1e-06 
0.0 0.0127999999998 0 2.0 1e-06 
0.0 0.0128999999998 0 2.0 1e-06 
0.0 0.0129999999998 0 2.0 1e-06 
0.0 0.0130999999998 0 2.0 1e-06 
0.0 0.0131999999998 0 2.0 1e-06 
0.0 0.0132999999998 0 2.0 1e-06 
0.0 0.0133999999998 0 2.0 1e-06 
0.0 0.0134999999998 0 2.0 1e-06 
0.0 0.0135999999998 0 2.0 1e-06 
0.0 0.0136999999998 0 2.0 1e-06 
0.0 0.0137999999998 0 2.0 1e-06 
0.0 0.0138999999998 0 2.0 1e-06 
0.0 0.0139999999998 0 2.0 1e-06 
0.0 0.0140999999998 0 2.0 1e-06 
0.0 0.0141999999998 0 2.0 1e-06 
0.0 0.0142999999998 0 2.0 1e-06 
0.0 0.0143999999998 0 2.0 1e-06 
0.0 0.0144999999998 0 2.0 1e-06 
0.0 0.0145999999998 0 2.0 1e-06 
0.0 0.0146999999998 0 2.0 1e-06 
0.0 0.0147999999998 0 2.0 1e-06 
0.0 0.0148999999998 0 2.0 1e-06 
0.0 0.0149999999998 0 2.0 1e-06 
0.0 0.0150999999998 0 2.0 1e-06 
0.0 0.0151999999998 0 2.0 1e-06 
0.0 0.0152999999998 0 2.0 1e-06 
0.0 0.0153999999998 0 2.0 1e-06 
0.0 0.0154999999998 0 2.0 1e-06 
0.0 0.0155999999998 0 2.0 1e-06 
0.0 0.0156999999998 0 2.0 1e-06 
0.0 0.0157999999998 0 2.0 1e-06 
0.0 0.0158999999998 0 2.0 1e-06 
0.0 0.0159999999998 0 2.0 1e-06 
0.0 0.0160999999998 0 2.0 1e-06 
0.0 0.0161999999998 0 2.0 1e-06 
0.0 0.0162999999998 0 2.0 1e-06 
0.0 0.0163999999998 0 2.0 1e-06 
0.0 0.0164999999998 0 2.0 1e-06 
0.0 0.0165999999998 0 2.0 1e-06 
0.0 0.0166999999998 0 2.0 1e-06 
0.0 0.0167999999998 0 2.0 1e-06 
0.0 0.0168999999998 0 2.0 1e-06 
0.0 0.0169999999998 0 2.0 1e-06 
0.0 0.0170999999998 0 2.0 1e-06 
0.0 0.0171999999998 0 2.0 1e-06 
0.0 0.0172999999998 0 2.0 1e-06 
0.0 0.0173999999998 0 2.0 1e-06 
0.0 0.0174999999998 0 2.0 1e-06 
0.0 0.0175999999998 0 2.0 1e-06 
0.0 0.0176999999998 0 2.0 1e-06 
0.0 0.0177999999998 0 2.0 1e-06 
0.0 0.0178999999998 0 2.0 1e-06 
0.0 0.0179999999998 0 2.0 1e-06 
0.0 0.0180999999998 0 2.0 1e-06 
0.0 0.0181999999998 0 2.0 1e-06 
0.0 0.0182999999998 0 2.0 1e-06 
0.0 0.0183999999998 0 2.0 1e-06 
0.0 0.0184999999998 0 2.0 1e-06 
0.0 0.0185999999998 0 2.0 1e-06 
0.0 0.0186999999998 0 2.0 1e-06 
0.0 0.0187999999998 0 2.0 1e-06 
0.0 0.0188999999998 0 2.0 1e-06 
0.0 0.0189999999998 0 2.0 1e-06 
0.0 0.0190999999998 0 2.0 1e-06 
0.0 0.0191999999998 0 2.0 1e-06 
0.0 0.0192999999998 0 2.0 1e-06 
0.0 0.0193999999998 0 2.0 1e-06 
0.0 0.0194999999998 0 2.0 1e-06 
0.0 0.0195999999998 0 2.0 1e-06 
0.0 0.0196999999998 0 2.0 1e-06 
0.0 0.0197999999998 0 2.0 1e-06 
0.0 0.0198999999998 0 2.0 1e-06 
0.0 0.0199999999998 0 2.0 1e-06 
0.0 0.0200999999998 0 2.0 1e-06 
0.0 0.0201999999998 0 2.0 1e-06 
0.0 0.0202999999998 0 2.0 1e-06 
0.0 0.0203999999998 0 2.0 1e-06 
0.0 0.0204999999998 0 2.0 1e-06 
0.0 0.0205999999998 0 2.0 1e-06 
0.0 0.0206999999998 0 2.0 1e-06 
0.0 0.0207999999998 0 2.0 1e-06 
0.0 0.0208999999998 0 2.0 1e-06 
0.0 0.0209999999998 0 2.0 1e-06 
0.0 0.0210999999998 0 2.0 1e-06 
0.0 0.0211999999998 0 2.0 1e-06 
0.0 0.0212999999998 0 2.0 1e-06 
0.0 0.0213999999998 0 2.0 1e-06 
0.0 0.0214999999998 0 2.0 1e-06 
0.0 0.0215999999998 0 2.0 1e-06 
0.0 0.0216999999998 0 2.0 1e-06 
0.0 0.0217999999998 0 2.0 1e-06 
0.0 0.0218999999998 0 2.0 1e-06 
0.0 0.0219999999998 0 2.0 1e-06 
0.0 0.0220999999998 0 2.0 1e-06 
0.0 0.0221999999998 0 2.0 1e-06 
0.0 0.0222999999998 0 2.0 1e-06 
0.0 0.0223999999998 0 2.0 1e-06 
0.0 0.0224999999998 0 2.0 1e-06 
0.0 0.0225999999998 0 2.0 1e-06 
0.0 0.0226999999998 0 2.0 1e-06 
0.0 0.0227999999998 0 2.0 1e-06 
0.0 0.0228999999998 0 2.0 1e-06 
0.0 0.0229999999998 0 2.0 1e-06 
0.0 0.0230999999998 0 2.0 1e-06 
0.0 0.0231999999998 0 2.0 1e-06 
0.0 0.0232999999998 0 2.0 1e-06 
0.0 0.0233999999998 0 2.0 1e-06 
0.0 0.0234999999998 0 2.0 1e-06 
0.0 0.0235999999998 0 2.0 1e-06 
0.0 0.0236999999998 0 2.0 1e-06 
0.0 0.0237999999998 0 2.0 1e-06 
0.0 0.0238999999998 0 2.0 1e-06 
0.0 0.0239999999998 0 2.0 1e-06 
0.0 0.0240999999998 0 2.0 1e-06 
0.0 0.0241999999998 0 2.0 1e-06 
0.0 0.0242999999998 0 2.0 1e-06 
0.0 0.0243999999998 0 2.0 1e-06 
0.0 0.0244999999998 0 2.0 1e-06 
0.0 0.0245999999998 0 2.0 1e-06 
0.0 0.0246999999998 0 2.0 1e-06 
0.0 0.0247999999998 0 2.0 1e-06 
0.0 0.0248999999998 0 2.0 1e-06 
0.0 0.0249999999998 0 2.0 1e-06 
0.0 0.0250999999998 0 2.0 1e-06 
0.0 0.0251999999998 0 2.0 1e-06 
0.0 0.0252999999998 0 2.0 1e-06 
0.0 0.0253999999998 0 2.0 1e-06 
0.0 0.0254999999998 0 2.0 1e-06 
0.0 0.0255999999998 0 2.0 1e-06 
0.0 0.0256999999998 0 2.0 1e-06 
0.0 0.0257999999998 0 2.0 1e-06 
0.0 0.0258999999998 0 2.0 1e-06 
0.0 0.0259999999998 0 2.0 1e-06 
0.0 0.0260999999998 0 2.0 1e-06 
0.0 0.0261999999998 0 2.0 1e-06 
0.0 0.0262999999998 0 2.0 1e-06 
0.0 0.0263999999998 0 2.0 1e-06 
0.0 0.0264999999998 0 2.0 1e-06 
0.0 0.0265999999998 0 2.0 1e-06 
0.0 0.0266999999998 0 2.0 1e-06 
0.0 0.0267999999998 0 2.0 1e-06 
0.0 0.0268999999998 0 2.0 1e-06 
0.0 0.0269999999998 0 2.0 1e-06 
0.0 0.0270999999998 0 2.0 1e-06 
0.0 0.0271999999998 0 2.0 1e-06 
0.0 0.0272999999998 0 2.0 1e-06 
0.0 0.0273999999998 0 2.0 1e-06 
0.0 0.0274999999998 0 2.0 1e-06 
0.0 0.0275999999998 0 2.0 1e-06 
0.0 0.0276999999998 0 2.0 1e-06 
0.0 0.0277999999998 0 2.0 1e-06 
0.0 0.0278999999998 0 2.0 1e-06 
0.0 0.0279999999998 0 2.0 1e-06 
0.0 0.0280999999998 0 2.0 1e-06 
0.0 0.0281999999998 0 2.0 1e-06 
0.0 0.0282999999998 0 2.0 1e-06 
0.0 0.0283999999998 0 2.0 1e-06 
0.0 0.0284999999998 0 2.0 1e-06 
0.0 0.0285999999998 0 2.0 1e-06 
0.0 0.0286999999998 0 2.0 1e-06 
0.0 0.0287999999998 0 2.0 1e-06 
0.0 0.0288999999998 0 2.0 1e-06 
0.0 0.0289999999998 0 2.0 1e-06 
0.0 0.0290999999998 0 2.0 1e-06 
0.0 0.0291999999998 0 2.0 1e-06 
0.0 0.0292999999998 0 2.0 1e-06 
0.0 0.0293999999998 0 2.0 1e-06 
0.0 0.0294999999998 0 2.0 1e-06 
0.0 0.0295999999998 0 2.0 1e-06 
0.0 0.0296999999998 0 2.0 1e-06 
0.0 0.0297999999998 0 2.0 1e-06 
0.0 0.0298999999998 0 2.0 1e-06 
0.0 0.0299999999998 0 2.0 1e-06 
0.0 0.0300999999998 0 2.0 1e-06 
0.0 0.0301999999998 0 2.0 1e-06 
0.0 0.0302999999998 0 2.0 1e-06 
0.0 0.0303999999998 0 2.0 1e-06 
0.0 0.0304999999998 0 2.0 1e-06 
0.0 0.0305999999998 0 2.0 1e-06 
0.0 0.0306999999998 0 2.0 1e-06 
0.0 0.0307999999998 0 2.0 1e-06 
0.0 0.0308999999998 0 2.0 1e-06 
0.0 0.0309999999998 0 2.0 1e-06 
0.0 0.0310999999998 0 2.0 1e-06 
0.0 0.0311999999998 0 2.0 1e-06 
0.0 0.0312999999998 0 2.0 1e-06 
0.0 0.0313999999998 0 2.0 1e-06 
0.0 0.0314999999998 0 2.0 1e-06 
0.0 0.0315999999998 0 2.0 1e-06 
0.0 0.0316999999998 0 2.0 1e-06 
0.0 0.0317999999998 0 2.0 1e-06 
0.0 0.0318999999998 0 2.0 1e-06 
0.0 0.0319999999998 0 2.0 1e-06 
0.0 0.0320999999998 0 2.0 1e-06 
0.0 0.0321999999998 0 2.0 1e-06 
0.0 0.0322999999998 0 2.0 1e-06 
0.0 0.0323999999998 0 2.0 1e-06 
0.0 0.0324999999998 0 2.0 1e-06 
0.0 0.0325999999998 0 2.0 1e-06 
0.0 0.0326999999998 0 2.0 1e-06 
0.0 0.0327999999998 0 2.0 1e-06 
0.0 0.0328999999998 0 2.0 1e-06 
0.0 0.0329999999998 0 2.0 1e-06 
0.0 0.0330999999998 0 2.0 1e-06 
0.0 0.0331999999998 0 2.0 1e-06 
0.0 0.0332999999998 0 2.0 1e-06 
0.0 0.0333999999998 0 2.0 1e-06 
0.0 0.0334999999998 0 2.0 1e-06 
0.0 0.0335999999998 0 2.0 1e-06 
0.0 0.0336999999998 0 2.0 1e-06 
0.0 0.0337999999998 0 2.0 1e-06 
0.0 0.0338999999998 0 2.0 1e-06 
0.0 0.0339999999998 0 2.0 1e-06 
0.0 0.0340999999998 0 2.0 1e-06 
0.0 0.0341999999998 0 2.0 1e-06 
0.0 0.0342999999998 0 2.0 1e-06 
0.0 0.0343999999998 0 2.0 1e-06 
0.0 0.0344999999998 0 2.0 1e-06 
0.0 0.0345999999998 0 2.0 1e-06 
0.0 0.0346999999998 0 2.0 1e-06 
0.0 0.0347999999998 0 2.0 1e-06 
0.0 0.0348999999998 0 2.0 1e-06 
0.0 0.0349999999998 0 2.0 1e-06 
0.0 0.0350999999998 0 2.0 1e-06 
0.0 0.0351999999998 0 2.0 1e-06 
0.0 0.0352999999998 0 2.0 1e-06 
0.0 0.0353999999998 0 2.0 1e-06 
0.0 0.0354999999998 0 2.0 1e-06 
0.0 0.0355999999998 0 2.0 1e-06 
0.0 0.0356999999998 0 2.0 1e-06 
0.0 0.0357999999998 0 2.0 1e-06 
0.0 0.0358999999998 0 2.0 1e-06 
0.0 0.0359999999998 0 2.0 1e-06 
0.0 0.0360999999998 0 2.0 1e-06 
0.0 0.0361999999998 0 2.0 1e-06 
0.0 0.0362999999998 0 2.0 1e-06 
0.0 0.0363999999998 0 2.0 1e-06 
0.0 0.0364999999998 0 2.0 1e-06 
0.0 0.0365999999998 0 2.0 1e-06 
0.0 0.0366999999998 0 2.0 1e-06 
0.0 0.0367999999998 0 2.0 1e-06 
0.0 0.0368999999998 0 2.0 1e-06 
0.0 0.0369999999998 0 2.0 1e-06 
0.0 0.0370999999998 0 2.0 1e-06 
0.0 0.0371999999998 0 2.0 1e-06 
0.0 0.0372999999998 0 2.0 1e-06 
0.0 0.0373999999998 0 2.0 1e-06 
0.0 0.0374999999998 0 2.0 1e-06 
0.0 0.0375999999998 0 2.0 1e-06 
0.0 0.0376999999998 0 2.0 1e-06 
0.0 0.0377999999998 0 2.0 1e-06 
0.0 0.0378999999998 0 2.0 1e-06 
0.0 0.0379999999998 0 2.0 1e-06 
0.0 0.0380999999998 0 2.0 1e-06 
0.0 0.0381999999998 0 2.0 1e-06 
0.0 0.0382999999998 0 2.0 1e-06 
0.0 0.0383999999998 0 2.0 1e-06 
0.0 0.0384999999998 0 2.0 1e-06 
0.0 0.0385999999998 0 2.0 1e-06 
0.0 0.0386999999998 0 2.0 1e-06 
0.0 0.0387999999998 0 2.0 1e-06 
0.0 0.0388999999998 0 2.0 1e-06 
0.0 0.0389999999998 0 2.0 1e-06 
0.0 0.0390999999998 0 2.0 1e-06 
0.0 0.0391999999998 0 2.0 1e-06 
0.0 0.0392999999998 0 2.0 1e-06 
0.0 0.0393999999998 0 2.0 1e-06 
0.0 0.0394999999998 0 2.0 1e-06 
0.0 0.0395999999998 0 2.0 1e-06 
0.0 0.0396999999998 0 2.0 1e-06 
0.0 0.0397999999998 0 2.0 1e-06 
0.0 0.0398999999998 0 2.0 1e-06 
0.0 0.0399999999998 0 2.0 1e-06 
0.0 0.0400999999998 0 2.0 1e-06 
0.0 0.0401999999998 0 2.0 1e-06 
0.0 0.0402999999998 0 2.0 1e-06 
0.0 0.0403999999998 0 2.0 1e-06 
0.0 0.0404999999998 0 2.0 1e-06 
0.0 0.0405999999998 0 2.0 1e-06 
0.0 0.0406999999998 0 2.0 1e-06 
0.0 0.0407999999998 0 2.0 1e-06 
0.0 0.0408999999998 0 2.0 1e-06 
0.0 0.0409999999998 0 2.0 1e-06 
0.0 0.0410999999998 0 2.0 1e-06 
0.0 0.0411999999998 0 2.0 1e-06 
0.0 0.0412999999998 0 2.0 1e-06 
0.0 0.0413999999998 0 2.0 1e-06 
0.0 0.0414999999998 0 2.0 1e-06 
0.0 0.0415999999998 0 2.0 1e-06 
0.0 0.0416999999998 0 2.0 1e-06 
0.0 0.0417999999998 0 2.0 1e-06 
0.0 0.0418999999998 0 2.0 1e-06 
0.0 0.0419999999998 0 2.0 1e-06 
0.0 0.0420999999998 0 2.0 1e-06 
0.0 0.0421999999998 0 2.0 1e-06 
0.0 0.0422999999998 0 2.0 1e-06 
0.0 0.0423999999998 0 2.0 1e-06 
0.0 0.0424999999998 0 2.0 1e-06 
0.0 0.0425999999998 0 2.0 1e-06 
0.0 0.0426999999998 0 2.0 1e-06 
0.0 0.0427999999998 0 2.0 1e-06 
0.0 0.0428999999998 0 2.0 1e-06 
0.0 0.0429999999998 0 2.0 1e-06 
0.0 0.0430999999998 0 2.0 1e-06 
0.0 0.0431999999998 0 2.0 1e-06 
0.0 0.0432999999998 0 2.0 1e-06 
0.0 0.0433999999998 0 2.0 1e-06 
0.0 0.0434999999998 0 2.0 1e-06 
0.0 0.0435999999998 0 2.0 1e-06 
0.0 0.0436999999998 0 2.0 1e-06 
0.0 0.0437999999998 0 2.0 1e-06 
0.0 0.0438999999998 0 2.0 1e-06 
0.0 0.0439999999998 0 2.0 1e-06 
0.0 0.0440999999998 0 2.0 1e-06 
0.0 0.0441999999998 0 2.0 1e-06 
0.0 0.0442999999998 0 2.0 1e-06 
0.0 0.0443999999998 0 2.0 1e-06 
0.0 0.0444999999998 0 2.0 1e-06 
0.0 0.0445999999998 0 2.0 1e-06 
0.0 0.0446999999998 0 2.0 1e-06 
0.0 0.0447999999998 0 2.0 1e-06 
0.0 0.0448999999998 0 2.0 1e-06 
0.0 0.0449999999998 0 2.0 1e-06 
0.0 0.0450999999998 0 2.0 1e-06 
0.0 0.0451999999998 0 2.0 1e-06 
0.0 0.0452999999998 0 2.0 1e-06 
0.0 0.0453999999998 0 2.0 1e-06 
0.0 0.0454999999998 0 2.0 1e-06 
0.0 0.0455999999998 0 2.0 1e-06 
0.0 0.0456999999998 0 2.0 1e-06 
0.0 0.0457999999998 0 2.0 1e-06 
0.0 0.0458999999998 0 2.0 1e-06 
0.0 0.0459999999998 0 2.0 1e-06 
0.0 0.0460999999998 0 2.0 1e-06 
0.0 0.0461999999998 0 2.0 1e-06 
0.0 0.0462999999998 0 2.0 1e-06 
0.0 0.0463999999998 0 2.0 1e-06 
0.0 0.0464999999998 0 2.0 1e-06 
0.0 0.0465999999998 0 2.0 1e-06 
0.0 0.0466999999998 0 2.0 1e-06 
0.0 0.0467999999998 0 2.0 1e-06 
0.0 0.0468999999998 0 2.0 1e-06 
0.0 0.0469999999998 0 2.0 1e-06 
0.0 0.0470999999998 0 2.0 1e-06 
0.0 0.0471999999998 0 2.0 1e-06 
0.0 0.0472999999998 0 2.0 1e-06 
0.0 0.0473999999998 0 2.0 1e-06 
0.0 0.0474999999998 0 2.0 1e-06 
0.0 0.0475999999998 0 2.0 1e-06 
0.0 0.0476999999998 0 2.0 1e-06 
0.0 0.0477999999998 0 2.0 1e-06 
0.0 0.0478999999998 0 2.0 1e-06 
0.0 0.0479999999998 0 2.0 1e-06 
0.0 0.0480999999998 0 2.0 1e-06 
0.0 0.0481999999998 0 2.0 1e-06 
0.0 0.0482999999998 0 2.0 1e-06 
0.0 0.0483999999998 0 2.0 1e-06 
0.0 0.0484999999998 0 2.0 1e-06 
0.0 0.0485999999998 0 2.0 1e-06 
0.0 0.0486999999998 0 2.0 1e-06 
0.0 0.0487999999998 0 2.0 1e-06 
0.0 0.0488999999998 0 2.0 1e-06 
0.0 0.0489999999998 0 2.0 1e-06 
0.0 0.0490999999998 0 2.0 1e-06 
0.0 0.0491999999998 0 2.0 1e-06 
0.0 0.0492999999998 0 2.0 1e-06 
0.0 0.0493999999998 0 2.0 1e-06 
0.0 0.0494999999998 0 2.0 1e-06 
0.0 0.0495999999998 0 2.0 1e-06 
0.0 0.0496999999998 0 2.0 1e-06 
0.0 0.0497999999998 0 2.0 1e-06 
0.0 0.0498999999998 0 2.0 1e-06 
0.0 0.0499999999998 0 2.0 1e-06 
0.0 0.0500999999998 0 2.0 1e-06 
0.0 0.0501999999998 0 2.0 1e-06 
0.0 0.0502999999998 0 2.0 1e-06 
0.0 0.0503999999998 0 2.0 1e-06 
0.0 0.0504999999998 0 2.0 1e-06 
0.0 0.0505999999998 0 2.0 1e-06 
0.0 0.0506999999998 0 2.0 1e-06 
0.0 0.0507999999998 0 2.0 1e-06 
0.0 0.0508999999998 0 2.0 1e-06 
0.0 0.0509999999998 0 2.0 1e-06 
0.0 0.0510999999998 0 2.0 1e-06 
0.0 0.0511999999998 0 2.0 1e-06 
0.0 0.0512999999998 0 2.0 1e-06 
0.0 0.0513999999998 0 2.0 1e-06 
0.0 0.0514999999998 0 2.0 1e-06 
0.0 0.0515999999998 0 2.0 1e-06 
0.0 0.0516999999998 0 2.0 1e-06 
0.0 0.0517999999998 0 2.0 1e-06 
0.0 0.0518999999998 0 2.0 1e-06 
0.0 0.0519999999998 0 2.0 1e-06 
0.0 0.0520999999998 0 2.0 1e-06 
0.0 0.0521999999998 0 2.0 1e-06 
0.0 0.0522999999998 0 2.0 1e-06 
0.0 0.0523999999998 0 2.0 1e-06 
0.0 0.0524999999998 0 2.0 1e-06 
0.0 0.0525999999998 0 2.0 1e-06 
0.0 0.0526999999998 0 2.0 1e-06 
0.0 0.0527999999998 0 2.0 1e-06 
0.0 0.0528999999998 0 2.0 1e-06 
0.0 0.0529999999998 0 2.0 1e-06 
0.0 0.0530999999998 0 2.0 1e-06 
0.0 0.0531999999998 0 2.0 1e-06 
0.0 0.0532999999998 0 2.0 1e-06 
0.0 0.0533999999998 0 2.0 1e-06 
0.0 0.0534999999998 0 2.0 1e-06 
0.0 0.0535999999998 0 2.0 1e-06 
0.0 0.0536999999998 0 2.0 1e-06 
0.0 0.0537999999998 0 2.0 1e-06 
0.0 0.0538999999998 0 2.0 1e-06 
0.0 0.0539999999998 0 2.0 1e-06 
0.0 0.0540999999998 0 2.0 1e-06 
0.0 0.0541999999998 0 2.0 1e-06 
0.0 0.0542999999998 0 2.0 1e-06 
0.0 0.0543999999998 0 2.0 1e-06 
0.0 0.0544999999998 0 2.0 1e-06 
0.0 0.0545999999998 0 2.0 1e-06 
0.0 0.0546999999998 0 2.0 1e-06 
0.0 0.0547999999998 0 2.0 1e-06 
0.0 0.0548999999998 0 2.0 1e-06 
0.0 0.0549999999998 0 2.0 1e-06 
0.0 0.0550999999998 0 2.0 1e-06 
0.0 0.0551999999998 0 2.0 1e-06 
0.0 0.0552999999998 0 2.0 1e-06 
0.0 0.0553999999998 0 2.0 1e-06 
0.0 0.0554999999998 0 2.0 1e-06 
0.0 0.0555999999998 0 2.0 1e-06 
0.0 0.0556999999998 0 2.0 1e-06 
0.0 0.0557999999998 0 2.0 1e-06 
0.0 0.0558999999998 0 2.0 1e-06 
0.0 0.0559999999998 0 2.0 1e-06 
0.0 0.0560999999998 0 2.0 1e-06 
0.0 0.0561999999998 0 2.0 1e-06 
0.0 0.0562999999998 0 2.0 1e-06 
0.0 0.0563999999998 0 2.0 1e-06 
0.0 0.0564999999998 0 2.0 1e-06 
0.0 0.0565999999998 0 2.0 1e-06 
0.0 0.0566999999998 0 2.0 1e-06 
0.0 0.0567999999998 0 2.0 1e-06 
0.0 0.0568999999998 0 2.0 1e-06 
0.0 0.0569999999998 0 2.0 1e-06 
0.0 0.0570999999998 0 2.0 1e-06 
0.0 0.0571999999998 0 2.0 1e-06 
0.0 0.0572999999998 0 2.0 1e-06 
0.0 0.0573999999998 0 2.0 1e-06 
0.0 0.0574999999998 0 2.0 1e-06 
0.0 0.0575999999998 0 2.0 1e-06 
0.0 0.0576999999998 0 2.0 1e-06 
0.0 0.0577999999998 0 2.0 1e-06 
0.0 0.0578999999998 0 2.0 1e-06 
0.0 0.0579999999998 0 2.0 1e-06 
0.0 0.0580999999998 0 2.0 1e-06 
0.0 0.0581999999998 0 2.0 1e-06 
0.0 0.0582999999998 0 2.0 1e-06 
0.0 0.0583999999998 0 2.0 1e-06 
0.0 0.0584999999998 0 2.0 1e-06 
0.0 0.0585999999998 0 2.0 1e-06 
0.0 0.0586999999998 0 2.0 1e-06 
0.0 0.0587999999998 0 2.0 1e-06 
0.0 0.0588999999998 0 2.0 1e-06 
0.0 0.0589999999998 0 2.0 1e-06 
0.0 0.0590999999998 0 2.0 1e-06 
0.0 0.0591999999998 0 2.0 1e-06 
0.0 0.0592999999998 0 2.0 1e-06 
0.0 0.0593999999998 0 2.0 1e-06 
0.0 0.0594999999998 0 2.0 1e-06 
0.0 0.0595999999998 0 2.0 1e-06 
0.0 0.0596999999998 0 2.0 1e-06 
0.0 0.0597999999998 0 2.0 1e-06 
0.0 0.0598999999998 0 2.0 1e-06 
0.0 0.0599999999998 0 2.0 1e-06 
0.0 0.0600999999998 0 2.0 1e-06 
0.0 0.0601999999998 0 2.0 1e-06 
0.0 0.0602999999998 0 2.0 1e-06 
0.0 0.0603999999998 0 2.0 1e-06 
0.0 0.0604999999998 0 2.0 1e-06 
0.0 0.0605999999998 0 2.0 1e-06 
0.0 0.0606999999998 0 2.0 1e-06 
0.0 0.0607999999998 0 2.0 1e-06 
0.0 0.0608999999998 0 2.0 1e-06 
0.0 0.0609999999998 0 2.0 1e-06 
0.0 0.0610999999998 0 2.0 1e-06 
0.0 0.0611999999998 0 2.0 1e-06 
0.0 0.0612999999998 0 2.0 1e-06 
0.0 0.0613999999998 0 2.0 1e-06 
0.0 0.0614999999998 0 2.0 1e-06 
0.0 0.0615999999998 0 2.0 1e-06 
0.0 0.0616999999998 0 2.0 1e-06 
0.0 0.0617999999998 0 2.0 1e-06 
0.0 0.0618999999998 0 2.0 1e-06 
0.0 0.0619999999998 0 2.0 1e-06 
0.0 0.0620999999998 0 2.0 1e-06 
0.0 0.0621999999998 0 2.0 1e-06 
0.0 0.0622999999998 0 2.0 1e-06 
0.0 0.0623999999998 0 2.0 1e-06 
0.0 0.0624999999998 0 2.0 1e-06 
0.0 0.0625999999998 0 2.0 1e-06 
0.0 0.0626999999998 0 2.0 1e-06 
0.0 0.0627999999998 0 2.0 1e-06 
0.0 0.0628999999998 0 2.0 1e-06 
0.0 0.0629999999998 0 2.0 1e-06 
0.0 0.0630999999998 0 2.0 1e-06 
0.0 0.0631999999998 0 2.0 1e-06 
0.0 0.0632999999998 0 2.0 1e-06 
0.0 0.0633999999998 0 2.0 1e-06 
0.0 0.0634999999998 0 2.0 1e-06 
0.0 0.0635999999998 0 2.0 1e-06 
0.0 0.0636999999998 0 2.0 1e-06 
0.0 0.0637999999998 0 2.0 1e-06 
0.0 0.0638999999998 0 2.0 1e-06 
0.0 0.0639999999998 0 2.0 1e-06 
0.0 0.0640999999998 0 2.0 1e-06 
0.0 0.0641999999998 0 2.0 1e-06 
0.0 0.0642999999998 0 2.0 1e-06 
0.0 0.0643999999998 0 2.0 1e-06 
0.0 0.0644999999998 0 2.0 1e-06 
0.0 0.0645999999998 0 2.0 1e-06 
0.0 0.0646999999998 0 2.0 1e-06 
0.0 0.0647999999998 0 2.0 1e-06 
0.0 0.0648999999998 0 2.0 1e-06 
0.0 0.0649999999998 0 2.0 1e-06 
0.0 0.0650999999998 0 2.0 1e-06 
0.0 0.0651999999998 0 2.0 1e-06 
0.0 0.0652999999998 0 2.0 1e-06 
0.0 0.0653999999998 0 2.0 1e-06 
0.0 0.0654999999998 0 2.0 1e-06 
0.0 0.0655999999998 0 2.0 1e-06 
0.0 0.0656999999998 0 2.0 1e-06 
0.0 0.0657999999998 0 2.0 1e-06 
0.0 0.0658999999998 0 2.0 1e-06 
0.0 0.0659999999998 0 2.0 1e-06 
0.0 0.0660999999998 0 2.0 1e-06 
0.0 0.0661999999998 0 2.0 1e-06 
0.0 0.0662999999998 0 2.0 1e-06 
0.0 0.0663999999998 0 2.0 1e-06 
0.0 0.0664999999998 0 2.0 1e-06 
0.0 0.0665999999998 0 2.0 1e-06 
0.0 0.0666999999998 0 2.0 1e-06 
0.0 0.0667999999998 0 2.0 1e-06 
0.0 0.0668999999998 0 2.0 1e-06 
0.0 0.0669999999998 0 2.0 1e-06 
0.0 0.0670999999998 0 2.0 1e-06 
0.0 0.0671999999998 0 2.0 1e-06 
0.0 0.0672999999998 0 2.0 1e-06 
0.0 0.0673999999998 0 2.0 1e-06 
0.0 0.0674999999998 0 2.0 1e-06 
0.0 0.0675999999998 0 2.0 1e-06 
0.0 0.0676999999998 0 2.0 1e-06 
0.0 0.0677999999998 0 2.0 1e-06 
0.0 0.0678999999998 0 2.0 1e-06 
0.0 0.0679999999998 0 2.0 1e-06 
0.0 0.0680999999998 0 2.0 1e-06 
0.0 0.0681999999998 0 2.0 1e-06 
0.0 0.0682999999998 0 2.0 1e-06 
0.0 0.0683999999998 0 2.0 1e-06 
0.0 0.0684999999998 0 2.0 1e-06 
0.0 0.0685999999998 0 2.0 1e-06 
0.0 0.0686999999998 0 2.0 1e-06 
0.0 0.0687999999998 0 2.0 1e-06 
0.0 0.0688999999998 0 2.0 1e-06 
0.0 0.0689999999998 0 2.0 1e-06 
0.0 0.0690999999998 0 2.0 1e-06 
0.0 0.0691999999998 0 2.0 1e-06 
0.0 0.0692999999998 0 2.0 1e-06 
0.0 0.0693999999998 0 2.0 1e-06 
0.0 0.0694999999998 0 2.0 1e-06 
0.0 0.0695999999998 0 2.0 1e-06 
0.0 0.0696999999998 0 2.0 1e-06 
0.0 0.0697999999998 0 2.0 1e-06 
0.0 0.0698999999998 0 2.0 1e-06 
0.0 0.0699999999998 0 2.0 1e-06 
0.0 0.0700999999998 0 2.0 1e-06 
0.0 0.0701999999998 0 2.0 1e-06 
0.0 0.0702999999998 0 2.0 1e-06 
0.0 0.0703999999998 0 2.0 1e-06 
0.0 0.0704999999998 0 2.0 1e-06 
0.0 0.0705999999998 0 2.0 1e-06 
0.0 0.0706999999998 0 2.0 1e-06 
0.0 0.0707999999998 0 2.0 1e-06 
0.0 0.0708999999998 0 2.0 1e-06 
0.0 0.0709999999998 0 2.0 1e-06 
0.0 0.0710999999998 0 2.0 1e-06 
0.0 0.0711999999998 0 2.0 1e-06 
0.0 0.0712999999998 0 2.0 1e-06 
0.0 0.0713999999998 0 2.0 1e-06 
0.0 0.0714999999998 0 2.0 1e-06 
0.0 0.0715999999998 0 2.0 1e-06 
0.0 0.0716999999998 0 2.0 1e-06 
0.0 0.0717999999998 0 2.0 1e-06 
0.0 0.0718999999998 0 2.0 1e-06 
0.0 0.0719999999998 0 2.0 1e-06 
0.0 0.0720999999998 0 2.0 1e-06 
0.0 0.0721999999998 0 2.0 1e-06 
0.0 0.0722999999998 0 2.0 1e-06 
0.0 0.0723999999998 0 2.0 1e-06 
0.0 0.0724999999998 0 2.0 1e-06 
0.0 0.0725999999998 0 2.0 1e-06 
0.0 0.0726999999998 0 2.0 1e-06 
0.0 0.0727999999998 0 2.0 1e-06 
0.0 0.0728999999998 0 2.0 1e-06 
0.0 0.0729999999998 0 2.0 1e-06 
0.0 0.0730999999998 0 2.0 1e-06 
0.0 0.0731999999998 0 2.0 1e-06 
0.0 0.0732999999998 0 2.0 1e-06 
0.0 0.0733999999998 0 2.0 1e-06 
0.0 0.0734999999998 0 2.0 1e-06 
0.0 0.0735999999998 0 2.0 1e-06 
0.0 0.0736999999998 0 2.0 1e-06 
0.0 0.0737999999998 0 2.0 1e-06 
0.0 0.0738999999998 0 2.0 1e-06 
0.0 0.0739999999998 0 2.0 1e-06 
0.0 0.0740999999998 0 2.0 1e-06 
0.0 0.0741999999998 0 2.0 1e-06 
0.0 0.0742999999998 0 2.0 1e-06 
0.0 0.0743999999998 0 2.0 1e-06 
0.0 0.0744999999998 0 2.0 1e-06 
0.0 0.0745999999998 0 2.0 1e-06 
0.0 0.0746999999998 0 2.0 1e-06 
0.0 0.0747999999998 0 2.0 1e-06 
0.0 0.0748999999998 0 2.0 1e-06 
0.0 0.0749999999998 0 2.0 1e-06 
0.0 0.0750999999998 0 2.0 1e-06 
0.0 0.0751999999998 0 2.0 1e-06 
0.0 0.0752999999998 0 2.0 1e-06 
0.0 0.0753999999998 0 2.0 1e-06 
0.0 0.0754999999998 0 2.0 1e-06 
0.0 0.0755999999998 0 2.0 1e-06 
0.0 0.0756999999998 0 2.0 1e-06 
0.0 0.0757999999998 0 2.0 1e-06 
0.0 0.0758999999998 0 2.0 1e-06 
0.0 0.0759999999998 0 2.0 1e-06 
0.0 0.0760999999998 0 2.0 1e-06 
0.0 0.0761999999998 0 2.0 1e-06 
0.0 0.0762999999998 0 2.0 1e-06 
0.0 0.0763999999998 0 2.0 1e-06 
0.0 0.0764999999998 0 2.0 1e-06 
0.0 0.0765999999998 0 2.0 1e-06 
0.0 0.0766999999998 0 2.0 1e-06 
0.0 0.0767999999998 0 2.0 1e-06 
0.0 0.0768999999998 0 2.0 1e-06 
0.0 0.0769999999998 0 2.0 1e-06 
0.0 0.0770999999998 0 2.0 1e-06 
0.0 0.0771999999998 0 2.0 1e-06 
0.0 0.0772999999998 0 2.0 1e-06 
0.0 0.0773999999998 0 2.0 1e-06 
0.0 0.0774999999998 0 2.0 1e-06 
0.0 0.0775999999998 0 2.0 1e-06 
0.0 0.0776999999998 0 2.0 1e-06 
0.0 0.0777999999998 0 2.0 1e-06 
0.0 0.0778999999998 0 2.0 1e-06 
0.0 0.0779999999998 0 2.0 1e-06 
0.0 0.0780999999998 0 2.0 1e-06 
0.0 0.0781999999998 0 2.0 1e-06 
0.0 0.0782999999998 0 2.0 1e-06 
0.0 0.0783999999998 0 2.0 1e-06 
0.0 0.0784999999998 0 2.0 1e-06 
0.0 0.0785999999998 0 2.0 1e-06 
0.0 0.0786999999998 0 2.0 1e-06 
0.0 0.0787999999998 0 2.0 1e-06 
0.0 0.0788999999998 0 2.0 1e-06 
0.0 0.0789999999998 0 2.0 1e-06 
0.0 0.0790999999998 0 2.0 1e-06 
0.0 0.0791999999998 0 2.0 1e-06 
0.0 0.0792999999998 0 2.0 1e-06 
0.0 0.0793999999998 0 2.0 1e-06 
0.0 0.0794999999998 0 2.0 1e-06 
0.0 0.0795999999998 0 2.0 1e-06 
0.0 0.0796999999998 0 2.0 1e-06 
0.0 0.0797999999998 0 2.0 1e-06 
0.0 0.0798999999998 0 2.0 1e-06 
0.0 0.0799999999998 0 2.0 1e-06 
0.0 0.0800999999998 0 2.0 1e-06 
0.0 0.0801999999998 0 2.0 1e-06 
0.0 0.0802999999998 0 2.0 1e-06 
0.0 0.0803999999998 0 2.0 1e-06 
0.0 0.0804999999998 0 2.0 1e-06 
0.0 0.0805999999998 0 2.0 1e-06 
0.0 0.0806999999998 0 2.0 1e-06 
0.0 0.0807999999998 0 2.0 1e-06 
0.0 0.0808999999998 0 2.0 1e-06 
0.0 0.0809999999998 0 2.0 1e-06 
0.0 0.0810999999998 0 2.0 1e-06 
0.0 0.0811999999998 0 2.0 1e-06 
0.0 0.0812999999998 0 2.0 1e-06 
0.0 0.0813999999998 0 2.0 1e-06 
0.0 0.0814999999998 0 2.0 1e-06 
0.0 0.0815999999998 0 2.0 1e-06 
0.0 0.0816999999998 0 2.0 1e-06 
0.0 0.0817999999998 0 2.0 1e-06 
0.0 0.0818999999998 0 2.0 1e-06 
0.0 0.0819999999998 0 2.0 1e-06 
0.0 0.0820999999998 0 2.0 1e-06 
0.0 0.0821999999998 0 2.0 1e-06 
0.0 0.0822999999998 0 2.0 1e-06 
0.0 0.0823999999998 0 2.0 1e-06 
0.0 0.0824999999998 0 2.0 1e-06 
0.0 0.0825999999998 0 2.0 1e-06 
0.0 0.0826999999998 0 2.0 1e-06 
0.0 0.0827999999998 0 2.0 1e-06 
0.0 0.0828999999998 0 2.0 1e-06 
0.0 0.0829999999998 0 2.0 1e-06 
0.0 0.0830999999998 0 2.0 1e-06 
0.0 0.0831999999998 0 2.0 1e-06 
0.0 0.0832999999998 0 2.0 1e-06 
0.0 0.0833999999998 0 2.0 1e-06 
0.0 0.0834999999998 0 2.0 1e-06 
0.0 0.0835999999998 0 2.0 1e-06 
0.0 0.0836999999998 0 2.0 1e-06 
0.0 0.0837999999998 0 2.0 1e-06 
0.0 0.0838999999998 0 2.0 1e-06 
0.0 0.0839999999998 0 2.0 1e-06 
0.0 0.0840999999998 0 2.0 1e-06 
0.0 0.0841999999998 0 2.0 1e-06 
0.0 0.0842999999998 0 2.0 1e-06 
0.0 0.0843999999998 0 2.0 1e-06 
0.0 0.0844999999998 0 2.0 1e-06 
0.0 0.0845999999998 0 2.0 1e-06 
0.0 0.0846999999998 0 2.0 1e-06 
0.0 0.0847999999998 0 2.0 1e-06 
0.0 0.0848999999998 0 2.0 1e-06 
0.0 0.0849999999998 0 2.0 1e-06 
0.0 0.0850999999998 0 2.0 1e-06 
0.0 0.0851999999998 0 2.0 1e-06 
0.0 0.0852999999998 0 2.0 1e-06 
0.0 0.0853999999998 0 2.0 1e-06 
0.0 0.0854999999998 0 2.0 1e-06 
0.0 0.0855999999998 0 2.0 1e-06 
0.0 0.0856999999998 0 2.0 1e-06 
0.0 0.0857999999998 0 2.0 1e-06 
0.0 0.0858999999998 0 2.0 1e-06 
0.0 0.0859999999998 0 2.0 1e-06 
0.0 0.0860999999998 0 2.0 1e-06 
0.0 0.0861999999998 0 2.0 1e-06 
0.0 0.0862999999998 0 2.0 1e-06 
0.0 0.0863999999998 0 2.0 1e-06 
0.0 0.0864999999998 0 2.0 1e-06 
0.0 0.0865999999998 0 2.0 1e-06 
0.0 0.0866999999998 0 2.0 1e-06 
0.0 0.0867999999998 0 2.0 1e-06 
0.0 0.0868999999998 0 2.0 1e-06 
0.0 0.0869999999998 0 2.0 1e-06 
0.0 0.0870999999998 0 2.0 1e-06 
0.0 0.0871999999998 0 2.0 1e-06 
0.0 0.0872999999998 0 2.0 1e-06 
0.0 0.0873999999998 0 2.0 1e-06 
0.0 0.0874999999998 0 2.0 1e-06 
0.0 0.0875999999998 0 2.0 1e-06 
0.0 0.0876999999998 0 2.0 1e-06 
0.0 0.0877999999998 0 2.0 1e-06 
0.0 0.0878999999998 0 2.0 1e-06 
0.0 0.0879999999998 0 2.0 1e-06 
0.0 0.0880999999998 0 2.0 1e-06 
0.0 0.0881999999998 0 2.0 1e-06 
0.0 0.0882999999998 0 2.0 1e-06 
0.0 0.0883999999998 0 2.0 1e-06 
0.0 0.0884999999998 0 2.0 1e-06 
0.0 0.0885999999998 0 2.0 1e-06 
0.0 0.0886999999998 0 2.0 1e-06 
0.0 0.0887999999998 0 2.0 1e-06 
0.0 0.0888999999998 0 2.0 1e-06 
0.0 0.0889999999998 0 2.0 1e-06 
0.0 0.0890999999998 0 2.0 1e-06 
0.0 0.0891999999998 0 2.0 1e-06 
0.0 0.0892999999998 0 2.0 1e-06 
0.0 0.0893999999998 0 2.0 1e-06 
0.0 0.0894999999998 0 2.0 1e-06 
0.0 0.0895999999998 0 2.0 1e-06 
0.0 0.0896999999998 0 2.0 1e-06 
0.0 0.0897999999998 0 2.0 1e-06 
0.0 0.0898999999998 0 2.0 1e-06 
0.0 0.0899999999998 0 2.0 1e-06 
0.0 0.0900999999998 0 2.0 1e-06 
0.0 0.0901999999998 0 2.0 1e-06 
0.0 0.0902999999998 0 2.0 1e-06 
0.0 0.0903999999998 0 2.0 1e-06 
0.0 0.0904999999998 0 2.0 1e-06 
0.0 0.0905999999998 0 2.0 1e-06 
0.0 0.0906999999998 0 2.0 1e-06 
0.0 0.0907999999998 0 2.0 1e-06 
0.0 0.0908999999998 0 2.0 1e-06 
0.0 0.0909999999998 0 2.0 1e-06 
0.0 0.0910999999998 0 2.0 1e-06 
0.0 0.0911999999998 0 2.0 1e-06 
0.0 0.0912999999998 0 2.0 1e-06 
0.0 0.0913999999998 0 2.0 1e-06 
0.0 0.0914999999998 0 2.0 1e-06 
0.0 0.0915999999998 0 2.0 1e-06 
0.0 0.0916999999998 0 2.0 1e-06 
0.0 0.0917999999998 0 2.0 1e-06 
0.0 0.0918999999998 0 2.0 1e-06 
0.0 0.0919999999998 0 2.0 1e-06 
0.0 0.0920999999998 0 2.0 1e-06 
0.0 0.0921999999998 0 2.0 1e-06 
0.0 0.0922999999998 0 2.0 1e-06 
0.0 0.0923999999998 0 2.0 1e-06 
0.0 0.0924999999998 0 2.0 1e-06 
0.0 0.0925999999998 0 2.0 1e-06 
0.0 0.0926999999998 0 2.0 1e-06 
0.0 0.0927999999998 0 2.0 1e-06 
0.0 0.0928999999998 0 2.0 1e-06 
0.0 0.0929999999998 0 2.0 1e-06 
0.0 0.0930999999998 0 2.0 1e-06 
0.0 0.0931999999998 0 2.0 1e-06 
0.0 0.0932999999998 0 2.0 1e-06 
0.0 0.0933999999998 0 2.0 1e-06 
0.0 0.0934999999998 0 2.0 1e-06 
0.0 0.0935999999998 0 2.0 1e-06 
0.0 0.0936999999998 0 2.0 1e-06 
0.0 0.0937999999998 0 2.0 1e-06 
0.0 0.0938999999998 0 2.0 1e-06 
0.0 0.0939999999998 0 2.0 1e-06 
0.0 0.0940999999998 0 2.0 1e-06 
0.0 0.0941999999998 0 2.0 1e-06 
0.0 0.0942999999998 0 2.0 1e-06 
0.0 0.0943999999998 0 2.0 1e-06 
0.0 0.0944999999998 0 2.0 1e-06 
0.0 0.0945999999998 0 2.0 1e-06 
0.0 0.0946999999998 0 2.0 1e-06 
0.0 0.0947999999998 0 2.0 1e-06 
0.0 0.0948999999998 0 2.0 1e-06 
0.0 0.0949999999998 0 2.0 1e-06 
0.0 0.0950999999998 0 2.0 1e-06 
0.0 0.0951999999998 0 2.0 1e-06 
0.0 0.0952999999998 0 2.0 1e-06 
0.0 0.0953999999998 0 2.0 1e-06 
0.0 0.0954999999998 0 2.0 1e-06 
0.0 0.0955999999998 0 2.0 1e-06 
0.0 0.0956999999998 0 2.0 1e-06 
0.0 0.0957999999998 0 2.0 1e-06 
0.0 0.0958999999998 0 2.0 1e-06 
0.0 0.0959999999998 0 2.0 1e-06 
0.0 0.0960999999998 0 2.0 1e-06 
0.0 0.0961999999998 0 2.0 1e-06 
0.0 0.0962999999998 0 2.0 1e-06 
0.0 0.0963999999998 0 2.0 1e-06 
0.0 0.0964999999998 0 2.0 1e-06 
0.0 0.0965999999998 0 2.0 1e-06 
0.0 0.0966999999998 0 2.0 1e-06 
0.0 0.0967999999998 0 2.0 1e-06 
0.0 0.0968999999998 0 2.0 1e-06 
0.0 0.0969999999998 0 2.0 1e-06 
0.0 0.0970999999998 0 2.0 1e-06 
0.0 0.0971999999998 0 2.0 1e-06 
0.0 0.0972999999998 0 2.0 1e-06 
0.0 0.0973999999998 0 2.0 1e-06 
0.0 0.0974999999998 0 2.0 1e-06 
0.0 0.0975999999998 0 2.0 1e-06 
0.0 0.0976999999998 0 2.0 1e-06 
0.0 0.0977999999998 0 2.0 1e-06 
0.0 0.0978999999998 0 2.0 1e-06 
0.0 0.0979999999998 0 2.0 1e-06 
0.0 0.0980999999998 0 2.0 1e-06 
0.0 0.0981999999998 0 2.0 1e-06 
0.0 0.0982999999998 0 2.0 1e-06 
0.0 0.0983999999998 0 2.0 1e-06 
0.0 0.0984999999998 0 2.0 1e-06 
0.0 0.0985999999998 0 2.0 1e-06 
0.0 0.0986999999998 0 2.0 1e-06 
0.0 0.0987999999998 0 2.0 1e-06 
0.0 0.0988999999998 0 2.0 1e-06 
0.0 0.0989999999998 0 2.0 1e-06 
0.0 0.0990999999998 0 2.0 1e-06 
0.0 0.0991999999998 0 2.0 1e-06 
0.0 0.0992999999998 0 2.0 1e-06 
0.0 0.0993999999998 0 2.0 1e-06 
0.0 0.0994999999998 0 2.0 1e-06 
0.0 0.0995999999998 0 2.0 1e-06 
0.0 0.0996999999998 0 2.0 1e-06 
0.0 0.0997999999998 0 2.0 1e-06 
0.0 0.0998999999998 0 2.0 1e-06 
0.0 0.0999999999998 0 2.0 1e-06 
0.0 0.1001 0 2.0 1e-06 
0.0 0.1002 0 2.0 1e-06 
0.0 0.1003 0 2.0 1e-06 
0.0 0.1004 0 2.0 1e-06 
0.0 0.1005 0 2.0 1e-06 
0.0 0.1006 0 2.0 1e-06 
0.0 0.1007 0 2.0 1e-06 
0.0 0.1008 0 2.0 1e-06 
0.0 0.1009 0 2.0 1e-06 
0.0 0.101 0 2.0 1e-06 
0.0 0.1011 0 2.0 1e-06 
0.0 0.1012 0 2.0 1e-06 
0.0 0.1013 0 2.0 1e-06 
0.0 0.1014 0 2.0 1e-06 
0.0 0.1015 0 2.0 1e-06 
0.0 0.1016 0 2.0 1e-06 
0.0 0.1017 0 2.0 1e-06 
0.0 0.1018 0 2.0 1e-06 
0.0 0.1019 0 2.0 1e-06 
0.0 0.102 0 2.0 1e-06 
0.0 0.1021 0 2.0 1e-06 
0.0 0.1022 0 2.0 1e-06 
0.0 0.1023 0 2.0 1e-06 
0.0 0.1024 0 2.0 1e-06 
0.0 0.1025 0 2.0 1e-06 
0.0 0.1026 0 2.0 1e-06 
0.0 0.1027 0 2.0 1e-06 
0.0 0.1028 0 2.0 1e-06 
0.0 0.1029 0 2.0 1e-06 
0.0 0.103 0 2.0 1e-06 
0.0 0.1031 0 2.0 1e-06 
0.0 0.1032 0 2.0 1e-06 
0.0 0.1033 0 2.0 1e-06 
0.0 0.1034 0 2.0 1e-06 
0.0 0.1035 0 2.0 1e-06 
0.0 0.1036 0 2.0 1e-06 
0.0 0.1037 0 2.0 1e-06 
0.0 0.1038 0 2.0 1e-06 
0.0 0.1039 0 2.0 1e-06 
0.0 0.104 0 2.0 1e-06 
0.0 0.1041 0 2.0 1e-06 
0.0 0.1042 0 2.0 1e-06 
0.0 0.1043 0 2.0 1e-06 
0.0 0.1044 0 2.0 1e-06 
0.0 0.1045 0 2.0 1e-06 
0.0 0.1046 0 2.0 1e-06 
0.0 0.1047 0 2.0 1e-06 
0.0 0.1048 0 2.0 1e-06 
0.0 0.1049 0 2.0 1e-06 
0.0 0.105 0 2.0 1e-06 
0.0 0.1051 0 2.0 1e-06 
0.0 0.1052 0 2.0 1e-06 
0.0 0.1053 0 2.0 1e-06 
0.0 0.1054 0 2.0 1e-06 
0.0 0.1055 0 2.0 1e-06 
0.0 0.1056 0 2.0 1e-06 
0.0 0.1057 0 2.0 1e-06 
0.0 0.1058 0 2.0 1e-06 
0.0 0.1059 0 2.0 1e-06 
0.0 0.106 0 2.0 1e-06 
0.0 0.1061 0 2.0 1e-06 
0.0 0.1062 0 2.0 1e-06 
0.0 0.1063 0 2.0 1e-06 
0.0 0.1064 0 2.0 1e-06 
0.0 0.1065 0 2.0 1e-06 
0.0 0.1066 0 2.0 1e-06 
0.0 0.1067 0 2.0 1e-06 
0.0 0.1068 0 2.0 1e-06 
0.0 0.1069 0 2.0 1e-06 
0.0 0.107 0 2.0 1e-06 
0.0 0.1071 0 2.0 1e-06 
0.0 0.1072 0 2.0 1e-06 
0.0 0.1073 0 2.0 1e-06 
0.0 0.1074 0 2.0 1e-06 
0.0 0.1075 0 2.0 1e-06 
0.0 0.1076 0 2.0 1e-06 
0.0 0.1077 0 2.0 1e-06 
0.0 0.1078 0 2.0 1e-06 
0.0 0.1079 0 2.0 1e-06 
0.0 0.108 0 2.0 1e-06 
0.0 0.1081 0 2.0 1e-06 
0.0 0.1082 0 2.0 1e-06 
0.0 0.1083 0 2.0 1e-06 
0.0 0.1084 0 2.0 1e-06 
0.0 0.1085 0 2.0 1e-06 
0.0 0.1086 0 2.0 1e-06 
0.0 0.1087 0 2.0 1e-06 
0.0 0.1088 0 2.0 1e-06 
0.0 0.1089 0 2.0 1e-06 
0.0 0.109 0 2.0 1e-06 
0.0 0.1091 0 2.0 1e-06 
0.0 0.1092 0 2.0 1e-06 
0.0 0.1093 0 2.0 1e-06 
0.0 0.1094 0 2.0 1e-06 
0.0 0.1095 0 2.0 1e-06 
0.0 0.1096 0 2.0 1e-06 
0.0 0.1097 0 2.0 1e-06 
0.0 0.1098 0 2.0 1e-06 
0.0 0.1099 0 2.0 1e-06 
0.0 0.11 0 2.0 1e-06 
0.0 0.1101 0 2.0 1e-06 
0.0 0.1102 0 2.0 1e-06 
0.0 0.1103 0 2.0 1e-06 
0.0 0.1104 0 2.0 1e-06 
0.0 0.1105 0 2.0 1e-06 
0.0 0.1106 0 2.0 1e-06 
0.0 0.1107 0 2.0 1e-06 
0.0 0.1108 0 2.0 1e-06 
0.0 0.1109 0 2.0 1e-06 
0.0 0.111 0 2.0 1e-06 
0.0 0.1111 0 2.0 1e-06 
0.0 0.1112 0 2.0 1e-06 
0.0 0.1113 0 2.0 1e-06 
0.0 0.1114 0 2.0 1e-06 
0.0 0.1115 0 2.0 1e-06 
0.0 0.1116 0 2.0 1e-06 
0.0 0.1117 0 2.0 1e-06 
0.0 0.1118 0 2.0 1e-06 
0.0 0.1119 0 2.0 1e-06 
0.0 0.112 0 2.0 1e-06 
0.0 0.1121 0 2.0 1e-06 
0.0 0.1122 0 2.0 1e-06 
0.0 0.1123 0 2.0 1e-06 
0.0 0.1124 0 2.0 1e-06 
0.0 0.1125 0 2.0 1e-06 
0.0 0.1126 0 2.0 1e-06 
0.0 0.1127 0 2.0 1e-06 
0.0 0.1128 0 2.0 1e-06 
0.0 0.1129 0 2.0 1e-06 
0.0 0.113 0 2.0 1e-06 
0.0 0.1131 0 2.0 1e-06 
0.0 0.1132 0 2.0 1e-06 
0.0 0.1133 0 2.0 1e-06 
0.0 0.1134 0 2.0 1e-06 
0.0 0.1135 0 2.0 1e-06 
0.0 0.1136 0 2.0 1e-06 
0.0 0.1137 0 2.0 1e-06 
0.0 0.1138 0 2.0 1e-06 
0.0 0.1139 0 2.0 1e-06 
0.0 0.114 0 2.0 1e-06 
0.0 0.1141 0 2.0 1e-06 
0.0 0.1142 0 2.0 1e-06 
0.0 0.1143 0 2.0 1e-06 
0.0 0.1144 0 2.0 1e-06 
0.0 0.1145 0 2.0 1e-06 
0.0 0.1146 0 2.0 1e-06 
0.0 0.1147 0 2.0 1e-06 
0.0 0.1148 0 2.0 1e-06 
0.0 0.1149 0 2.0 1e-06 
0.0 0.115 0 2.0 1e-06 
0.0 0.1151 0 2.0 1e-06 
0.0 0.1152 0 2.0 1e-06 
0.0 0.1153 0 2.0 1e-06 
0.0 0.1154 0 2.0 1e-06 
0.0 0.1155 0 2.0 1e-06 
0.0 0.1156 0 2.0 1e-06 
0.0 0.1157 0 2.0 1e-06 
0.0 0.1158 0 2.0 1e-06 
0.0 0.1159 0 2.0 1e-06 
0.0 0.116 0 2.0 1e-06 
0.0 0.1161 0 2.0 1e-06 
0.0 0.1162 0 2.0 1e-06 
0.0 0.1163 0 2.0 1e-06 
0.0 0.1164 0 2.0 1e-06 
0.0 0.1165 0 2.0 1e-06 
0.0 0.1166 0 2.0 1e-06 
0.0 0.1167 0 2.0 1e-06 
0.0 0.1168 0 2.0 1e-06 
0.0 0.1169 0 2.0 1e-06 
0.0 0.117 0 2.0 1e-06 
0.0 0.1171 0 2.0 1e-06 
0.0 0.1172 0 2.0 1e-06 
0.0 0.1173 0 2.0 1e-06 
0.0 0.1174 0 2.0 1e-06 
0.0 0.1175 0 2.0 1e-06 
0.0 0.1176 0 2.0 1e-06 
0.0 0.1177 0 2.0 1e-06 
0.0 0.1178 0 2.0 1e-06 
0.0 0.1179 0 2.0 1e-06 
0.0 0.118 0 2.0 1e-06 
0.0 0.1181 0 2.0 1e-06 
0.0 0.1182 0 2.0 1e-06 
0.0 0.1183 0 2.0 1e-06 
0.0 0.1184 0 2.0 1e-06 
0.0 0.1185 0 2.0 1e-06 
0.0 0.1186 0 2.0 1e-06 
0.0 0.1187 0 2.0 1e-06 
0.0 0.1188 0 2.0 1e-06 
0.0 0.1189 0 2.0 1e-06 
0.0 0.119 0 2.0 1e-06 
0.0 0.1191 0 2.0 1e-06 
0.0 0.1192 0 2.0 1e-06 
0.0 0.1193 0 2.0 1e-06 
0.0 0.1194 0 2.0 1e-06 
0.0 0.1195 0 2.0 1e-06 
0.0 0.1196 0 2.0 1e-06 
0.0 0.1197 0 2.0 1e-06 
0.0 0.1198 0 2.0 1e-06 
0.0 0.1199 0 2.0 1e-06 
0.0 0.12 0 2.0 1e-06 
0.0 0.1201 0 2.0 1e-06 
0.0 0.1202 0 2.0 1e-06 
0.0 0.1203 0 2.0 1e-06 
0.0 0.1204 0 2.0 1e-06 
0.0 0.1205 0 2.0 1e-06 
0.0 0.1206 0 2.0 1e-06 
0.0 0.1207 0 2.0 1e-06 
0.0 0.1208 0 2.0 1e-06 
0.0 0.1209 0 2.0 1e-06 
0.0 0.121 0 2.0 1e-06 
0.0 0.1211 0 2.0 1e-06 
0.0 0.1212 0 2.0 1e-06 
0.0 0.1213 0 2.0 1e-06 
0.0 0.1214 0 2.0 1e-06 
0.0 0.1215 0 2.0 1e-06 
0.0 0.1216 0 2.0 1e-06 
0.0 0.1217 0 2.0 1e-06 
0.0 0.1218 0 2.0 1e-06 
0.0 0.1219 0 2.0 1e-06 
0.0 0.122 0 2.0 1e-06 
0.0 0.1221 0 2.0 1e-06 
0.0 0.1222 0 2.0 1e-06 
0.0 0.1223 0 2.0 1e-06 
0.0 0.1224 0 2.0 1e-06 
0.0 0.1225 0 2.0 1e-06 
0.0 0.1226 0 2.0 1e-06 
0.0 0.1227 0 2.0 1e-06 
0.0 0.1228 0 2.0 1e-06 
0.0 0.1229 0 2.0 1e-06 
0.0 0.123 0 2.0 1e-06 
0.0 0.1231 0 2.0 1e-06 
0.0 0.1232 0 2.0 1e-06 
0.0 0.1233 0 2.0 1e-06 
0.0 0.1234 0 2.0 1e-06 
0.0 0.1235 0 2.0 1e-06 
0.0 0.1236 0 2.0 1e-06 
0.0 0.1237 0 2.0 1e-06 
0.0 0.1238 0 2.0 1e-06 
0.0 0.1239 0 2.0 1e-06 
0.0 0.124 0 2.0 1e-06 
0.0 0.1241 0 2.0 1e-06 
0.0 0.1242 0 2.0 1e-06 
0.0 0.1243 0 2.0 1e-06 
0.0 0.1244 0 2.0 1e-06 
0.0 0.1245 0 2.0 1e-06 
0.0 0.1246 0 2.0 1e-06 
0.0 0.1247 0 2.0 1e-06 
0.0 0.1248 0 2.0 1e-06 
0.0 0.1249 0 2.0 1e-06 
0.0 0.125 0 2.0 1e-06 
0.0 0.1251 0 2.0 1e-06 
0.0 0.1252 0 2.0 1e-06 
0.0 0.1253 0 2.0 1e-06 
0.0 0.1254 0 2.0 1e-06 
0.0 0.1255 0 2.0 1e-06 
0.0 0.1256 0 2.0 1e-06 
0.0 0.1257 0 2.0 1e-06 
0.0 0.1258 0 2.0 1e-06 
0.0 0.1259 0 2.0 1e-06 
0.0 0.126 0 2.0 1e-06 
0.0 0.1261 0 2.0 1e-06 
0.0 0.1262 0 2.0 1e-06 
0.0 0.1263 0 2.0 1e-06 
0.0 0.1264 0 2.0 1e-06 
0.0 0.1265 0 2.0 1e-06 
0.0 0.1266 0 2.0 1e-06 
0.0 0.1267 0 2.0 1e-06 
0.0 0.1268 0 2.0 1e-06 
0.0 0.1269 0 2.0 1e-06 
0.0 0.127 0 2.0 1e-06 
0.0 0.1271 0 2.0 1e-06 
0.0 0.1272 0 2.0 1e-06 
0.0 0.1273 0 2.0 1e-06 
0.0 0.1274 0 2.0 1e-06 
0.0 0.1275 0 2.0 1e-06 
0.0 0.1276 0 2.0 1e-06 
0.0 0.1277 0 2.0 1e-06 
0.0 0.1278 0 2.0 1e-06 
0.0 0.1279 0 2.0 1e-06 
0.0 0.128 0 2.0 1e-06 
0.0 0.1281 0 2.0 1e-06 
0.0 0.1282 0 2.0 1e-06 
0.0 0.1283 0 2.0 1e-06 
0.0 0.1284 0 2.0 1e-06 
0.0 0.1285 0 2.0 1e-06 
0.0 0.1286 0 2.0 1e-06 
0.0 0.1287 0 2.0 1e-06 
0.0 0.1288 0 2.0 1e-06 
0.0 0.1289 0 2.0 1e-06 
0.0 0.129 0 2.0 1e-06 
0.0 0.1291 0 2.0 1e-06 
0.0 0.1292 0 2.0 1e-06 
0.0 0.1293 0 2.0 1e-06 
0.0 0.1294 0 2.0 1e-06 
0.0 0.1295 0 2.0 1e-06 
0.0 0.1296 0 2.0 1e-06 
0.0 0.1297 0 2.0 1e-06 
0.0 0.1298 0 2.0 1e-06 
0.0 0.1299 0 2.0 1e-06 
0.0 0.13 0 2.0 1e-06 
0.0 0.1301 0 2.0 1e-06 
0.0 0.1302 0 2.0 1e-06 
0.0 0.1303 0 2.0 1e-06 
0.0 0.1304 0 2.0 1e-06 
0.0 0.1305 0 2.0 1e-06 
0.0 0.1306 0 2.0 1e-06 
0.0 0.1307 0 2.0 1e-06 
0.0 0.1308 0 2.0 1e-06 
0.0 0.1309 0 2.0 1e-06 
0.0 0.131 0 2.0 1e-06 
0.0 0.1311 0 2.0 1e-06 
0.0 0.1312 0 2.0 1e-06 
0.0 0.1313 0 2.0 1e-06 
0.0 0.1314 0 2.0 1e-06 
0.0 0.1315 0 2.0 1e-06 
0.0 0.1316 0 2.0 1e-06 
0.0 0.1317 0 2.0 1e-06 
0.0 0.1318 0 2.0 1e-06 
0.0 0.1319 0 2.0 1e-06 
0.0 0.132 0 2.0 1e-06 
0.0 0.1321 0 2.0 1e-06 
0.0 0.1322 0 2.0 1e-06 
0.0 0.1323 0 2.0 1e-06 
0.0 0.1324 0 2.0 1e-06 
0.0 0.1325 0 2.0 1e-06 
0.0 0.1326 0 2.0 1e-06 
0.0 0.1327 0 2.0 1e-06 
0.0 0.1328 0 2.0 1e-06 
0.0 0.1329 0 2.0 1e-06 
0.0 0.133 0 2.0 1e-06 
0.0 0.1331 0 2.0 1e-06 
0.0 0.1332 0 2.0 1e-06 
0.0 0.1333 0 2.0 1e-06 
0.0 0.1334 0 2.0 1e-06 
0.0 0.1335 0 2.0 1e-06 
0.0 0.1336 0 2.0 1e-06 
0.0 0.1337 0 2.0 1e-06 
0.0 0.1338 0 2.0 1e-06 
0.0 0.1339 0 2.0 1e-06 
0.0 0.134 0 2.0 1e-06 
0.0 0.1341 0 2.0 1e-06 
0.0 0.1342 0 2.0 1e-06 
0.0 0.1343 0 2.0 1e-06 
0.0 0.1344 0 2.0 1e-06 
0.0 0.1345 0 2.0 1e-06 
0.0 0.1346 0 2.0 1e-06 
0.0 0.1347 0 2.0 1e-06 
0.0 0.1348 0 2.0 1e-06 
0.0 0.1349 0 2.0 1e-06 
0.0 0.135 0 2.0 1e-06 
0.0 0.1351 0 2.0 1e-06 
0.0 0.1352 0 2.0 1e-06 
0.0 0.1353 0 2.0 1e-06 
0.0 0.1354 0 2.0 1e-06 
0.0 0.1355 0 2.0 1e-06 
0.0 0.1356 0 2.0 1e-06 
0.0 0.1357 0 2.0 1e-06 
0.0 0.1358 0 2.0 1e-06 
0.0 0.1359 0 2.0 1e-06 
0.0 0.136 0 2.0 1e-06 
0.0 0.1361 0 2.0 1e-06 
0.0 0.1362 0 2.0 1e-06 
0.0 0.1363 0 2.0 1e-06 
0.0 0.1364 0 2.0 1e-06 
0.0 0.1365 0 2.0 1e-06 
0.0 0.1366 0 2.0 1e-06 
0.0 0.1367 0 2.0 1e-06 
0.0 0.1368 0 2.0 1e-06 
0.0 0.1369 0 2.0 1e-06 
0.0 0.137 0 2.0 1e-06 
0.0 0.1371 0 2.0 1e-06 
0.0 0.1372 0 2.0 1e-06 
0.0 0.1373 0 2.0 1e-06 
0.0 0.1374 0 2.0 1e-06 
0.0 0.1375 0 2.0 1e-06 
0.0 0.1376 0 2.0 1e-06 
0.0 0.1377 0 2.0 1e-06 
0.0 0.1378 0 2.0 1e-06 
0.0 0.1379 0 2.0 1e-06 
0.0 0.138 0 2.0 1e-06 
0.0 0.1381 0 2.0 1e-06 
0.0 0.1382 0 2.0 1e-06 
0.0 0.1383 0 2.0 1e-06 
0.0 0.1384 0 2.0 1e-06 
0.0 0.1385 0 2.0 1e-06 
0.0 0.1386 0 2.0 1e-06 
0.0 0.1387 0 2.0 1e-06 
0.0 0.1388 0 2.0 1e-06 
0.0 0.1389 0 2.0 1e-06 
0.0 0.139 0 2.0 1e-06 
0.0 0.1391 0 2.0 1e-06 
0.0 0.1392 0 2.0 1e-06 
0.0 0.1393 0 2.0 1e-06 
0.0 0.1394 0 2.0 1e-06 
0.0 0.1395 0 2.0 1e-06 
0.0 0.1396 0 2.0 1e-06 
0.0 0.1397 0 2.0 1e-06 
0.0 0.1398 0 2.0 1e-06 
0.0 0.1399 0 2.0 1e-06 
0.0 0.14 0 2.0 1e-06 
0.0 0.1401 0 2.0 1e-06 
0.0 0.1402 0 2.0 1e-06 
0.0 0.1403 0 2.0 1e-06 
0.0 0.1404 0 2.0 1e-06 
0.0 0.1405 0 2.0 1e-06 
0.0 0.1406 0 2.0 1e-06 
0.0 0.1407 0 2.0 1e-06 
0.0 0.1408 0 2.0 1e-06 
0.0 0.1409 0 2.0 1e-06 
0.0 0.141 0 2.0 1e-06 
0.0 0.1411 0 2.0 1e-06 
0.0 0.1412 0 2.0 1e-06 
0.0 0.1413 0 2.0 1e-06 
0.0 0.1414 0 2.0 1e-06 
0.0 0.1415 0 2.0 1e-06 
0.0 0.1416 0 2.0 1e-06 
0.0 0.1417 0 2.0 1e-06 
0.0 0.1418 0 2.0 1e-06 
0.0 0.1419 0 2.0 1e-06 
0.0 0.142 0 2.0 1e-06 
0.0 0.1421 0 2.0 1e-06 
0.0 0.1422 0 2.0 1e-06 
0.0 0.1423 0 2.0 1e-06 
0.0 0.1424 0 2.0 1e-06 
0.0 0.1425 0 2.0 1e-06 
0.0 0.1426 0 2.0 1e-06 
0.0 0.1427 0 2.0 1e-06 
0.0 0.1428 0 2.0 1e-06 
0.0 0.1429 0 2.0 1e-06 
0.0 0.143 0 2.0 1e-06 
0.0 0.1431 0 2.0 1e-06 
0.0 0.1432 0 2.0 1e-06 
0.0 0.1433 0 2.0 1e-06 
0.0 0.1434 0 2.0 1e-06 
0.0 0.1435 0 2.0 1e-06 
0.0 0.1436 0 2.0 1e-06 
0.0 0.1437 0 2.0 1e-06 
0.0 0.1438 0 2.0 1e-06 
0.0 0.1439 0 2.0 1e-06 
0.0 0.144 0 2.0 1e-06 
0.0 0.1441 0 2.0 1e-06 
0.0 0.1442 0 2.0 1e-06 
0.0 0.1443 0 2.0 1e-06 
0.0 0.1444 0 2.0 1e-06 
0.0 0.1445 0 2.0 1e-06 
0.0 0.1446 0 2.0 1e-06 
0.0 0.1447 0 2.0 1e-06 
0.0 0.1448 0 2.0 1e-06 
0.0 0.1449 0 2.0 1e-06 
0.0 0.145 0 2.0 1e-06 
0.0 0.1451 0 2.0 1e-06 
0.0 0.1452 0 2.0 1e-06 
0.0 0.1453 0 2.0 1e-06 
0.0 0.1454 0 2.0 1e-06 
0.0 0.1455 0 2.0 1e-06 
0.0 0.1456 0 2.0 1e-06 
0.0 0.1457 0 2.0 1e-06 
0.0 0.1458 0 2.0 1e-06 
0.0 0.1459 0 2.0 1e-06 
0.0 0.146 0 2.0 1e-06 
0.0 0.1461 0 2.0 1e-06 
0.0 0.1462 0 2.0 1e-06 
0.0 0.1463 0 2.0 1e-06 
0.0 0.1464 0 2.0 1e-06 
0.0 0.1465 0 2.0 1e-06 
0.0 0.1466 0 2.0 1e-06 
0.0 0.1467 0 2.0 1e-06 
0.0 0.1468 0 2.0 1e-06 
0.0 0.1469 0 2.0 1e-06 
0.0 0.147 0 2.0 1e-06 
0.0 0.1471 0 2.0 1e-06 
0.0 0.1472 0 2.0 1e-06 
0.0 0.1473 0 2.0 1e-06 
0.0 0.1474 0 2.0 1e-06 
0.0 0.1475 0 2.0 1e-06 
0.0 0.1476 0 2.0 1e-06 
0.0 0.1477 0 2.0 1e-06 
0.0 0.1478 0 2.0 1e-06 
0.0 0.1479 0 2.0 1e-06 
0.0 0.148 0 2.0 1e-06 
0.0 0.1481 0 2.0 1e-06 
0.0 0.1482 0 2.0 1e-06 
0.0 0.1483 0 2.0 1e-06 
0.0 0.1484 0 2.0 1e-06 
0.0 0.1485 0 2.0 1e-06 
0.0 0.1486 0 2.0 1e-06 
0.0 0.1487 0 2.0 1e-06 
0.0 0.1488 0 2.0 1e-06 
0.0 0.1489 0 2.0 1e-06 
0.0 0.149 0 2.0 1e-06 
0.0 0.1491 0 2.0 1e-06 
0.0 0.1492 0 2.0 1e-06 
0.0 0.1493 0 2.0 1e-06 
0.0 0.1494 0 2.0 1e-06 
0.0 0.1495 0 2.0 1e-06 
0.0 0.1496 0 2.0 1e-06 
0.0 0.1497 0 2.0 1e-06 
0.0 0.1498 0 2.0 1e-06 
0.0 0.1499 0 2.0 1e-06 
0.0 0.15 0 2.0 1e-06 
0.0 0.1501 0 2.0 1e-06 
0.0 0.1502 0 2.0 1e-06 
0.0 0.1503 0 2.0 1e-06 
0.0 0.1504 0 2.0 1e-06 
0.0 0.1505 0 2.0 1e-06 
0.0 0.1506 0 2.0 1e-06 
0.0 0.1507 0 2.0 1e-06 
0.0 0.1508 0 2.0 1e-06 
0.0 0.1509 0 2.0 1e-06 
0.0 0.151 0 2.0 1e-06 
0.0 0.1511 0 2.0 1e-06 
0.0 0.1512 0 2.0 1e-06 
0.0 0.1513 0 2.0 1e-06 
0.0 0.1514 0 2.0 1e-06 
0.0 0.1515 0 2.0 1e-06 
0.0 0.1516 0 2.0 1e-06 
0.0 0.1517 0 2.0 1e-06 
0.0 0.1518 0 2.0 1e-06 
0.0 0.1519 0 2.0 1e-06 
0.0 0.152 0 2.0 1e-06 
0.0 0.1521 0 2.0 1e-06 
0.0 0.1522 0 2.0 1e-06 
0.0 0.1523 0 2.0 1e-06 
0.0 0.1524 0 2.0 1e-06 
0.0 0.1525 0 2.0 1e-06 
0.0 0.1526 0 2.0 1e-06 
0.0 0.1527 0 2.0 1e-06 
0.0 0.1528 0 2.0 1e-06 
0.0 0.1529 0 2.0 1e-06 
0.0 0.153 0 2.0 1e-06 
0.0 0.1531 0 2.0 1e-06 
0.0 0.1532 0 2.0 1e-06 
0.0 0.1533 0 2.0 1e-06 
0.0 0.1534 0 2.0 1e-06 
0.0 0.1535 0 2.0 1e-06 
0.0 0.1536 0 2.0 1e-06 
0.0 0.1537 0 2.0 1e-06 
0.0 0.1538 0 2.0 1e-06 
0.0 0.1539 0 2.0 1e-06 
0.0 0.154 0 2.0 1e-06 
0.0 0.1541 0 2.0 1e-06 
0.0 0.1542 0 2.0 1e-06 
0.0 0.1543 0 2.0 1e-06 
0.0 0.1544 0 2.0 1e-06 
0.0 0.1545 0 2.0 1e-06 
0.0 0.1546 0 2.0 1e-06 
0.0 0.1547 0 2.0 1e-06 
0.0 0.1548 0 2.0 1e-06 
0.0 0.1549 0 2.0 1e-06 
0.0 0.155 0 2.0 1e-06 
0.0 0.1551 0 2.0 1e-06 
0.0 0.1552 0 2.0 1e-06 
0.0 0.1553 0 2.0 1e-06 
0.0 0.1554 0 2.0 1e-06 
0.0 0.1555 0 2.0 1e-06 
0.0 0.1556 0 2.0 1e-06 
0.0 0.1557 0 2.0 1e-06 
0.0 0.1558 0 2.0 1e-06 
0.0 0.1559 0 2.0 1e-06 
0.0 0.156 0 2.0 1e-06 
0.0 0.1561 0 2.0 1e-06 
0.0 0.1562 0 2.0 1e-06 
0.0 0.1563 0 2.0 1e-06 
0.0 0.1564 0 2.0 1e-06 
0.0 0.1565 0 2.0 1e-06 
0.0 0.1566 0 2.0 1e-06 
0.0 0.1567 0 2.0 1e-06 
0.0 0.1568 0 2.0 1e-06 
0.0 0.1569 0 2.0 1e-06 
0.0 0.157 0 2.0 1e-06 
0.0 0.1571 0 2.0 1e-06 
0.0 0.1572 0 2.0 1e-06 
0.0 0.1573 0 2.0 1e-06 
0.0 0.1574 0 2.0 1e-06 
0.0 0.1575 0 2.0 1e-06 
0.0 0.1576 0 2.0 1e-06 
0.0 0.1577 0 2.0 1e-06 
0.0 0.1578 0 2.0 1e-06 
0.0 0.1579 0 2.0 1e-06 
0.0 0.158 0 2.0 1e-06 
0.0 0.1581 0 2.0 1e-06 
0.0 0.1582 0 2.0 1e-06 
0.0 0.1583 0 2.0 1e-06 
0.0 0.1584 0 2.0 1e-06 
0.0 0.1585 0 2.0 1e-06 
0.0 0.1586 0 2.0 1e-06 
0.0 0.1587 0 2.0 1e-06 
0.0 0.1588 0 2.0 1e-06 
0.0 0.1589 0 2.0 1e-06 
0.0 0.159 0 2.0 1e-06 
0.0 0.1591 0 2.0 1e-06 
0.0 0.1592 0 2.0 1e-06 
0.0 0.1593 0 2.0 1e-06 
0.0 0.1594 0 2.0 1e-06 
0.0 0.1595 0 2.0 1e-06 
0.0 0.1596 0 2.0 1e-06 
0.0 0.1597 0 2.0 1e-06 
0.0 0.1598 0 2.0 1e-06 
0.0 0.1599 0 2.0 1e-06 
0.0 0.16 0 2.0 1e-06 
0.0 0.1601 0 2.0 1e-06 
0.0 0.1602 0 2.0 1e-06 
0.0 0.1603 0 2.0 1e-06 
0.0 0.1604 0 2.0 1e-06 
0.0 0.1605 0 2.0 1e-06 
0.0 0.1606 0 2.0 1e-06 
0.0 0.1607 0 2.0 1e-06 
0.0 0.1608 0 2.0 1e-06 
0.0 0.1609 0 2.0 1e-06 
0.0 0.161 0 2.0 1e-06 
0.0 0.1611 0 2.0 1e-06 
0.0 0.1612 0 2.0 1e-06 
0.0 0.1613 0 2.0 1e-06 
0.0 0.1614 0 2.0 1e-06 
0.0 0.1615 0 2.0 1e-06 
0.0 0.1616 0 2.0 1e-06 
0.0 0.1617 0 2.0 1e-06 
0.0 0.1618 0 2.0 1e-06 
0.0 0.1619 0 2.0 1e-06 
0.0 0.162 0 2.0 1e-06 
0.0 0.1621 0 2.0 1e-06 
0.0 0.1622 0 2.0 1e-06 
0.0 0.1623 0 2.0 1e-06 
0.0 0.1624 0 2.0 1e-06 
0.0 0.1625 0 2.0 1e-06 
0.0 0.1626 0 2.0 1e-06 
0.0 0.1627 0 2.0 1e-06 
0.0 0.1628 0 2.0 1e-06 
0.0 0.1629 0 2.0 1e-06 
0.0 0.163 0 2.0 1e-06 
0.0 0.1631 0 2.0 1e-06 
0.0 0.1632 0 2.0 1e-06 
0.0 0.1633 0 2.0 1e-06 
0.0 0.1634 0 2.0 1e-06 
0.0 0.1635 0 2.0 1e-06 
0.0 0.1636 0 2.0 1e-06 
0.0 0.1637 0 2.0 1e-06 
0.0 0.1638 0 2.0 1e-06 
0.0 0.1639 0 2.0 1e-06 
0.0 0.164 0 2.0 1e-06 
0.0 0.1641 0 2.0 1e-06 
0.0 0.1642 0 2.0 1e-06 
0.0 0.1643 0 2.0 1e-06 
0.0 0.1644 0 2.0 1e-06 
0.0 0.1645 0 2.0 1e-06 
0.0 0.1646 0 2.0 1e-06 
0.0 0.1647 0 2.0 1e-06 
0.0 0.1648 0 2.0 1e-06 
0.0 0.1649 0 2.0 1e-06 
0.0 0.165 0 2.0 1e-06 
0.0 0.1651 0 2.0 1e-06 
0.0 0.1652 0 2.0 1e-06 
0.0 0.1653 0 2.0 1e-06 
0.0 0.1654 0 2.0 1e-06 
0.0 0.1655 0 2.0 1e-06 
0.0 0.1656 0 2.0 1e-06 
0.0 0.1657 0 2.0 1e-06 
0.0 0.1658 0 2.0 1e-06 
0.0 0.1659 0 2.0 1e-06 
0.0 0.166 0 2.0 1e-06 
0.0 0.1661 0 2.0 1e-06 
0.0 0.1662 0 2.0 1e-06 
0.0 0.1663 0 2.0 1e-06 
0.0 0.1664 0 2.0 1e-06 
0.0 0.1665 0 2.0 1e-06 
0.0 0.1666 0 2.0 1e-06 
0.0 0.1667 0 2.0 1e-06 
0.0 0.1668 0 2.0 1e-06 
0.0 0.1669 0 2.0 1e-06 
0.0 0.167 0 2.0 1e-06 
0.0 0.1671 0 2.0 1e-06 
0.0 0.1672 0 2.0 1e-06 
0.0 0.1673 0 2.0 1e-06 
0.0 0.1674 0 2.0 1e-06 
0.0 0.1675 0 2.0 1e-06 
0.0 0.1676 0 2.0 1e-06 
0.0 0.1677 0 2.0 1e-06 
0.0 0.1678 0 2.0 1e-06 
0.0 0.1679 0 2.0 1e-06 
0.0 0.168 0 2.0 1e-06 
0.0 0.1681 0 2.0 1e-06 
0.0 0.1682 0 2.0 1e-06 
0.0 0.1683 0 2.0 1e-06 
0.0 0.1684 0 2.0 1e-06 
0.0 0.1685 0 2.0 1e-06 
0.0 0.1686 0 2.0 1e-06 
0.0 0.1687 0 2.0 1e-06 
0.0 0.1688 0 2.0 1e-06 
0.0 0.1689 0 2.0 1e-06 
0.0 0.169 0 2.0 1e-06 
0.0 0.1691 0 2.0 1e-06 
0.0 0.1692 0 2.0 1e-06 
0.0 0.1693 0 2.0 1e-06 
0.0 0.1694 0 2.0 1e-06 
0.0 0.1695 0 2.0 1e-06 
0.0 0.1696 0 2.0 1e-06 
0.0 0.1697 0 2.0 1e-06 
0.0 0.1698 0 2.0 1e-06 
0.0 0.1699 0 2.0 1e-06 
0.0 0.17 0 2.0 1e-06 
0.0 0.1701 0 2.0 1e-06 
0.0 0.1702 0 2.0 1e-06 
0.0 0.1703 0 2.0 1e-06 
0.0 0.1704 0 2.0 1e-06 
0.0 0.1705 0 2.0 1e-06 
0.0 0.1706 0 2.0 1e-06 
0.0 0.1707 0 2.0 1e-06 
0.0 0.1708 0 2.0 1e-06 
0.0 0.1709 0 2.0 1e-06 
0.0 0.171 0 2.0 1e-06 
0.0 0.1711 0 2.0 1e-06 
0.0 0.1712 0 2.0 1e-06 
0.0 0.1713 0 2.0 1e-06 
0.0 0.1714 0 2.0 1e-06 
0.0 0.1715 0 2.0 1e-06 
0.0 0.1716 0 2.0 1e-06 
0.0 0.1717 0 2.0 1e-06 
0.0 0.1718 0 2.0 1e-06 
0.0 0.1719 0 2.0 1e-06 
0.0 0.172 0 2.0 1e-06 
0.0 0.1721 0 2.0 1e-06 
0.0 0.1722 0 2.0 1e-06 
0.0 0.1723 0 2.0 1e-06 
0.0 0.1724 0 2.0 1e-06 
0.0 0.1725 0 2.0 1e-06 
0.0 0.1726 0 2.0 1e-06 
0.0 0.1727 0 2.0 1e-06 
0.0 0.1728 0 2.0 1e-06 
0.0 0.1729 0 2.0 1e-06 
0.0 0.173 0 2.0 1e-06 
0.0 0.1731 0 2.0 1e-06 
0.0 0.1732 0 2.0 1e-06 
0.0 0.1733 0 2.0 1e-06 
0.0 0.1734 0 2.0 1e-06 
0.0 0.1735 0 2.0 1e-06 
0.0 0.1736 0 2.0 1e-06 
0.0 0.1737 0 2.0 1e-06 
0.0 0.1738 0 2.0 1e-06 
0.0 0.1739 0 2.0 1e-06 
0.0 0.174 0 2.0 1e-06 
0.0 0.1741 0 2.0 1e-06 
0.0 0.1742 0 2.0 1e-06 
0.0 0.1743 0 2.0 1e-06 
0.0 0.1744 0 2.0 1e-06 
0.0 0.1745 0 2.0 1e-06 
0.0 0.1746 0 2.0 1e-06 
0.0 0.1747 0 2.0 1e-06 
0.0 0.1748 0 2.0 1e-06 
0.0 0.1749 0 2.0 1e-06 
0.0 0.175 0 2.0 1e-06 
0.0 0.1751 0 2.0 1e-06 
0.0 0.1752 0 2.0 1e-06 
0.0 0.1753 0 2.0 1e-06 
0.0 0.1754 0 2.0 1e-06 
0.0 0.1755 0 2.0 1e-06 
0.0 0.1756 0 2.0 1e-06 
0.0 0.1757 0 2.0 1e-06 
0.0 0.1758 0 2.0 1e-06 
0.0 0.1759 0 2.0 1e-06 
0.0 0.176 0 2.0 1e-06 
0.0 0.1761 0 2.0 1e-06 
0.0 0.1762 0 2.0 1e-06 
0.0 0.1763 0 2.0 1e-06 
0.0 0.1764 0 2.0 1e-06 
0.0 0.1765 0 2.0 1e-06 
0.0 0.1766 0 2.0 1e-06 
0.0 0.1767 0 2.0 1e-06 
0.0 0.1768 0 2.0 1e-06 
0.0 0.1769 0 2.0 1e-06 
0.0 0.177 0 2.0 1e-06 
0.0 0.1771 0 2.0 1e-06 
0.0 0.1772 0 2.0 1e-06 
0.0 0.1773 0 2.0 1e-06 
0.0 0.1774 0 2.0 1e-06 
0.0 0.1775 0 2.0 1e-06 
0.0 0.1776 0 2.0 1e-06 
0.0 0.1777 0 2.0 1e-06 
0.0 0.1778 0 2.0 1e-06 
0.0 0.1779 0 2.0 1e-06 
0.0 0.178 0 2.0 1e-06 
0.0 0.1781 0 2.0 1e-06 
0.0 0.1782 0 2.0 1e-06 
0.0 0.1783 0 2.0 1e-06 
0.0 0.1784 0 2.0 1e-06 
0.0 0.1785 0 2.0 1e-06 
0.0 0.1786 0 2.0 1e-06 
0.0 0.1787 0 2.0 1e-06 
0.0 0.1788 0 2.0 1e-06 
0.0 0.1789 0 2.0 1e-06 
0.0 0.179 0 2.0 1e-06 
0.0 0.1791 0 2.0 1e-06 
0.0 0.1792 0 2.0 1e-06 
0.0 0.1793 0 2.0 1e-06 
0.0 0.1794 0 2.0 1e-06 
0.0 0.1795 0 2.0 1e-06 
0.0 0.1796 0 2.0 1e-06 
0.0 0.1797 0 2.0 1e-06 
0.0 0.1798 0 2.0 1e-06 
0.0 0.1799 0 2.0 1e-06 
0.0 0.18 0 2.0 1e-06 
0.0 0.1801 0 2.0 1e-06 
0.0 0.1802 0 2.0 1e-06 
0.0 0.1803 0 2.0 1e-06 
0.0 0.1804 0 2.0 1e-06 
0.0 0.1805 0 2.0 1e-06 
0.0 0.1806 0 2.0 1e-06 
0.0 0.1807 0 2.0 1e-06 
0.0 0.1808 0 2.0 1e-06 
0.0 0.1809 0 2.0 1e-06 
0.0 0.181 0 2.0 1e-06 
0.0 0.1811 0 2.0 1e-06 
0.0 0.1812 0 2.0 1e-06 
0.0 0.1813 0 2.0 1e-06 
0.0 0.1814 0 2.0 1e-06 
0.0 0.1815 0 2.0 1e-06 
0.0 0.1816 0 2.0 1e-06 
0.0 0.1817 0 2.0 1e-06 
0.0 0.1818 0 2.0 1e-06 
0.0 0.1819 0 2.0 1e-06 
0.0 0.182 0 2.0 1e-06 
0.0 0.1821 0 2.0 1e-06 
0.0 0.1822 0 2.0 1e-06 
0.0 0.1823 0 2.0 1e-06 
0.0 0.1824 0 2.0 1e-06 
0.0 0.1825 0 2.0 1e-06 
0.0 0.1826 0 2.0 1e-06 
0.0 0.1827 0 2.0 1e-06 
0.0 0.1828 0 2.0 1e-06 
0.0 0.1829 0 2.0 1e-06 
0.0 0.183 0 2.0 1e-06 
0.0 0.1831 0 2.0 1e-06 
0.0 0.1832 0 2.0 1e-06 
0.0 0.1833 0 2.0 1e-06 
0.0 0.1834 0 2.0 1e-06 
0.0 0.1835 0 2.0 1e-06 
0.0 0.1836 0 2.0 1e-06 
0.0 0.1837 0 2.0 1e-06 
0.0 0.1838 0 2.0 1e-06 
0.0 0.1839 0 2.0 1e-06 
0.0 0.184 0 2.0 1e-06 
0.0 0.1841 0 2.0 1e-06 
0.0 0.1842 0 2.0 1e-06 
0.0 0.1843 0 2.0 1e-06 
0.0 0.1844 0 2.0 1e-06 
0.0 0.1845 0 2.0 1e-06 
0.0 0.1846 0 2.0 1e-06 
0.0 0.1847 0 2.0 1e-06 
0.0 0.1848 0 2.0 1e-06 
0.0 0.1849 0 2.0 1e-06 
0.0 0.185 0 2.0 1e-06 
0.0 0.1851 0 2.0 1e-06 
0.0 0.1852 0 2.0 1e-06 
0.0 0.1853 0 2.0 1e-06 
0.0 0.1854 0 2.0 1e-06 
0.0 0.1855 0 2.0 1e-06 
0.0 0.1856 0 2.0 1e-06 
0.0 0.1857 0 2.0 1e-06 
0.0 0.1858 0 2.0 1e-06 
0.0 0.1859 0 2.0 1e-06 
0.0 0.186 0 2.0 1e-06 
0.0 0.1861 0 2.0 1e-06 
0.0 0.1862 0 2.0 1e-06 
0.0 0.1863 0 2.0 1e-06 
0.0 0.1864 0 2.0 1e-06 
0.0 0.1865 0 2.0 1e-06 
0.0 0.1866 0 2.0 1e-06 
0.0 0.1867 0 2.0 1e-06 
0.0 0.1868 0 2.0 1e-06 
0.0 0.1869 0 2.0 1e-06 
0.0 0.187 0 2.0 1e-06 
0.0 0.1871 0 2.0 1e-06 
0.0 0.1872 0 2.0 1e-06 
0.0 0.1873 0 2.0 1e-06 
0.0 0.1874 0 2.0 1e-06 
0.0 0.1875 0 2.0 1e-06 
0.0 0.1876 0 2.0 1e-06 
0.0 0.1877 0 2.0 1e-06 
0.0 0.1878 0 2.0 1e-06 
0.0 0.1879 0 2.0 1e-06 
0.0 0.188 0 2.0 1e-06 
0.0 0.1881 0 2.0 1e-06 
0.0 0.1882 0 2.0 1e-06 
0.0 0.1883 0 2.0 1e-06 
0.0 0.1884 0 2.0 1e-06 
0.0 0.1885 0 2.0 1e-06 
0.0 0.1886 0 2.0 1e-06 
0.0 0.1887 0 2.0 1e-06 
0.0 0.1888 0 2.0 1e-06 
0.0 0.1889 0 2.0 1e-06 
0.0 0.189 0 2.0 1e-06 
0.0 0.1891 0 2.0 1e-06 
0.0 0.1892 0 2.0 1e-06 
0.0 0.1893 0 2.0 1e-06 
0.0 0.1894 0 2.0 1e-06 
0.0 0.1895 0 2.0 1e-06 
0.0 0.1896 0 2.0 1e-06 
0.0 0.1897 0 2.0 1e-06 
0.0 0.1898 0 2.0 1e-06 
0.0 0.1899 0 2.0 1e-06 
0.0 0.19 0 2.0 1e-06 
0.0 0.1901 0 2.0 1e-06 
0.0 0.1902 0 2.0 1e-06 
0.0 0.1903 0 2.0 1e-06 
0.0 0.1904 0 2.0 1e-06 
0.0 0.1905 0 2.0 1e-06 
0.0 0.1906 0 2.0 1e-06 
0.0 0.1907 0 2.0 1e-06 
0.0 0.1908 0 2.0 1e-06 
0.0 0.1909 0 2.0 1e-06 
0.0 0.191 0 2.0 1e-06 
0.0 0.1911 0 2.0 1e-06 
0.0 0.1912 0 2.0 1e-06 
0.0 0.1913 0 2.0 1e-06 
0.0 0.1914 0 2.0 1e-06 
0.0 0.1915 0 2.0 1e-06 
0.0 0.1916 0 2.0 1e-06 
0.0 0.1917 0 2.0 1e-06 
0.0 0.1918 0 2.0 1e-06 
0.0 0.1919 0 2.0 1e-06 
0.0 0.192 0 2.0 1e-06 
0.0 0.1921 0 2.0 1e-06 
0.0 0.1922 0 2.0 1e-06 
0.0 0.1923 0 2.0 1e-06 
0.0 0.1924 0 2.0 1e-06 
0.0 0.1925 0 2.0 1e-06 
0.0 0.1926 0 2.0 1e-06 
0.0 0.1927 0 2.0 1e-06 
0.0 0.1928 0 2.0 1e-06 
0.0 0.1929 0 2.0 1e-06 
0.0 0.193 0 2.0 1e-06 
0.0 0.1931 0 2.0 1e-06 
0.0 0.1932 0 2.0 1e-06 
0.0 0.1933 0 2.0 1e-06 
0.0 0.1934 0 2.0 1e-06 
0.0 0.1935 0 2.0 1e-06 
0.0 0.1936 0 2.0 1e-06 
0.0 0.1937 0 2.0 1e-06 
0.0 0.1938 0 2.0 1e-06 
0.0 0.1939 0 2.0 1e-06 
0.0 0.194 0 2.0 1e-06 
0.0 0.1941 0 2.0 1e-06 
0.0 0.1942 0 2.0 1e-06 
0.0 0.1943 0 2.0 1e-06 
0.0 0.1944 0 2.0 1e-06 
0.0 0.1945 0 2.0 1e-06 
0.0 0.1946 0 2.0 1e-06 
0.0 0.1947 0 2.0 1e-06 
0.0 0.1948 0 2.0 1e-06 
0.0 0.1949 0 2.0 1e-06 
0.0 0.195 0 2.0 1e-06 
0.0 0.1951 0 2.0 1e-06 
0.0 0.1952 0 2.0 1e-06 
0.0 0.1953 0 2.0 1e-06 
0.0 0.1954 0 2.0 1e-06 
0.0 0.1955 0 2.0 1e-06 
0.0 0.1956 0 2.0 1e-06 
0.0 0.1957 0 2.0 1e-06 
0.0 0.1958 0 2.0 1e-06 
0.0 0.1959 0 2.0 1e-06 
0.0 0.196 0 2.0 1e-06 
0.0 0.1961 0 2.0 1e-06 
0.0 0.1962 0 2.0 1e-06 
0.0 0.1963 0 2.0 1e-06 
0.0 0.1964 0 2.0 1e-06 
0.0 0.1965 0 2.0 1e-06 
0.0 0.1966 0 2.0 1e-06 
0.0 0.1967 0 2.0 1e-06 
0.0 0.1968 0 2.0 1e-06 
0.0 0.1969 0 2.0 1e-06 
0.0 0.197 0 2.0 1e-06 
0.0 0.1971 0 2.0 1e-06 
0.0 0.1972 0 2.0 1e-06 
0.0 0.1973 0 2.0 1e-06 
0.0 0.1974 0 2.0 1e-06 
0.0 0.1975 0 2.0 1e-06 
0.0 0.1976 0 2.0 1e-06 
0.0 0.1977 0 2.0 1e-06 
0.0 0.1978 0 2.0 1e-06 
0.0 0.1979 0 2.0 1e-06 
0.0 0.198 0 2.0 1e-06 
0.0 0.1981 0 2.0 1e-06 
0.0 0.1982 0 2.0 1e-06 
0.0 0.1983 0 2.0 1e-06 
0.0 0.1984 0 2.0 1e-06 
0.0 0.1985 0 2.0 1e-06 
0.0 0.1986 0 2.0 1e-06 
0.0 0.1987 0 2.0 1e-06 
0.0 0.1988 0 2.0 1e-06 
0.0 0.1989 0 2.0 1e-06 
0.0 0.199 0 2.0 1e-06 
0.0 0.1991 0 2.0 1e-06 
0.0 0.1992 0 2.0 1e-06 
0.0 0.1993 0 2.0 1e-06 
0.0 0.1994 0 2.0 1e-06 
0.0 0.1995 0 2.0 1e-06 
0.0 0.1996 0 2.0 1e-06 
0.0 0.1997 0 2.0 1e-06 
0.0 0.1998 0 2.0 1e-06 
0.0 0.1999 0 2.0 1e-06 
0.0 0.2 0 2.0 1e-06 
0.0 0.2001 0 2.0 1e-06 
0.0 0.2002 0 2.0 1e-06 
0.0 0.2003 0 2.0 1e-06 
0.0 0.2004 0 2.0 1e-06 
0.0 0.2005 0 2.0 1e-06 
0.0 0.2006 0 2.0 1e-06 
0.0 0.2007 0 2.0 1e-06 
0.0 0.2008 0 2.0 1e-06 
0.0 0.2009 0 2.0 1e-06 
0.0 0.201 0 2.0 1e-06 
0.0 0.2011 0 2.0 1e-06 
0.0 0.2012 0 2.0 1e-06 
0.0 0.2013 0 2.0 1e-06 
0.0 0.2014 0 2.0 1e-06 
0.0 0.2015 0 2.0 1e-06 
0.0 0.2016 0 2.0 1e-06 
0.0 0.2017 0 2.0 1e-06 
0.0 0.2018 0 2.0 1e-06 
0.0 0.2019 0 2.0 1e-06 
0.0 0.202 0 2.0 1e-06 
0.0 0.2021 0 2.0 1e-06 
0.0 0.2022 0 2.0 1e-06 
0.0 0.2023 0 2.0 1e-06 
0.0 0.2024 0 2.0 1e-06 
0.0 0.2025 0 2.0 1e-06 
0.0 0.2026 0 2.0 1e-06 
0.0 0.2027 0 2.0 1e-06 
0.0 0.2028 0 2.0 1e-06 
0.0 0.2029 0 2.0 1e-06 
0.0 0.203 0 2.0 1e-06 
0.0 0.2031 0 2.0 1e-06 
0.0 0.2032 0 2.0 1e-06 
0.0 0.2033 0 2.0 1e-06 
0.0 0.2034 0 2.0 1e-06 
0.0 0.2035 0 2.0 1e-06 
0.0 0.2036 0 2.0 1e-06 
0.0 0.2037 0 2.0 1e-06 
0.0 0.2038 0 2.0 1e-06 
0.0 0.2039 0 2.0 1e-06 
0.0 0.204 0 2.0 1e-06 
0.0 0.2041 0 2.0 1e-06 
0.0 0.2042 0 2.0 1e-06 
0.0 0.2043 0 2.0 1e-06 
0.0 0.2044 0 2.0 1e-06 
0.0 0.2045 0 2.0 1e-06 
0.0 0.2046 0 2.0 1e-06 
0.0 0.2047 0 2.0 1e-06 
0.0 0.2048 0 2.0 1e-06 
0.0 0.2049 0 2.0 1e-06 
0.0 0.205 0 2.0 1e-06 
0.0 0.2051 0 2.0 1e-06 
0.0 0.2052 0 2.0 1e-06 
0.0 0.2053 0 2.0 1e-06 
0.0 0.2054 0 2.0 1e-06 
0.0 0.2055 0 2.0 1e-06 
0.0 0.2056 0 2.0 1e-06 
0.0 0.2057 0 2.0 1e-06 
0.0 0.2058 0 2.0 1e-06 
0.0 0.2059 0 2.0 1e-06 
0.0 0.206 0 2.0 1e-06 
0.0 0.2061 0 2.0 1e-06 
0.0 0.2062 0 2.0 1e-06 
0.0 0.2063 0 2.0 1e-06 
0.0 0.2064 0 2.0 1e-06 
0.0 0.2065 0 2.0 1e-06 
0.0 0.2066 0 2.0 1e-06 
0.0 0.2067 0 2.0 1e-06 
0.0 0.2068 0 2.0 1e-06 
0.0 0.2069 0 2.0 1e-06 
0.0 0.207 0 2.0 1e-06 
0.0 0.2071 0 2.0 1e-06 
0.0 0.2072 0 2.0 1e-06 
0.0 0.2073 0 2.0 1e-06 
0.0 0.2074 0 2.0 1e-06 
0.0 0.2075 0 2.0 1e-06 
0.0 0.2076 0 2.0 1e-06 
0.0 0.2077 0 2.0 1e-06 
0.0 0.2078 0 2.0 1e-06 
0.0 0.2079 0 2.0 1e-06 
0.0 0.208 0 2.0 1e-06 
0.0 0.2081 0 2.0 1e-06 
0.0 0.2082 0 2.0 1e-06 
0.0 0.2083 0 2.0 1e-06 
0.0 0.2084 0 2.0 1e-06 
0.0 0.2085 0 2.0 1e-06 
0.0 0.2086 0 2.0 1e-06 
0.0 0.2087 0 2.0 1e-06 
0.0 0.2088 0 2.0 1e-06 
0.0 0.2089 0 2.0 1e-06 
0.0 0.209 0 2.0 1e-06 
0.0 0.2091 0 2.0 1e-06 
0.0 0.2092 0 2.0 1e-06 
0.0 0.2093 0 2.0 1e-06 
0.0 0.2094 0 2.0 1e-06 
0.0 0.2095 0 2.0 1e-06 
0.0 0.2096 0 2.0 1e-06 
0.0 0.2097 0 2.0 1e-06 
0.0 0.2098 0 2.0 1e-06 
0.0 0.2099 0 2.0 1e-06 
0.0 0.21 0 2.0 1e-06 
0.0 0.2101 0 2.0 1e-06 
0.0 0.2102 0 2.0 1e-06 
0.0 0.2103 0 2.0 1e-06 
0.0 0.2104 0 2.0 1e-06 
0.0 0.2105 0 2.0 1e-06 
0.0 0.2106 0 2.0 1e-06 
0.0 0.2107 0 2.0 1e-06 
0.0 0.2108 0 2.0 1e-06 
0.0 0.2109 0 2.0 1e-06 
0.0 0.211 0 2.0 1e-06 
0.0 0.2111 0 2.0 1e-06 
0.0 0.2112 0 2.0 1e-06 
0.0 0.2113 0 2.0 1e-06 
0.0 0.2114 0 2.0 1e-06 
0.0 0.2115 0 2.0 1e-06 
0.0 0.2116 0 2.0 1e-06 
0.0 0.2117 0 2.0 1e-06 
0.0 0.2118 0 2.0 1e-06 
0.0 0.2119 0 2.0 1e-06 
0.0 0.212 0 2.0 1e-06 
0.0 0.2121 0 2.0 1e-06 
0.0 0.2122 0 2.0 1e-06 
0.0 0.2123 0 2.0 1e-06 
0.0 0.2124 0 2.0 1e-06 
0.0 0.2125 0 2.0 1e-06 
0.0 0.2126 0 2.0 1e-06 
0.0 0.2127 0 2.0 1e-06 
0.0 0.2128 0 2.0 1e-06 
0.0 0.2129 0 2.0 1e-06 
0.0 0.213 0 2.0 1e-06 
0.0 0.2131 0 2.0 1e-06 
0.0 0.2132 0 2.0 1e-06 
0.0 0.2133 0 2.0 1e-06 
0.0 0.2134 0 2.0 1e-06 
0.0 0.2135 0 2.0 1e-06 
0.0 0.2136 0 2.0 1e-06 
0.0 0.2137 0 2.0 1e-06 
0.0 0.2138 0 2.0 1e-06 
0.0 0.2139 0 2.0 1e-06 
0.0 0.214 0 2.0 1e-06 
0.0 0.2141 0 2.0 1e-06 
0.0 0.2142 0 2.0 1e-06 
0.0 0.2143 0 2.0 1e-06 
0.0 0.2144 0 2.0 1e-06 
0.0 0.2145 0 2.0 1e-06 
0.0 0.2146 0 2.0 1e-06 
0.0 0.2147 0 2.0 1e-06 
0.0 0.2148 0 2.0 1e-06 
0.0 0.2149 0 2.0 1e-06 
0.0 0.215 0 2.0 1e-06 
0.0 0.2151 0 2.0 1e-06 
0.0 0.2152 0 2.0 1e-06 
0.0 0.2153 0 2.0 1e-06 
0.0 0.2154 0 2.0 1e-06 
0.0 0.2155 0 2.0 1e-06 
0.0 0.2156 0 2.0 1e-06 
0.0 0.2157 0 2.0 1e-06 
0.0 0.2158 0 2.0 1e-06 
0.0 0.2159 0 2.0 1e-06 
0.0 0.216 0 2.0 1e-06 
0.0 0.2161 0 2.0 1e-06 
0.0 0.2162 0 2.0 1e-06 
0.0 0.2163 0 2.0 1e-06 
0.0 0.2164 0 2.0 1e-06 
0.0 0.2165 0 2.0 1e-06 
0.0 0.2166 0 2.0 1e-06 
0.0 0.2167 0 2.0 1e-06 
0.0 0.2168 0 2.0 1e-06 
0.0 0.2169 0 2.0 1e-06 
0.0 0.217 0 2.0 1e-06 
0.0 0.2171 0 2.0 1e-06 
0.0 0.2172 0 2.0 1e-06 
0.0 0.2173 0 2.0 1e-06 
0.0 0.2174 0 2.0 1e-06 
0.0 0.2175 0 2.0 1e-06 
0.0 0.2176 0 2.0 1e-06 
0.0 0.2177 0 2.0 1e-06 
0.0 0.2178 0 2.0 1e-06 
0.0 0.2179 0 2.0 1e-06 
0.0 0.218 0 2.0 1e-06 
0.0 0.2181 0 2.0 1e-06 
0.0 0.2182 0 2.0 1e-06 
0.0 0.2183 0 2.0 1e-06 
0.0 0.2184 0 2.0 1e-06 
0.0 0.2185 0 2.0 1e-06 
0.0 0.2186 0 2.0 1e-06 
0.0 0.2187 0 2.0 1e-06 
0.0 0.2188 0 2.0 1e-06 
0.0 0.2189 0 2.0 1e-06 
0.0 0.219 0 2.0 1e-06 
0.0 0.2191 0 2.0 1e-06 
0.0 0.2192 0 2.0 1e-06 
0.0 0.2193 0 2.0 1e-06 
0.0 0.2194 0 2.0 1e-06 
0.0 0.2195 0 2.0 1e-06 
0.0 0.2196 0 2.0 1e-06 
0.0 0.2197 0 2.0 1e-06 
0.0 0.2198 0 2.0 1e-06 
0.0 0.2199 0 2.0 1e-06 
0.0 0.22 0 2.0 1e-06 
0.0 0.2201 0 2.0 1e-06 
0.0 0.2202 0 2.0 1e-06 
0.0 0.2203 0 2.0 1e-06 
0.0 0.2204 0 2.0 1e-06 
0.0 0.2205 0 2.0 1e-06 
0.0 0.2206 0 2.0 1e-06 
0.0 0.2207 0 2.0 1e-06 
0.0 0.2208 0 2.0 1e-06 
0.0 0.2209 0 2.0 1e-06 
0.0 0.221 0 2.0 1e-06 
0.0 0.2211 0 2.0 1e-06 
0.0 0.2212 0 2.0 1e-06 
0.0 0.2213 0 2.0 1e-06 
0.0 0.2214 0 2.0 1e-06 
0.0 0.2215 0 2.0 1e-06 
0.0 0.2216 0 2.0 1e-06 
0.0 0.2217 0 2.0 1e-06 
0.0 0.2218 0 2.0 1e-06 
0.0 0.2219 0 2.0 1e-06 
0.0 0.222 0 2.0 1e-06 
0.0 0.2221 0 2.0 1e-06 
0.0 0.2222 0 2.0 1e-06 
0.0 0.2223 0 2.0 1e-06 
0.0 0.2224 0 2.0 1e-06 
0.0 0.2225 0 2.0 1e-06 
0.0 0.2226 0 2.0 1e-06 
0.0 0.2227 0 2.0 1e-06 
0.0 0.2228 0 2.0 1e-06 
0.0 0.2229 0 2.0 1e-06 
0.0 0.223 0 2.0 1e-06 
0.0 0.2231 0 2.0 1e-06 
0.0 0.2232 0 2.0 1e-06 
0.0 0.2233 0 2.0 1e-06 
0.0 0.2234 0 2.0 1e-06 
0.0 0.2235 0 2.0 1e-06 
0.0 0.2236 0 2.0 1e-06 
0.0 0.2237 0 2.0 1e-06 
0.0 0.2238 0 2.0 1e-06 
0.0 0.2239 0 2.0 1e-06 
0.0 0.224 0 2.0 1e-06 
0.0 0.2241 0 2.0 1e-06 
0.0 0.2242 0 2.0 1e-06 
0.0 0.2243 0 2.0 1e-06 
0.0 0.2244 0 2.0 1e-06 
0.0 0.2245 0 2.0 1e-06 
0.0 0.2246 0 2.0 1e-06 
0.0 0.2247 0 2.0 1e-06 
0.0 0.2248 0 2.0 1e-06 
0.0 0.2249 0 2.0 1e-06 
0.0 0.225 0 2.0 1e-06 
0.0 0.2251 0 2.0 1e-06 
0.0 0.2252 0 2.0 1e-06 
0.0 0.2253 0 2.0 1e-06 
0.0 0.2254 0 2.0 1e-06 
0.0 0.2255 0 2.0 1e-06 
0.0 0.2256 0 2.0 1e-06 
0.0 0.2257 0 2.0 1e-06 
0.0 0.2258 0 2.0 1e-06 
0.0 0.2259 0 2.0 1e-06 
0.0 0.226 0 2.0 1e-06 
0.0 0.2261 0 2.0 1e-06 
0.0 0.2262 0 2.0 1e-06 
0.0 0.2263 0 2.0 1e-06 
0.0 0.2264 0 2.0 1e-06 
0.0 0.2265 0 2.0 1e-06 
0.0 0.2266 0 2.0 1e-06 
0.0 0.2267 0 2.0 1e-06 
0.0 0.2268 0 2.0 1e-06 
0.0 0.2269 0 2.0 1e-06 
0.0 0.227 0 2.0 1e-06 
0.0 0.2271 0 2.0 1e-06 
0.0 0.2272 0 2.0 1e-06 
0.0 0.2273 0 2.0 1e-06 
0.0 0.2274 0 2.0 1e-06 
0.0 0.2275 0 2.0 1e-06 
0.0 0.2276 0 2.0 1e-06 
0.0 0.2277 0 2.0 1e-06 
0.0 0.2278 0 2.0 1e-06 
0.0 0.2279 0 2.0 1e-06 
0.0 0.228 0 2.0 1e-06 
0.0 0.2281 0 2.0 1e-06 
0.0 0.2282 0 2.0 1e-06 
0.0 0.2283 0 2.0 1e-06 
0.0 0.2284 0 2.0 1e-06 
0.0 0.2285 0 2.0 1e-06 
0.0 0.2286 0 2.0 1e-06 
0.0 0.2287 0 2.0 1e-06 
0.0 0.2288 0 2.0 1e-06 
0.0 0.2289 0 2.0 1e-06 
0.0 0.229 0 2.0 1e-06 
0.0 0.2291 0 2.0 1e-06 
0.0 0.2292 0 2.0 1e-06 
0.0 0.2293 0 2.0 1e-06 
0.0 0.2294 0 2.0 1e-06 
0.0 0.2295 0 2.0 1e-06 
0.0 0.2296 0 2.0 1e-06 
0.0 0.2297 0 2.0 1e-06 
0.0 0.2298 0 2.0 1e-06 
0.0 0.2299 0 2.0 1e-06 
0.0 0.23 0 2.0 1e-06 
0.0 0.2301 0 2.0 1e-06 
0.0 0.2302 0 2.0 1e-06 
0.0 0.2303 0 2.0 1e-06 
0.0 0.2304 0 2.0 1e-06 
0.0 0.2305 0 2.0 1e-06 
0.0 0.2306 0 2.0 1e-06 
0.0 0.2307 0 2.0 1e-06 
0.0 0.2308 0 2.0 1e-06 
0.0 0.2309 0 2.0 1e-06 
0.0 0.231 0 2.0 1e-06 
0.0 0.2311 0 2.0 1e-06 
0.0 0.2312 0 2.0 1e-06 
0.0 0.2313 0 2.0 1e-06 
0.0 0.2314 0 2.0 1e-06 
0.0 0.2315 0 2.0 1e-06 
0.0 0.2316 0 2.0 1e-06 
0.0 0.2317 0 2.0 1e-06 
0.0 0.2318 0 2.0 1e-06 
0.0 0.2319 0 2.0 1e-06 
0.0 0.232 0 2.0 1e-06 
0.0 0.2321 0 2.0 1e-06 
0.0 0.2322 0 2.0 1e-06 
0.0 0.2323 0 2.0 1e-06 
0.0 0.2324 0 2.0 1e-06 
0.0 0.2325 0 2.0 1e-06 
0.0 0.2326 0 2.0 1e-06 
0.0 0.2327 0 2.0 1e-06 
0.0 0.2328 0 2.0 1e-06 
0.0 0.2329 0 2.0 1e-06 
0.0 0.233 0 2.0 1e-06 
0.0 0.2331 0 2.0 1e-06 
0.0 0.2332 0 2.0 1e-06 
0.0 0.2333 0 2.0 1e-06 
0.0 0.2334 0 2.0 1e-06 
0.0 0.2335 0 2.0 1e-06 
0.0 0.2336 0 2.0 1e-06 
0.0 0.2337 0 2.0 1e-06 
0.0 0.2338 0 2.0 1e-06 
0.0 0.2339 0 2.0 1e-06 
0.0 0.234 0 2.0 1e-06 
0.0 0.2341 0 2.0 1e-06 
0.0 0.2342 0 2.0 1e-06 
0.0 0.2343 0 2.0 1e-06 
0.0 0.2344 0 2.0 1e-06 
0.0 0.2345 0 2.0 1e-06 
0.0 0.2346 0 2.0 1e-06 
0.0 0.2347 0 2.0 1e-06 
0.0 0.2348 0 2.0 1e-06 
0.0 0.2349 0 2.0 1e-06 
0.0 0.235 0 2.0 1e-06 
0.0 0.2351 0 2.0 1e-06 
0.0 0.2352 0 2.0 1e-06 
0.0 0.2353 0 2.0 1e-06 
0.0 0.2354 0 2.0 1e-06 
0.0 0.2355 0 2.0 1e-06 
0.0 0.2356 0 2.0 1e-06 
0.0 0.2357 0 2.0 1e-06 
0.0 0.2358 0 2.0 1e-06 
0.0 0.2359 0 2.0 1e-06 
0.0 0.236 0 2.0 1e-06 
0.0 0.2361 0 2.0 1e-06 
0.0 0.2362 0 2.0 1e-06 
0.0 0.2363 0 2.0 1e-06 
0.0 0.2364 0 2.0 1e-06 
0.0 0.2365 0 2.0 1e-06 
0.0 0.2366 0 2.0 1e-06 
0.0 0.2367 0 2.0 1e-06 
0.0 0.2368 0 2.0 1e-06 
0.0 0.2369 0 2.0 1e-06 
0.0 0.237 0 2.0 1e-06 
0.0 0.2371 0 2.0 1e-06 
0.0 0.2372 0 2.0 1e-06 
0.0 0.2373 0 2.0 1e-06 
0.0 0.2374 0 2.0 1e-06 
0.0 0.2375 0 2.0 1e-06 
0.0 0.2376 0 2.0 1e-06 
0.0 0.2377 0 2.0 1e-06 
0.0 0.2378 0 2.0 1e-06 
0.0 0.2379 0 2.0 1e-06 
0.0 0.238 0 2.0 1e-06 
0.0 0.2381 0 2.0 1e-06 
0.0 0.2382 0 2.0 1e-06 
0.0 0.2383 0 2.0 1e-06 
0.0 0.2384 0 2.0 1e-06 
0.0 0.2385 0 2.0 1e-06 
0.0 0.2386 0 2.0 1e-06 
0.0 0.2387 0 2.0 1e-06 
0.0 0.2388 0 2.0 1e-06 
0.0 0.2389 0 2.0 1e-06 
0.0 0.239 0 2.0 1e-06 
0.0 0.2391 0 2.0 1e-06 
0.0 0.2392 0 2.0 1e-06 
0.0 0.2393 0 2.0 1e-06 
0.0 0.2394 0 2.0 1e-06 
0.0 0.2395 0 2.0 1e-06 
0.0 0.2396 0 2.0 1e-06 
0.0 0.2397 0 2.0 1e-06 
0.0 0.2398 0 2.0 1e-06 
0.0 0.2399 0 2.0 1e-06 
0.0 0.24 0 2.0 1e-06 
0.0 0.2401 0 2.0 1e-06 
0.0 0.2402 0 2.0 1e-06 
0.0 0.2403 0 2.0 1e-06 
0.0 0.2404 0 2.0 1e-06 
0.0 0.2405 0 2.0 1e-06 
0.0 0.2406 0 2.0 1e-06 
0.0 0.2407 0 2.0 1e-06 
0.0 0.2408 0 2.0 1e-06 
0.0 0.2409 0 2.0 1e-06 
0.0 0.241 0 2.0 1e-06 
0.0 0.2411 0 2.0 1e-06 
0.0 0.2412 0 2.0 1e-06 
0.0 0.2413 0 2.0 1e-06 
0.0 0.2414 0 2.0 1e-06 
0.0 0.2415 0 2.0 1e-06 
0.0 0.2416 0 2.0 1e-06 
0.0 0.2417 0 2.0 1e-06 
0.0 0.2418 0 2.0 1e-06 
0.0 0.2419 0 2.0 1e-06 
0.0 0.242 0 2.0 1e-06 
0.0 0.2421 0 2.0 1e-06 
0.0 0.2422 0 2.0 1e-06 
0.0 0.2423 0 2.0 1e-06 
0.0 0.2424 0 2.0 1e-06 
0.0 0.2425 0 2.0 1e-06 
0.0 0.2426 0 2.0 1e-06 
0.0 0.2427 0 2.0 1e-06 
0.0 0.2428 0 2.0 1e-06 
0.0 0.2429 0 2.0 1e-06 
0.0 0.243 0 2.0 1e-06 
0.0 0.2431 0 2.0 1e-06 
0.0 0.2432 0 2.0 1e-06 
0.0 0.2433 0 2.0 1e-06 
0.0 0.2434 0 2.0 1e-06 
0.0 0.2435 0 2.0 1e-06 
0.0 0.2436 0 2.0 1e-06 
0.0 0.2437 0 2.0 1e-06 
0.0 0.2438 0 2.0 1e-06 
0.0 0.2439 0 2.0 1e-06 
0.0 0.244 0 2.0 1e-06 
0.0 0.2441 0 2.0 1e-06 
0.0 0.2442 0 2.0 1e-06 
0.0 0.2443 0 2.0 1e-06 
0.0 0.2444 0 2.0 1e-06 
0.0 0.2445 0 2.0 1e-06 
0.0 0.2446 0 2.0 1e-06 
0.0 0.2447 0 2.0 1e-06 
0.0 0.2448 0 2.0 1e-06 
0.0 0.2449 0 2.0 1e-06 
0.0 0.245 0 2.0 1e-06 
0.0 0.2451 0 2.0 1e-06 
0.0 0.2452 0 2.0 1e-06 
0.0 0.2453 0 2.0 1e-06 
0.0 0.2454 0 2.0 1e-06 
0.0 0.2455 0 2.0 1e-06 
0.0 0.2456 0 2.0 1e-06 
0.0 0.2457 0 2.0 1e-06 
0.0 0.2458 0 2.0 1e-06 
0.0 0.2459 0 2.0 1e-06 
0.0 0.246 0 2.0 1e-06 
0.0 0.2461 0 2.0 1e-06 
0.0 0.2462 0 2.0 1e-06 
0.0 0.2463 0 2.0 1e-06 
0.0 0.2464 0 2.0 1e-06 
0.0 0.2465 0 2.0 1e-06 
0.0 0.2466 0 2.0 1e-06 
0.0 0.2467 0 2.0 1e-06 
0.0 0.2468 0 2.0 1e-06 
0.0 0.2469 0 2.0 1e-06 
0.0 0.247 0 2.0 1e-06 
0.0 0.2471 0 2.0 1e-06 
0.0 0.2472 0 2.0 1e-06 
0.0 0.2473 0 2.0 1e-06 
0.0 0.2474 0 2.0 1e-06 
0.0 0.2475 0 2.0 1e-06 
0.0 0.2476 0 2.0 1e-06 
0.0 0.2477 0 2.0 1e-06 
0.0 0.2478 0 2.0 1e-06 
0.0 0.2479 0 2.0 1e-06 
0.0 0.248 0 2.0 1e-06 
0.0 0.2481 0 2.0 1e-06 
0.0 0.2482 0 2.0 1e-06 
0.0 0.2483 0 2.0 1e-06 
0.0 0.2484 0 2.0 1e-06 
0.0 0.2485 0 2.0 1e-06 
0.0 0.2486 0 2.0 1e-06 
0.0 0.2487 0 2.0 1e-06 
0.0 0.2488 0 2.0 1e-06 
0.0 0.2489 0 2.0 1e-06 
0.0 0.249 0 2.0 1e-06 
0.0 0.2491 0 2.0 1e-06 
0.0 0.2492 0 2.0 1e-06 
0.0 0.2493 0 2.0 1e-06 
0.0 0.2494 0 2.0 1e-06 
0.0 0.2495 0 2.0 1e-06 
0.0 0.2496 0 2.0 1e-06 
0.0 0.2497 0 2.0 1e-06 
0.0 0.2498 0 2.0 1e-06 
0.0 0.2499 0 2.0 1e-06 
0.0 0.25 0 2.0 1e-06 
0.0 0.2501 0 2.0 1e-06 
0.0 0.2502 0 2.0 1e-06 
0.0 0.2503 0 2.0 1e-06 
0.0 0.2504 0 2.0 1e-06 
0.0 0.2505 0 2.0 1e-06 
0.0 0.2506 0 2.0 1e-06 
0.0 0.2507 0 2.0 1e-06 
0.0 0.2508 0 2.0 1e-06 
0.0 0.2509 0 2.0 1e-06 
0.0 0.251 0 2.0 1e-06 
0.0 0.2511 0 2.0 1e-06 
0.0 0.2512 0 2.0 1e-06 
0.0 0.2513 0 2.0 1e-06 
0.0 0.2514 0 2.0 1e-06 
0.0 0.2515 0 2.0 1e-06 
0.0 0.2516 0 2.0 1e-06 
0.0 0.2517 0 2.0 1e-06 
0.0 0.2518 0 2.0 1e-06 
0.0 0.2519 0 2.0 1e-06 
0.0 0.252 0 2.0 1e-06 
0.0 0.2521 0 2.0 1e-06 
0.0 0.2522 0 2.0 1e-06 
0.0 0.2523 0 2.0 1e-06 
0.0 0.2524 0 2.0 1e-06 
0.0 0.2525 0 2.0 1e-06 
0.0 0.2526 0 2.0 1e-06 
0.0 0.2527 0 2.0 1e-06 
0.0 0.2528 0 2.0 1e-06 
0.0 0.2529 0 2.0 1e-06 
0.0 0.253 0 2.0 1e-06 
0.0 0.2531 0 2.0 1e-06 
0.0 0.2532 0 2.0 1e-06 
0.0 0.2533 0 2.0 1e-06 
0.0 0.2534 0 2.0 1e-06 
0.0 0.2535 0 2.0 1e-06 
0.0 0.2536 0 2.0 1e-06 
0.0 0.2537 0 2.0 1e-06 
0.0 0.2538 0 2.0 1e-06 
0.0 0.2539 0 2.0 1e-06 
0.0 0.254 0 2.0 1e-06 
0.0 0.2541 0 2.0 1e-06 
0.0 0.2542 0 2.0 1e-06 
0.0 0.2543 0 2.0 1e-06 
0.0 0.2544 0 2.0 1e-06 
0.0 0.2545 0 2.0 1e-06 
0.0 0.2546 0 2.0 1e-06 
0.0 0.2547 0 2.0 1e-06 
0.0 0.2548 0 2.0 1e-06 
0.0 0.2549 0 2.0 1e-06 
0.0 0.255 0 2.0 1e-06 
0.0 0.2551 0 2.0 1e-06 
0.0 0.2552 0 2.0 1e-06 
0.0 0.2553 0 2.0 1e-06 
0.0 0.2554 0 2.0 1e-06 
0.0 0.2555 0 2.0 1e-06 
0.0 0.2556 0 2.0 1e-06 
0.0 0.2557 0 2.0 1e-06 
0.0 0.2558 0 2.0 1e-06 
0.0 0.2559 0 2.0 1e-06 
0.0 0.256 0 2.0 1e-06 
0.0 0.2561 0 2.0 1e-06 
0.0 0.2562 0 2.0 1e-06 
0.0 0.2563 0 2.0 1e-06 
0.0 0.2564 0 2.0 1e-06 
0.0 0.2565 0 2.0 1e-06 
0.0 0.2566 0 2.0 1e-06 
0.0 0.2567 0 2.0 1e-06 
0.0 0.2568 0 2.0 1e-06 
0.0 0.2569 0 2.0 1e-06 
0.0 0.257 0 2.0 1e-06 
0.0 0.2571 0 2.0 1e-06 
0.0 0.2572 0 2.0 1e-06 
0.0 0.2573 0 2.0 1e-06 
0.0 0.2574 0 2.0 1e-06 
0.0 0.2575 0 2.0 1e-06 
0.0 0.2576 0 2.0 1e-06 
0.0 0.2577 0 2.0 1e-06 
0.0 0.2578 0 2.0 1e-06 
0.0 0.2579 0 2.0 1e-06 
0.0 0.258 0 2.0 1e-06 
0.0 0.2581 0 2.0 1e-06 
0.0 0.2582 0 2.0 1e-06 
0.0 0.2583 0 2.0 1e-06 
0.0 0.2584 0 2.0 1e-06 
0.0 0.2585 0 2.0 1e-06 
0.0 0.2586 0 2.0 1e-06 
0.0 0.2587 0 2.0 1e-06 
0.0 0.2588 0 2.0 1e-06 
0.0 0.2589 0 2.0 1e-06 
0.0 0.259 0 2.0 1e-06 
0.0 0.2591 0 2.0 1e-06 
0.0 0.2592 0 2.0 1e-06 
0.0 0.2593 0 2.0 1e-06 
0.0 0.2594 0 2.0 1e-06 
0.0 0.2595 0 2.0 1e-06 
0.0 0.2596 0 2.0 1e-06 
0.0 0.2597 0 2.0 1e-06 
0.0 0.2598 0 2.0 1e-06 
0.0 0.2599 0 2.0 1e-06 
0.0 0.26 0 2.0 1e-06 
0.0 0.2601 0 2.0 1e-06 
0.0 0.2602 0 2.0 1e-06 
0.0 0.2603 0 2.0 1e-06 
0.0 0.2604 0 2.0 1e-06 
0.0 0.2605 0 2.0 1e-06 
0.0 0.2606 0 2.0 1e-06 
0.0 0.2607 0 2.0 1e-06 
0.0 0.2608 0 2.0 1e-06 
0.0 0.2609 0 2.0 1e-06 
0.0 0.261 0 2.0 1e-06 
0.0 0.2611 0 2.0 1e-06 
0.0 0.2612 0 2.0 1e-06 
0.0 0.2613 0 2.0 1e-06 
0.0 0.2614 0 2.0 1e-06 
0.0 0.2615 0 2.0 1e-06 
0.0 0.2616 0 2.0 1e-06 
0.0 0.2617 0 2.0 1e-06 
0.0 0.2618 0 2.0 1e-06 
0.0 0.2619 0 2.0 1e-06 
0.0 0.262 0 2.0 1e-06 
0.0 0.2621 0 2.0 1e-06 
0.0 0.2622 0 2.0 1e-06 
0.0 0.2623 0 2.0 1e-06 
0.0 0.2624 0 2.0 1e-06 
0.0 0.2625 0 2.0 1e-06 
0.0 0.2626 0 2.0 1e-06 
0.0 0.2627 0 2.0 1e-06 
0.0 0.2628 0 2.0 1e-06 
0.0 0.2629 0 2.0 1e-06 
0.0 0.263 0 2.0 1e-06 
0.0 0.2631 0 2.0 1e-06 
0.0 0.2632 0 2.0 1e-06 
0.0 0.2633 0 2.0 1e-06 
0.0 0.2634 0 2.0 1e-06 
0.0 0.2635 0 2.0 1e-06 
0.0 0.2636 0 2.0 1e-06 
0.0 0.2637 0 2.0 1e-06 
0.0 0.2638 0 2.0 1e-06 
0.0 0.2639 0 2.0 1e-06 
0.0 0.264 0 2.0 1e-06 
0.0 0.2641 0 2.0 1e-06 
0.0 0.2642 0 2.0 1e-06 
0.0 0.2643 0 2.0 1e-06 
0.0 0.2644 0 2.0 1e-06 
0.0 0.2645 0 2.0 1e-06 
0.0 0.2646 0 2.0 1e-06 
0.0 0.2647 0 2.0 1e-06 
0.0 0.2648 0 2.0 1e-06 
0.0 0.2649 0 2.0 1e-06 
0.0 0.265 0 2.0 1e-06 
0.0 0.2651 0 2.0 1e-06 
0.0 0.2652 0 2.0 1e-06 
0.0 0.2653 0 2.0 1e-06 
0.0 0.2654 0 2.0 1e-06 
0.0 0.2655 0 2.0 1e-06 
0.0 0.2656 0 2.0 1e-06 
0.0 0.2657 0 2.0 1e-06 
0.0 0.2658 0 2.0 1e-06 
0.0 0.2659 0 2.0 1e-06 
0.0 0.266 0 2.0 1e-06 
0.0 0.2661 0 2.0 1e-06 
0.0 0.2662 0 2.0 1e-06 
0.0 0.2663 0 2.0 1e-06 
0.0 0.2664 0 2.0 1e-06 
0.0 0.2665 0 2.0 1e-06 
0.0 0.2666 0 2.0 1e-06 
0.0 0.2667 0 2.0 1e-06 
0.0 0.2668 0 2.0 1e-06 
0.0 0.2669 0 2.0 1e-06 
0.0 0.267 0 2.0 1e-06 
0.0 0.2671 0 2.0 1e-06 
0.0 0.2672 0 2.0 1e-06 
0.0 0.2673 0 2.0 1e-06 
0.0 0.2674 0 2.0 1e-06 
0.0 0.2675 0 2.0 1e-06 
0.0 0.2676 0 2.0 1e-06 
0.0 0.2677 0 2.0 1e-06 
0.0 0.2678 0 2.0 1e-06 
0.0 0.2679 0 2.0 1e-06 
0.0 0.268 0 2.0 1e-06 
0.0 0.2681 0 2.0 1e-06 
0.0 0.2682 0 2.0 1e-06 
0.0 0.2683 0 2.0 1e-06 
0.0 0.2684 0 2.0 1e-06 
0.0 0.2685 0 2.0 1e-06 
0.0 0.2686 0 2.0 1e-06 
0.0 0.2687 0 2.0 1e-06 
0.0 0.2688 0 2.0 1e-06 
0.0 0.2689 0 2.0 1e-06 
0.0 0.269 0 2.0 1e-06 
0.0 0.2691 0 2.0 1e-06 
0.0 0.2692 0 2.0 1e-06 
0.0 0.2693 0 2.0 1e-06 
0.0 0.2694 0 2.0 1e-06 
0.0 0.2695 0 2.0 1e-06 
0.0 0.2696 0 2.0 1e-06 
0.0 0.2697 0 2.0 1e-06 
0.0 0.2698 0 2.0 1e-06 
0.0 0.2699 0 2.0 1e-06 
0.0 0.27 0 2.0 1e-06 
0.0 0.2701 0 2.0 1e-06 
0.0 0.2702 0 2.0 1e-06 
0.0 0.2703 0 2.0 1e-06 
0.0 0.2704 0 2.0 1e-06 
0.0 0.2705 0 2.0 1e-06 
0.0 0.2706 0 2.0 1e-06 
0.0 0.2707 0 2.0 1e-06 
0.0 0.2708 0 2.0 1e-06 
0.0 0.2709 0 2.0 1e-06 
0.0 0.271 0 2.0 1e-06 
0.0 0.2711 0 2.0 1e-06 
0.0 0.2712 0 2.0 1e-06 
0.0 0.2713 0 2.0 1e-06 
0.0 0.2714 0 2.0 1e-06 
0.0 0.2715 0 2.0 1e-06 
0.0 0.2716 0 2.0 1e-06 
0.0 0.2717 0 2.0 1e-06 
0.0 0.2718 0 2.0 1e-06 
0.0 0.2719 0 2.0 1e-06 
0.0 0.272 0 2.0 1e-06 
0.0 0.2721 0 2.0 1e-06 
0.0 0.2722 0 2.0 1e-06 
0.0 0.2723 0 2.0 1e-06 
0.0 0.2724 0 2.0 1e-06 
0.0 0.2725 0 2.0 1e-06 
0.0 0.2726 0 2.0 1e-06 
0.0 0.2727 0 2.0 1e-06 
0.0 0.2728 0 2.0 1e-06 
0.0 0.2729 0 2.0 1e-06 
0.0 0.273 0 2.0 1e-06 
0.0 0.2731 0 2.0 1e-06 
0.0 0.2732 0 2.0 1e-06 
0.0 0.2733 0 2.0 1e-06 
0.0 0.2734 0 2.0 1e-06 
0.0 0.2735 0 2.0 1e-06 
0.0 0.2736 0 2.0 1e-06 
0.0 0.2737 0 2.0 1e-06 
0.0 0.2738 0 2.0 1e-06 
0.0 0.2739 0 2.0 1e-06 
0.0 0.274 0 2.0 1e-06 
0.0 0.2741 0 2.0 1e-06 
0.0 0.2742 0 2.0 1e-06 
0.0 0.2743 0 2.0 1e-06 
0.0 0.2744 0 2.0 1e-06 
0.0 0.2745 0 2.0 1e-06 
0.0 0.2746 0 2.0 1e-06 
0.0 0.2747 0 2.0 1e-06 
0.0 0.2748 0 2.0 1e-06 
0.0 0.2749 0 2.0 1e-06 
0.0 0.275 0 2.0 1e-06 
0.0 0.2751 0 2.0 1e-06 
0.0 0.2752 0 2.0 1e-06 
0.0 0.2753 0 2.0 1e-06 
0.0 0.2754 0 2.0 1e-06 
0.0 0.2755 0 2.0 1e-06 
0.0 0.2756 0 2.0 1e-06 
0.0 0.2757 0 2.0 1e-06 
0.0 0.2758 0 2.0 1e-06 
0.0 0.2759 0 2.0 1e-06 
0.0 0.276 0 2.0 1e-06 
0.0 0.2761 0 2.0 1e-06 
0.0 0.2762 0 2.0 1e-06 
0.0 0.2763 0 2.0 1e-06 
0.0 0.2764 0 2.0 1e-06 
0.0 0.2765 0 2.0 1e-06 
0.0 0.2766 0 2.0 1e-06 
0.0 0.2767 0 2.0 1e-06 
0.0 0.2768 0 2.0 1e-06 
0.0 0.2769 0 2.0 1e-06 
0.0 0.277 0 2.0 1e-06 
0.0 0.2771 0 2.0 1e-06 
0.0 0.2772 0 2.0 1e-06 
0.0 0.2773 0 2.0 1e-06 
0.0 0.2774 0 2.0 1e-06 
0.0 0.2775 0 2.0 1e-06 
0.0 0.2776 0 2.0 1e-06 
0.0 0.2777 0 2.0 1e-06 
0.0 0.2778 0 2.0 1e-06 
0.0 0.2779 0 2.0 1e-06 
0.0 0.278 0 2.0 1e-06 
0.0 0.2781 0 2.0 1e-06 
0.0 0.2782 0 2.0 1e-06 
0.0 0.2783 0 2.0 1e-06 
0.0 0.2784 0 2.0 1e-06 
0.0 0.2785 0 2.0 1e-06 
0.0 0.2786 0 2.0 1e-06 
0.0 0.2787 0 2.0 1e-06 
0.0 0.2788 0 2.0 1e-06 
0.0 0.2789 0 2.0 1e-06 
0.0 0.279 0 2.0 1e-06 
0.0 0.2791 0 2.0 1e-06 
0.0 0.2792 0 2.0 1e-06 
0.0 0.2793 0 2.0 1e-06 
0.0 0.2794 0 2.0 1e-06 
0.0 0.2795 0 2.0 1e-06 
0.0 0.2796 0 2.0 1e-06 
0.0 0.2797 0 2.0 1e-06 
0.0 0.2798 0 2.0 1e-06 
0.0 0.2799 0 2.0 1e-06 
0.0 0.28 0 2.0 1e-06 
0.0 0.2801 0 2.0 1e-06 
0.0 0.2802 0 2.0 1e-06 
0.0 0.2803 0 2.0 1e-06 
0.0 0.2804 0 2.0 1e-06 
0.0 0.2805 0 2.0 1e-06 
0.0 0.2806 0 2.0 1e-06 
0.0 0.2807 0 2.0 1e-06 
0.0 0.2808 0 2.0 1e-06 
0.0 0.2809 0 2.0 1e-06 
0.0 0.281 0 2.0 1e-06 
0.0 0.2811 0 2.0 1e-06 
0.0 0.2812 0 2.0 1e-06 
0.0 0.2813 0 2.0 1e-06 
0.0 0.2814 0 2.0 1e-06 
0.0 0.2815 0 2.0 1e-06 
0.0 0.2816 0 2.0 1e-06 
0.0 0.2817 0 2.0 1e-06 
0.0 0.2818 0 2.0 1e-06 
0.0 0.2819 0 2.0 1e-06 
0.0 0.282 0 2.0 1e-06 
0.0 0.2821 0 2.0 1e-06 
0.0 0.2822 0 2.0 1e-06 
0.0 0.2823 0 2.0 1e-06 
0.0 0.2824 0 2.0 1e-06 
0.0 0.2825 0 2.0 1e-06 
0.0 0.2826 0 2.0 1e-06 
0.0 0.2827 0 2.0 1e-06 
0.0 0.2828 0 2.0 1e-06 
0.0 0.2829 0 2.0 1e-06 
0.0 0.283 0 2.0 1e-06 
0.0 0.2831 0 2.0 1e-06 
0.0 0.2832 0 2.0 1e-06 
0.0 0.2833 0 2.0 1e-06 
0.0 0.2834 0 2.0 1e-06 
0.0 0.2835 0 2.0 1e-06 
0.0 0.2836 0 2.0 1e-06 
0.0 0.2837 0 2.0 1e-06 
0.0 0.2838 0 2.0 1e-06 
0.0 0.2839 0 2.0 1e-06 
0.0 0.284 0 2.0 1e-06 
0.0 0.2841 0 2.0 1e-06 
0.0 0.2842 0 2.0 1e-06 
0.0 0.2843 0 2.0 1e-06 
0.0 0.2844 0 2.0 1e-06 
0.0 0.2845 0 2.0 1e-06 
0.0 0.2846 0 2.0 1e-06 
0.0 0.2847 0 2.0 1e-06 
0.0 0.2848 0 2.0 1e-06 
0.0 0.2849 0 2.0 1e-06 
0.0 0.285 0 2.0 1e-06 
0.0 0.2851 0 2.0 1e-06 
0.0 0.2852 0 2.0 1e-06 
0.0 0.2853 0 2.0 1e-06 
0.0 0.2854 0 2.0 1e-06 
0.0 0.2855 0 2.0 1e-06 
0.0 0.2856 0 2.0 1e-06 
0.0 0.2857 0 2.0 1e-06 
0.0 0.2858 0 2.0 1e-06 
0.0 0.2859 0 2.0 1e-06 
0.0 0.286 0 2.0 1e-06 
0.0 0.2861 0 2.0 1e-06 
0.0 0.2862 0 2.0 1e-06 
0.0 0.2863 0 2.0 1e-06 
0.0 0.2864 0 2.0 1e-06 
0.0 0.2865 0 2.0 1e-06 
0.0 0.2866 0 2.0 1e-06 
0.0 0.2867 0 2.0 1e-06 
0.0 0.2868 0 2.0 1e-06 
0.0 0.2869 0 2.0 1e-06 
0.0 0.287 0 2.0 1e-06 
0.0 0.2871 0 2.0 1e-06 
0.0 0.2872 0 2.0 1e-06 
0.0 0.2873 0 2.0 1e-06 
0.0 0.2874 0 2.0 1e-06 
0.0 0.2875 0 2.0 1e-06 
0.0 0.2876 0 2.0 1e-06 
0.0 0.2877 0 2.0 1e-06 
0.0 0.2878 0 2.0 1e-06 
0.0 0.2879 0 2.0 1e-06 
0.0 0.288 0 2.0 1e-06 
0.0 0.2881 0 2.0 1e-06 
0.0 0.2882 0 2.0 1e-06 
0.0 0.2883 0 2.0 1e-06 
0.0 0.2884 0 2.0 1e-06 
0.0 0.2885 0 2.0 1e-06 
0.0 0.2886 0 2.0 1e-06 
0.0 0.2887 0 2.0 1e-06 
0.0 0.2888 0 2.0 1e-06 
0.0 0.2889 0 2.0 1e-06 
0.0 0.289 0 2.0 1e-06 
0.0 0.2891 0 2.0 1e-06 
0.0 0.2892 0 2.0 1e-06 
0.0 0.2893 0 2.0 1e-06 
0.0 0.2894 0 2.0 1e-06 
0.0 0.2895 0 2.0 1e-06 
0.0 0.2896 0 2.0 1e-06 
0.0 0.2897 0 2.0 1e-06 
0.0 0.2898 0 2.0 1e-06 
0.0 0.2899 0 2.0 1e-06 
0.0 0.29 0 2.0 1e-06 
0.0 0.2901 0 2.0 1e-06 
0.0 0.2902 0 2.0 1e-06 
0.0 0.2903 0 2.0 1e-06 
0.0 0.2904 0 2.0 1e-06 
0.0 0.2905 0 2.0 1e-06 
0.0 0.2906 0 2.0 1e-06 
0.0 0.2907 0 2.0 1e-06 
0.0 0.2908 0 2.0 1e-06 
0.0 0.2909 0 2.0 1e-06 
0.0 0.291 0 2.0 1e-06 
0.0 0.2911 0 2.0 1e-06 
0.0 0.2912 0 2.0 1e-06 
0.0 0.2913 0 2.0 1e-06 
0.0 0.2914 0 2.0 1e-06 
0.0 0.2915 0 2.0 1e-06 
0.0 0.2916 0 2.0 1e-06 
0.0 0.2917 0 2.0 1e-06 
0.0 0.2918 0 2.0 1e-06 
0.0 0.2919 0 2.0 1e-06 
0.0 0.292 0 2.0 1e-06 
0.0 0.2921 0 2.0 1e-06 
0.0 0.2922 0 2.0 1e-06 
0.0 0.2923 0 2.0 1e-06 
0.0 0.2924 0 2.0 1e-06 
0.0 0.2925 0 2.0 1e-06 
0.0 0.2926 0 2.0 1e-06 
0.0 0.2927 0 2.0 1e-06 
0.0 0.2928 0 2.0 1e-06 
0.0 0.2929 0 2.0 1e-06 
0.0 0.293 0 2.0 1e-06 
0.0 0.2931 0 2.0 1e-06 
0.0 0.2932 0 2.0 1e-06 
0.0 0.2933 0 2.0 1e-06 
0.0 0.2934 0 2.0 1e-06 
0.0 0.2935 0 2.0 1e-06 
0.0 0.2936 0 2.0 1e-06 
0.0 0.2937 0 2.0 1e-06 
0.0 0.2938 0 2.0 1e-06 
0.0 0.2939 0 2.0 1e-06 
0.0 0.294 0 2.0 1e-06 
0.0 0.2941 0 2.0 1e-06 
0.0 0.2942 0 2.0 1e-06 
0.0 0.2943 0 2.0 1e-06 
0.0 0.2944 0 2.0 1e-06 
0.0 0.2945 0 2.0 1e-06 
0.0 0.2946 0 2.0 1e-06 
0.0 0.2947 0 2.0 1e-06 
0.0 0.2948 0 2.0 1e-06 
0.0 0.2949 0 2.0 1e-06 
0.0 0.295 0 2.0 1e-06 
0.0 0.2951 0 2.0 1e-06 
0.0 0.2952 0 2.0 1e-06 
0.0 0.2953 0 2.0 1e-06 
0.0 0.2954 0 2.0 1e-06 
0.0 0.2955 0 2.0 1e-06 
0.0 0.2956 0 2.0 1e-06 
0.0 0.2957 0 2.0 1e-06 
0.0 0.2958 0 2.0 1e-06 
0.0 0.2959 0 2.0 1e-06 
0.0 0.296 0 2.0 1e-06 
0.0 0.2961 0 2.0 1e-06 
0.0 0.2962 0 2.0 1e-06 
0.0 0.2963 0 2.0 1e-06 
0.0 0.2964 0 2.0 1e-06 
0.0 0.2965 0 2.0 1e-06 
0.0 0.2966 0 2.0 1e-06 
0.0 0.2967 0 2.0 1e-06 
0.0 0.2968 0 2.0 1e-06 
0.0 0.2969 0 2.0 1e-06 
0.0 0.297 0 2.0 1e-06 
0.0 0.2971 0 2.0 1e-06 
0.0 0.2972 0 2.0 1e-06 
0.0 0.2973 0 2.0 1e-06 
0.0 0.2974 0 2.0 1e-06 
0.0 0.2975 0 2.0 1e-06 
0.0 0.2976 0 2.0 1e-06 
0.0 0.2977 0 2.0 1e-06 
0.0 0.2978 0 2.0 1e-06 
0.0 0.2979 0 2.0 1e-06 
0.0 0.298 0 2.0 1e-06 
0.0 0.2981 0 2.0 1e-06 
0.0 0.2982 0 2.0 1e-06 
0.0 0.2983 0 2.0 1e-06 
0.0 0.2984 0 2.0 1e-06 
0.0 0.2985 0 2.0 1e-06 
0.0 0.2986 0 2.0 1e-06 
0.0 0.2987 0 2.0 1e-06 
0.0 0.2988 0 2.0 1e-06 
0.0 0.2989 0 2.0 1e-06 
0.0 0.299 0 2.0 1e-06 
0.0 0.2991 0 2.0 1e-06 
0.0 0.2992 0 2.0 1e-06 
0.0 0.2993 0 2.0 1e-06 
0.0 0.2994 0 2.0 1e-06 
0.0 0.2995 0 2.0 1e-06 
0.0 0.2996 0 2.0 1e-06 
0.0 0.2997 0 2.0 1e-06 
0.0 0.2998 0 2.0 1e-06 
0.0 0.2999 0 2.0 1e-06 
0.0 0.3 0 2.0 1e-06 
0.0 0.3001 0 2.0 1e-06 
0.0 0.3002 0 2.0 1e-06 
0.0 0.3003 0 2.0 1e-06 
0.0 0.3004 0 2.0 1e-06 
0.0 0.3005 0 2.0 1e-06 
0.0 0.3006 0 2.0 1e-06 
0.0 0.3007 0 2.0 1e-06 
0.0 0.3008 0 2.0 1e-06 
0.0 0.3009 0 2.0 1e-06 
0.0 0.301 0 2.0 1e-06 
0.0 0.3011 0 2.0 1e-06 
0.0 0.3012 0 2.0 1e-06 
0.0 0.3013 0 2.0 1e-06 
0.0 0.3014 0 2.0 1e-06 
0.0 0.3015 0 2.0 1e-06 
0.0 0.3016 0 2.0 1e-06 
0.0 0.3017 0 2.0 1e-06 
0.0 0.3018 0 2.0 1e-06 
0.0 0.3019 0 2.0 1e-06 
0.0 0.302 0 2.0 1e-06 
0.0 0.3021 0 2.0 1e-06 
0.0 0.3022 0 2.0 1e-06 
0.0 0.3023 0 2.0 1e-06 
0.0 0.3024 0 2.0 1e-06 
0.0 0.3025 0 2.0 1e-06 
0.0 0.3026 0 2.0 1e-06 
0.0 0.3027 0 2.0 1e-06 
0.0 0.3028 0 2.0 1e-06 
0.0 0.3029 0 2.0 1e-06 
0.0 0.303 0 2.0 1e-06 
0.0 0.3031 0 2.0 1e-06 
0.0 0.3032 0 2.0 1e-06 
0.0 0.3033 0 2.0 1e-06 
0.0 0.3034 0 2.0 1e-06 
0.0 0.3035 0 2.0 1e-06 
0.0 0.3036 0 2.0 1e-06 
0.0 0.3037 0 2.0 1e-06 
0.0 0.3038 0 2.0 1e-06 
0.0 0.3039 0 2.0 1e-06 
0.0 0.304 0 2.0 1e-06 
0.0 0.3041 0 2.0 1e-06 
0.0 0.3042 0 2.0 1e-06 
0.0 0.3043 0 2.0 1e-06 
0.0 0.3044 0 2.0 1e-06 
0.0 0.3045 0 2.0 1e-06 
0.0 0.3046 0 2.0 1e-06 
0.0 0.3047 0 2.0 1e-06 
0.0 0.3048 0 2.0 1e-06 
0.0 0.3049 0 2.0 1e-06 
0.0 0.305 0 2.0 1e-06 
0.0 0.3051 0 2.0 1e-06 
0.0 0.3052 0 2.0 1e-06 
0.0 0.3053 0 2.0 1e-06 
0.0 0.3054 0 2.0 1e-06 
0.0 0.3055 0 2.0 1e-06 
0.0 0.3056 0 2.0 1e-06 
0.0 0.3057 0 2.0 1e-06 
0.0 0.3058 0 2.0 1e-06 
0.0 0.3059 0 2.0 1e-06 
0.0 0.306 0 2.0 1e-06 
0.0 0.3061 0 2.0 1e-06 
0.0 0.3062 0 2.0 1e-06 
0.0 0.3063 0 2.0 1e-06 
0.0 0.3064 0 2.0 1e-06 
0.0 0.3065 0 2.0 1e-06 
0.0 0.3066 0 2.0 1e-06 
0.0 0.3067 0 2.0 1e-06 
0.0 0.3068 0 2.0 1e-06 
0.0 0.3069 0 2.0 1e-06 
0.0 0.307 0 2.0 1e-06 
0.0 0.3071 0 2.0 1e-06 
0.0 0.3072 0 2.0 1e-06 
0.0 0.3073 0 2.0 1e-06 
0.0 0.3074 0 2.0 1e-06 
0.0 0.3075 0 2.0 1e-06 
0.0 0.3076 0 2.0 1e-06 
0.0 0.3077 0 2.0 1e-06 
0.0 0.3078 0 2.0 1e-06 
0.0 0.3079 0 2.0 1e-06 
0.0 0.308 0 2.0 1e-06 
0.0 0.3081 0 2.0 1e-06 
0.0 0.3082 0 2.0 1e-06 
0.0 0.3083 0 2.0 1e-06 
0.0 0.3084 0 2.0 1e-06 
0.0 0.3085 0 2.0 1e-06 
0.0 0.3086 0 2.0 1e-06 
0.0 0.3087 0 2.0 1e-06 
0.0 0.3088 0 2.0 1e-06 
0.0 0.3089 0 2.0 1e-06 
0.0 0.309 0 2.0 1e-06 
0.0 0.3091 0 2.0 1e-06 
0.0 0.3092 0 2.0 1e-06 
0.0 0.3093 0 2.0 1e-06 
0.0 0.3094 0 2.0 1e-06 
0.0 0.3095 0 2.0 1e-06 
0.0 0.3096 0 2.0 1e-06 
0.0 0.3097 0 2.0 1e-06 
0.0 0.3098 0 2.0 1e-06 
0.0 0.3099 0 2.0 1e-06 
0.0 0.31 0 2.0 1e-06 
0.0 0.3101 0 2.0 1e-06 
0.0 0.3102 0 2.0 1e-06 
0.0 0.3103 0 2.0 1e-06 
0.0 0.3104 0 2.0 1e-06 
0.0 0.3105 0 2.0 1e-06 
0.0 0.3106 0 2.0 1e-06 
0.0 0.3107 0 2.0 1e-06 
0.0 0.3108 0 2.0 1e-06 
0.0 0.3109 0 2.0 1e-06 
0.0 0.311 0 2.0 1e-06 
0.0 0.3111 0 2.0 1e-06 
0.0 0.3112 0 2.0 1e-06 
0.0 0.3113 0 2.0 1e-06 
0.0 0.3114 0 2.0 1e-06 
0.0 0.3115 0 2.0 1e-06 
0.0 0.3116 0 2.0 1e-06 
0.0 0.3117 0 2.0 1e-06 
0.0 0.3118 0 2.0 1e-06 
0.0 0.3119 0 2.0 1e-06 
0.0 0.312 0 2.0 1e-06 
0.0 0.3121 0 2.0 1e-06 
0.0 0.3122 0 2.0 1e-06 
0.0 0.3123 0 2.0 1e-06 
0.0 0.3124 0 2.0 1e-06 
0.0 0.3125 0 2.0 1e-06 
0.0 0.3126 0 2.0 1e-06 
0.0 0.3127 0 2.0 1e-06 
0.0 0.3128 0 2.0 1e-06 
0.0 0.3129 0 2.0 1e-06 
0.0 0.313 0 2.0 1e-06 
0.0 0.3131 0 2.0 1e-06 
0.0 0.3132 0 2.0 1e-06 
0.0 0.3133 0 2.0 1e-06 
0.0 0.3134 0 2.0 1e-06 
0.0 0.3135 0 2.0 1e-06 
0.0 0.3136 0 2.0 1e-06 
0.0 0.3137 0 2.0 1e-06 
0.0 0.3138 0 2.0 1e-06 
0.0 0.3139 0 2.0 1e-06 
0.0 0.314 0 2.0 1e-06 
0.0 0.3141 0 2.0 1e-06 
0.0 0.3142 0 2.0 1e-06 
0.0 0.3143 0 2.0 1e-06 
0.0 0.3144 0 2.0 1e-06 
0.0 0.3145 0 2.0 1e-06 
0.0 0.3146 0 2.0 1e-06 
0.0 0.3147 0 2.0 1e-06 
0.0 0.3148 0 2.0 1e-06 
0.0 0.3149 0 2.0 1e-06 
0.0 0.315 0 2.0 1e-06 
0.0 0.3151 0 2.0 1e-06 
0.0 0.3152 0 2.0 1e-06 
0.0 0.3153 0 2.0 1e-06 
0.0 0.3154 0 2.0 1e-06 
0.0 0.3155 0 2.0 1e-06 
0.0 0.3156 0 2.0 1e-06 
0.0 0.3157 0 2.0 1e-06 
0.0 0.3158 0 2.0 1e-06 
0.0 0.3159 0 2.0 1e-06 
0.0 0.316 0 2.0 1e-06 
0.0 0.3161 0 2.0 1e-06 
0.0 0.3162 0 2.0 1e-06 
0.0 0.3163 0 2.0 1e-06 
0.0 0.3164 0 2.0 1e-06 
0.0 0.3165 0 2.0 1e-06 
0.0 0.3166 0 2.0 1e-06 
0.0 0.3167 0 2.0 1e-06 
0.0 0.3168 0 2.0 1e-06 
0.0 0.3169 0 2.0 1e-06 
0.0 0.317 0 2.0 1e-06 
0.0 0.3171 0 2.0 1e-06 
0.0 0.3172 0 2.0 1e-06 
0.0 0.3173 0 2.0 1e-06 
0.0 0.3174 0 2.0 1e-06 
0.0 0.3175 0 2.0 1e-06 
0.0 0.3176 0 2.0 1e-06 
0.0 0.3177 0 2.0 1e-06 
0.0 0.3178 0 2.0 1e-06 
0.0 0.3179 0 2.0 1e-06 
0.0 0.318 0 2.0 1e-06 
0.0 0.3181 0 2.0 1e-06 
0.0 0.3182 0 2.0 1e-06 
0.0 0.3183 0 2.0 1e-06 
0.0 0.3184 0 2.0 1e-06 
0.0 0.3185 0 2.0 1e-06 
0.0 0.3186 0 2.0 1e-06 
0.0 0.3187 0 2.0 1e-06 
0.0 0.3188 0 2.0 1e-06 
0.0 0.3189 0 2.0 1e-06 
0.0 0.319 0 2.0 1e-06 
0.0 0.3191 0 2.0 1e-06 
0.0 0.3192 0 2.0 1e-06 
0.0 0.3193 0 2.0 1e-06 
0.0 0.3194 0 2.0 1e-06 
0.0 0.3195 0 2.0 1e-06 
0.0 0.3196 0 2.0 1e-06 
0.0 0.3197 0 2.0 1e-06 
0.0 0.3198 0 2.0 1e-06 
0.0 0.3199 0 2.0 1e-06 
0.0 0.32 0 2.0 1e-06 
0.0 0.3201 0 2.0 1e-06 
0.0 0.3202 0 2.0 1e-06 
0.0 0.3203 0 2.0 1e-06 
0.0 0.3204 0 2.0 1e-06 
0.0 0.3205 0 2.0 1e-06 
0.0 0.3206 0 2.0 1e-06 
0.0 0.3207 0 2.0 1e-06 
0.0 0.3208 0 2.0 1e-06 
0.0 0.3209 0 2.0 1e-06 
0.0 0.321 0 2.0 1e-06 
0.0 0.3211 0 2.0 1e-06 
0.0 0.3212 0 2.0 1e-06 
0.0 0.3213 0 2.0 1e-06 
0.0 0.3214 0 2.0 1e-06 
0.0 0.3215 0 2.0 1e-06 
0.0 0.3216 0 2.0 1e-06 
0.0 0.3217 0 2.0 1e-06 
0.0 0.3218 0 2.0 1e-06 
0.0 0.3219 0 2.0 1e-06 
0.0 0.322 0 2.0 1e-06 
0.0 0.3221 0 2.0 1e-06 
0.0 0.3222 0 2.0 1e-06 
0.0 0.3223 0 2.0 1e-06 
0.0 0.3224 0 2.0 1e-06 
0.0 0.3225 0 2.0 1e-06 
0.0 0.3226 0 2.0 1e-06 
0.0 0.3227 0 2.0 1e-06 
0.0 0.3228 0 2.0 1e-06 
0.0 0.3229 0 2.0 1e-06 
0.0 0.323 0 2.0 1e-06 
0.0 0.3231 0 2.0 1e-06 
0.0 0.3232 0 2.0 1e-06 
0.0 0.3233 0 2.0 1e-06 
0.0 0.3234 0 2.0 1e-06 
0.0 0.3235 0 2.0 1e-06 
0.0 0.3236 0 2.0 1e-06 
0.0 0.3237 0 2.0 1e-06 
0.0 0.3238 0 2.0 1e-06 
0.0 0.3239 0 2.0 1e-06 
0.0 0.324 0 2.0 1e-06 
0.0 0.3241 0 2.0 1e-06 
0.0 0.3242 0 2.0 1e-06 
0.0 0.3243 0 2.0 1e-06 
0.0 0.3244 0 2.0 1e-06 
0.0 0.3245 0 2.0 1e-06 
0.0 0.3246 0 2.0 1e-06 
0.0 0.3247 0 2.0 1e-06 
0.0 0.3248 0 2.0 1e-06 
0.0 0.3249 0 2.0 1e-06 
0.0 0.325 0 2.0 1e-06 
0.0 0.3251 0 2.0 1e-06 
0.0 0.3252 0 2.0 1e-06 
0.0 0.3253 0 2.0 1e-06 
0.0 0.3254 0 2.0 1e-06 
0.0 0.3255 0 2.0 1e-06 
0.0 0.3256 0 2.0 1e-06 
0.0 0.3257 0 2.0 1e-06 
0.0 0.3258 0 2.0 1e-06 
0.0 0.3259 0 2.0 1e-06 
0.0 0.326 0 2.0 1e-06 
0.0 0.3261 0 2.0 1e-06 
0.0 0.3262 0 2.0 1e-06 
0.0 0.3263 0 2.0 1e-06 
0.0 0.3264 0 2.0 1e-06 
0.0 0.3265 0 2.0 1e-06 
0.0 0.3266 0 2.0 1e-06 
0.0 0.3267 0 2.0 1e-06 
0.0 0.3268 0 2.0 1e-06 
0.0 0.3269 0 2.0 1e-06 
0.0 0.327 0 2.0 1e-06 
0.0 0.3271 0 2.0 1e-06 
0.0 0.3272 0 2.0 1e-06 
0.0 0.3273 0 2.0 1e-06 
0.0 0.3274 0 2.0 1e-06 
0.0 0.3275 0 2.0 1e-06 
0.0 0.3276 0 2.0 1e-06 
0.0 0.3277 0 2.0 1e-06 
0.0 0.3278 0 2.0 1e-06 
0.0 0.3279 0 2.0 1e-06 
0.0 0.328 0 2.0 1e-06 
0.0 0.3281 0 2.0 1e-06 
0.0 0.3282 0 2.0 1e-06 
0.0 0.3283 0 2.0 1e-06 
0.0 0.3284 0 2.0 1e-06 
0.0 0.3285 0 2.0 1e-06 
0.0 0.3286 0 2.0 1e-06 
0.0 0.3287 0 2.0 1e-06 
0.0 0.3288 0 2.0 1e-06 
0.0 0.3289 0 2.0 1e-06 
0.0 0.329 0 2.0 1e-06 
0.0 0.3291 0 2.0 1e-06 
0.0 0.3292 0 2.0 1e-06 
0.0 0.3293 0 2.0 1e-06 
0.0 0.3294 0 2.0 1e-06 
0.0 0.3295 0 2.0 1e-06 
0.0 0.3296 0 2.0 1e-06 
0.0 0.3297 0 2.0 1e-06 
0.0 0.3298 0 2.0 1e-06 
0.0 0.3299 0 2.0 1e-06 
0.0 0.33 0 2.0 1e-06 
0.0 0.3301 0 2.0 1e-06 
0.0 0.3302 0 2.0 1e-06 
0.0 0.3303 0 2.0 1e-06 
0.0 0.3304 0 2.0 1e-06 
0.0 0.3305 0 2.0 1e-06 
0.0 0.3306 0 2.0 1e-06 
0.0 0.3307 0 2.0 1e-06 
0.0 0.3308 0 2.0 1e-06 
0.0 0.3309 0 2.0 1e-06 
0.0 0.331 0 2.0 1e-06 
0.0 0.3311 0 2.0 1e-06 
0.0 0.3312 0 2.0 1e-06 
0.0 0.3313 0 2.0 1e-06 
0.0 0.3314 0 2.0 1e-06 
0.0 0.3315 0 2.0 1e-06 
0.0 0.3316 0 2.0 1e-06 
0.0 0.3317 0 2.0 1e-06 
0.0 0.3318 0 2.0 1e-06 
0.0 0.3319 0 2.0 1e-06 
0.0 0.332 0 2.0 1e-06 
0.0 0.3321 0 2.0 1e-06 
0.0 0.3322 0 2.0 1e-06 
0.0 0.3323 0 2.0 1e-06 
0.0 0.3324 0 2.0 1e-06 
0.0 0.3325 0 2.0 1e-06 
0.0 0.3326 0 2.0 1e-06 
0.0 0.3327 0 2.0 1e-06 
0.0 0.3328 0 2.0 1e-06 
0.0 0.3329 0 2.0 1e-06 
0.0 0.333 0 2.0 1e-06 
0.0 0.3331 0 2.0 1e-06 
0.0 0.3332 0 2.0 1e-06 
0.0 0.3333 0 2.0 1e-06 
0.0 0.3334 0 2.0 1e-06 
0.0 0.3335 0 2.0 1e-06 
0.0 0.3336 0 2.0 1e-06 
0.0 0.3337 0 2.0 1e-06 
0.0 0.3338 0 2.0 1e-06 
0.0 0.3339 0 2.0 1e-06 
0.0 0.334 0 2.0 1e-06 
0.0 0.3341 0 2.0 1e-06 
0.0 0.3342 0 2.0 1e-06 
0.0 0.3343 0 2.0 1e-06 
0.0 0.3344 0 2.0 1e-06 
0.0 0.3345 0 2.0 1e-06 
0.0 0.3346 0 2.0 1e-06 
0.0 0.3347 0 2.0 1e-06 
0.0 0.3348 0 2.0 1e-06 
0.0 0.3349 0 2.0 1e-06 
0.0 0.335 0 2.0 1e-06 
0.0 0.3351 0 2.0 1e-06 
0.0 0.3352 0 2.0 1e-06 
0.0 0.3353 0 2.0 1e-06 
0.0 0.3354 0 2.0 1e-06 
0.0 0.3355 0 2.0 1e-06 
0.0 0.3356 0 2.0 1e-06 
0.0 0.3357 0 2.0 1e-06 
0.0 0.3358 0 2.0 1e-06 
0.0 0.3359 0 2.0 1e-06 
0.0 0.336 0 2.0 1e-06 
0.0 0.3361 0 2.0 1e-06 
0.0 0.3362 0 2.0 1e-06 
0.0 0.3363 0 2.0 1e-06 
0.0 0.3364 0 2.0 1e-06 
0.0 0.3365 0 2.0 1e-06 
0.0 0.3366 0 2.0 1e-06 
0.0 0.3367 0 2.0 1e-06 
0.0 0.3368 0 2.0 1e-06 
0.0 0.3369 0 2.0 1e-06 
0.0 0.337 0 2.0 1e-06 
0.0 0.3371 0 2.0 1e-06 
0.0 0.3372 0 2.0 1e-06 
0.0 0.3373 0 2.0 1e-06 
0.0 0.3374 0 2.0 1e-06 
0.0 0.3375 0 2.0 1e-06 
0.0 0.3376 0 2.0 1e-06 
0.0 0.3377 0 2.0 1e-06 
0.0 0.3378 0 2.0 1e-06 
0.0 0.3379 0 2.0 1e-06 
0.0 0.338 0 2.0 1e-06 
0.0 0.3381 0 2.0 1e-06 
0.0 0.3382 0 2.0 1e-06 
0.0 0.3383 0 2.0 1e-06 
0.0 0.3384 0 2.0 1e-06 
0.0 0.3385 0 2.0 1e-06 
0.0 0.3386 0 2.0 1e-06 
0.0 0.3387 0 2.0 1e-06 
0.0 0.3388 0 2.0 1e-06 
0.0 0.3389 0 2.0 1e-06 
0.0 0.339 0 2.0 1e-06 
0.0 0.3391 0 2.0 1e-06 
0.0 0.3392 0 2.0 1e-06 
0.0 0.3393 0 2.0 1e-06 
0.0 0.3394 0 2.0 1e-06 
0.0 0.3395 0 2.0 1e-06 
0.0 0.3396 0 2.0 1e-06 
0.0 0.3397 0 2.0 1e-06 
0.0 0.3398 0 2.0 1e-06 
0.0 0.3399 0 2.0 1e-06 
0.0 0.34 0 2.0 1e-06 
0.0 0.3401 0 2.0 1e-06 
0.0 0.3402 0 2.0 1e-06 
0.0 0.3403 0 2.0 1e-06 
0.0 0.3404 0 2.0 1e-06 
0.0 0.3405 0 2.0 1e-06 
0.0 0.3406 0 2.0 1e-06 
0.0 0.3407 0 2.0 1e-06 
0.0 0.3408 0 2.0 1e-06 
0.0 0.3409 0 2.0 1e-06 
0.0 0.341 0 2.0 1e-06 
0.0 0.3411 0 2.0 1e-06 
0.0 0.3412 0 2.0 1e-06 
0.0 0.3413 0 2.0 1e-06 
0.0 0.3414 0 2.0 1e-06 
0.0 0.3415 0 2.0 1e-06 
0.0 0.3416 0 2.0 1e-06 
0.0 0.3417 0 2.0 1e-06 
0.0 0.3418 0 2.0 1e-06 
0.0 0.3419 0 2.0 1e-06 
0.0 0.342 0 2.0 1e-06 
0.0 0.3421 0 2.0 1e-06 
0.0 0.3422 0 2.0 1e-06 
0.0 0.3423 0 2.0 1e-06 
0.0 0.3424 0 2.0 1e-06 
0.0 0.3425 0 2.0 1e-06 
0.0 0.3426 0 2.0 1e-06 
0.0 0.3427 0 2.0 1e-06 
0.0 0.3428 0 2.0 1e-06 
0.0 0.3429 0 2.0 1e-06 
0.0 0.343 0 2.0 1e-06 
0.0 0.3431 0 2.0 1e-06 
0.0 0.3432 0 2.0 1e-06 
0.0 0.3433 0 2.0 1e-06 
0.0 0.3434 0 2.0 1e-06 
0.0 0.3435 0 2.0 1e-06 
0.0 0.3436 0 2.0 1e-06 
0.0 0.3437 0 2.0 1e-06 
0.0 0.3438 0 2.0 1e-06 
0.0 0.3439 0 2.0 1e-06 
0.0 0.344 0 2.0 1e-06 
0.0 0.3441 0 2.0 1e-06 
0.0 0.3442 0 2.0 1e-06 
0.0 0.3443 0 2.0 1e-06 
0.0 0.3444 0 2.0 1e-06 
0.0 0.3445 0 2.0 1e-06 
0.0 0.3446 0 2.0 1e-06 
0.0 0.3447 0 2.0 1e-06 
0.0 0.3448 0 2.0 1e-06 
0.0 0.3449 0 2.0 1e-06 
0.0 0.345 0 2.0 1e-06 
0.0 0.3451 0 2.0 1e-06 
0.0 0.3452 0 2.0 1e-06 
0.0 0.3453 0 2.0 1e-06 
0.0 0.3454 0 2.0 1e-06 
0.0 0.3455 0 2.0 1e-06 
0.0 0.3456 0 2.0 1e-06 
0.0 0.3457 0 2.0 1e-06 
0.0 0.3458 0 2.0 1e-06 
0.0 0.3459 0 2.0 1e-06 
0.0 0.346 0 2.0 1e-06 
0.0 0.3461 0 2.0 1e-06 
0.0 0.3462 0 2.0 1e-06 
0.0 0.3463 0 2.0 1e-06 
0.0 0.3464 0 2.0 1e-06 
0.0 0.3465 0 2.0 1e-06 
0.0 0.3466 0 2.0 1e-06 
0.0 0.3467 0 2.0 1e-06 
0.0 0.3468 0 2.0 1e-06 
0.0 0.3469 0 2.0 1e-06 
0.0 0.347 0 2.0 1e-06 
0.0 0.3471 0 2.0 1e-06 
0.0 0.3472 0 2.0 1e-06 
0.0 0.3473 0 2.0 1e-06 
0.0 0.3474 0 2.0 1e-06 
0.0 0.3475 0 2.0 1e-06 
0.0 0.3476 0 2.0 1e-06 
0.0 0.3477 0 2.0 1e-06 
0.0 0.3478 0 2.0 1e-06 
0.0 0.3479 0 2.0 1e-06 
0.0 0.348 0 2.0 1e-06 
0.0 0.3481 0 2.0 1e-06 
0.0 0.3482 0 2.0 1e-06 
0.0 0.3483 0 2.0 1e-06 
0.0 0.3484 0 2.0 1e-06 
0.0 0.3485 0 2.0 1e-06 
0.0 0.3486 0 2.0 1e-06 
0.0 0.3487 0 2.0 1e-06 
0.0 0.3488 0 2.0 1e-06 
0.0 0.3489 0 2.0 1e-06 
0.0 0.349 0 2.0 1e-06 
0.0 0.3491 0 2.0 1e-06 
0.0 0.3492 0 2.0 1e-06 
0.0 0.3493 0 2.0 1e-06 
0.0 0.3494 0 2.0 1e-06 
0.0 0.3495 0 2.0 1e-06 
0.0 0.3496 0 2.0 1e-06 
0.0 0.3497 0 2.0 1e-06 
0.0 0.3498 0 2.0 1e-06 
0.0 0.3499 0 2.0 1e-06 
0.0 0.35 0 2.0 1e-06 
0.0 0.3501 0 2.0 1e-06 
0.0 0.3502 0 2.0 1e-06 
0.0 0.3503 0 2.0 1e-06 
0.0 0.3504 0 2.0 1e-06 
0.0 0.3505 0 2.0 1e-06 
0.0 0.3506 0 2.0 1e-06 
0.0 0.3507 0 2.0 1e-06 
0.0 0.3508 0 2.0 1e-06 
0.0 0.3509 0 2.0 1e-06 
0.0 0.351 0 2.0 1e-06 
0.0 0.3511 0 2.0 1e-06 
0.0 0.3512 0 2.0 1e-06 
0.0 0.3513 0 2.0 1e-06 
0.0 0.3514 0 2.0 1e-06 
0.0 0.3515 0 2.0 1e-06 
0.0 0.3516 0 2.0 1e-06 
0.0 0.3517 0 2.0 1e-06 
0.0 0.3518 0 2.0 1e-06 
0.0 0.3519 0 2.0 1e-06 
0.0 0.352 0 2.0 1e-06 
0.0 0.3521 0 2.0 1e-06 
0.0 0.3522 0 2.0 1e-06 
0.0 0.3523 0 2.0 1e-06 
0.0 0.3524 0 2.0 1e-06 
0.0 0.3525 0 2.0 1e-06 
0.0 0.3526 0 2.0 1e-06 
0.0 0.3527 0 2.0 1e-06 
0.0 0.3528 0 2.0 1e-06 
0.0 0.3529 0 2.0 1e-06 
0.0 0.353 0 2.0 1e-06 
0.0 0.3531 0 2.0 1e-06 
0.0 0.3532 0 2.0 1e-06 
0.0 0.3533 0 2.0 1e-06 
0.0 0.3534 0 2.0 1e-06 
0.0 0.3535 0 2.0 1e-06 
0.0 0.3536 0 2.0 1e-06 
0.0 0.3537 0 2.0 1e-06 
0.0 0.3538 0 2.0 1e-06 
0.0 0.3539 0 2.0 1e-06 
0.0 0.354 0 2.0 1e-06 
0.0 0.3541 0 2.0 1e-06 
0.0 0.3542 0 2.0 1e-06 
0.0 0.3543 0 2.0 1e-06 
0.0 0.3544 0 2.0 1e-06 
0.0 0.3545 0 2.0 1e-06 
0.0 0.3546 0 2.0 1e-06 
0.0 0.3547 0 2.0 1e-06 
0.0 0.3548 0 2.0 1e-06 
0.0 0.3549 0 2.0 1e-06 
0.0 0.355 0 2.0 1e-06 
0.0 0.3551 0 2.0 1e-06 
0.0 0.3552 0 2.0 1e-06 
0.0 0.3553 0 2.0 1e-06 
0.0 0.3554 0 2.0 1e-06 
0.0 0.3555 0 2.0 1e-06 
0.0 0.3556 0 2.0 1e-06 
0.0 0.3557 0 2.0 1e-06 
0.0 0.3558 0 2.0 1e-06 
0.0 0.3559 0 2.0 1e-06 
0.0 0.356 0 2.0 1e-06 
0.0 0.3561 0 2.0 1e-06 
0.0 0.3562 0 2.0 1e-06 
0.0 0.3563 0 2.0 1e-06 
0.0 0.3564 0 2.0 1e-06 
0.0 0.3565 0 2.0 1e-06 
0.0 0.3566 0 2.0 1e-06 
0.0 0.3567 0 2.0 1e-06 
0.0 0.3568 0 2.0 1e-06 
0.0 0.3569 0 2.0 1e-06 
0.0 0.357 0 2.0 1e-06 
0.0 0.3571 0 2.0 1e-06 
0.0 0.3572 0 2.0 1e-06 
0.0 0.3573 0 2.0 1e-06 
0.0 0.3574 0 2.0 1e-06 
0.0 0.3575 0 2.0 1e-06 
0.0 0.3576 0 2.0 1e-06 
0.0 0.3577 0 2.0 1e-06 
0.0 0.3578 0 2.0 1e-06 
0.0 0.3579 0 2.0 1e-06 
0.0 0.358 0 2.0 1e-06 
0.0 0.3581 0 2.0 1e-06 
0.0 0.3582 0 2.0 1e-06 
0.0 0.3583 0 2.0 1e-06 
0.0 0.3584 0 2.0 1e-06 
0.0 0.3585 0 2.0 1e-06 
0.0 0.3586 0 2.0 1e-06 
0.0 0.3587 0 2.0 1e-06 
0.0 0.3588 0 2.0 1e-06 
0.0 0.3589 0 2.0 1e-06 
0.0 0.359 0 2.0 1e-06 
0.0 0.3591 0 2.0 1e-06 
0.0 0.3592 0 2.0 1e-06 
0.0 0.3593 0 2.0 1e-06 
0.0 0.3594 0 2.0 1e-06 
0.0 0.3595 0 2.0 1e-06 
0.0 0.3596 0 2.0 1e-06 
0.0 0.3597 0 2.0 1e-06 
0.0 0.3598 0 2.0 1e-06 
0.0 0.3599 0 2.0 1e-06 
0.0 0.36 0 2.0 1e-06 
0.0 0.3601 0 2.0 1e-06 
0.0 0.3602 0 2.0 1e-06 
0.0 0.3603 0 2.0 1e-06 
0.0 0.3604 0 2.0 1e-06 
0.0 0.3605 0 2.0 1e-06 
0.0 0.3606 0 2.0 1e-06 
0.0 0.3607 0 2.0 1e-06 
0.0 0.3608 0 2.0 1e-06 
0.0 0.3609 0 2.0 1e-06 
0.0 0.361 0 2.0 1e-06 
0.0 0.3611 0 2.0 1e-06 
0.0 0.3612 0 2.0 1e-06 
0.0 0.3613 0 2.0 1e-06 
0.0 0.3614 0 2.0 1e-06 
0.0 0.3615 0 2.0 1e-06 
0.0 0.3616 0 2.0 1e-06 
0.0 0.3617 0 2.0 1e-06 
0.0 0.3618 0 2.0 1e-06 
0.0 0.3619 0 2.0 1e-06 
0.0 0.362 0 2.0 1e-06 
0.0 0.3621 0 2.0 1e-06 
0.0 0.3622 0 2.0 1e-06 
0.0 0.3623 0 2.0 1e-06 
0.0 0.3624 0 2.0 1e-06 
0.0 0.3625 0 2.0 1e-06 
0.0 0.3626 0 2.0 1e-06 
0.0 0.3627 0 2.0 1e-06 
0.0 0.3628 0 2.0 1e-06 
0.0 0.3629 0 2.0 1e-06 
0.0 0.363 0 2.0 1e-06 
0.0 0.3631 0 2.0 1e-06 
0.0 0.3632 0 2.0 1e-06 
0.0 0.3633 0 2.0 1e-06 
0.0 0.3634 0 2.0 1e-06 
0.0 0.3635 0 2.0 1e-06 
0.0 0.3636 0 2.0 1e-06 
0.0 0.3637 0 2.0 1e-06 
0.0 0.3638 0 2.0 1e-06 
0.0 0.3639 0 2.0 1e-06 
0.0 0.364 0 2.0 1e-06 
0.0 0.3641 0 2.0 1e-06 
0.0 0.3642 0 2.0 1e-06 
0.0 0.3643 0 2.0 1e-06 
0.0 0.3644 0 2.0 1e-06 
0.0 0.3645 0 2.0 1e-06 
0.0 0.3646 0 2.0 1e-06 
0.0 0.3647 0 2.0 1e-06 
0.0 0.3648 0 2.0 1e-06 
0.0 0.3649 0 2.0 1e-06 
0.0 0.365 0 2.0 1e-06 
0.0 0.3651 0 2.0 1e-06 
0.0 0.3652 0 2.0 1e-06 
0.0 0.3653 0 2.0 1e-06 
0.0 0.3654 0 2.0 1e-06 
0.0 0.3655 0 2.0 1e-06 
0.0 0.3656 0 2.0 1e-06 
0.0 0.3657 0 2.0 1e-06 
0.0 0.3658 0 2.0 1e-06 
0.0 0.3659 0 2.0 1e-06 
0.0 0.366 0 2.0 1e-06 
0.0 0.3661 0 2.0 1e-06 
0.0 0.3662 0 2.0 1e-06 
0.0 0.3663 0 2.0 1e-06 
0.0 0.3664 0 2.0 1e-06 
0.0 0.3665 0 2.0 1e-06 
0.0 0.3666 0 2.0 1e-06 
0.0 0.3667 0 2.0 1e-06 
0.0 0.3668 0 2.0 1e-06 
0.0 0.3669 0 2.0 1e-06 
0.0 0.367 0 2.0 1e-06 
0.0 0.3671 0 2.0 1e-06 
0.0 0.3672 0 2.0 1e-06 
0.0 0.3673 0 2.0 1e-06 
0.0 0.3674 0 2.0 1e-06 
0.0 0.3675 0 2.0 1e-06 
0.0 0.3676 0 2.0 1e-06 
0.0 0.3677 0 2.0 1e-06 
0.0 0.3678 0 2.0 1e-06 
0.0 0.3679 0 2.0 1e-06 
0.0 0.368 0 2.0 1e-06 
0.0 0.3681 0 2.0 1e-06 
0.0 0.3682 0 2.0 1e-06 
0.0 0.3683 0 2.0 1e-06 
0.0 0.3684 0 2.0 1e-06 
0.0 0.3685 0 2.0 1e-06 
0.0 0.3686 0 2.0 1e-06 
0.0 0.3687 0 2.0 1e-06 
0.0 0.3688 0 2.0 1e-06 
0.0 0.3689 0 2.0 1e-06 
0.0 0.369 0 2.0 1e-06 
0.0 0.3691 0 2.0 1e-06 
0.0 0.3692 0 2.0 1e-06 
0.0 0.3693 0 2.0 1e-06 
0.0 0.3694 0 2.0 1e-06 
0.0 0.3695 0 2.0 1e-06 
0.0 0.3696 0 2.0 1e-06 
0.0 0.3697 0 2.0 1e-06 
0.0 0.3698 0 2.0 1e-06 
0.0 0.3699 0 2.0 1e-06 
0.0 0.37 0 2.0 1e-06 
0.0 0.3701 0 2.0 1e-06 
0.0 0.3702 0 2.0 1e-06 
0.0 0.3703 0 2.0 1e-06 
0.0 0.3704 0 2.0 1e-06 
0.0 0.3705 0 2.0 1e-06 
0.0 0.3706 0 2.0 1e-06 
0.0 0.3707 0 2.0 1e-06 
0.0 0.3708 0 2.0 1e-06 
0.0 0.3709 0 2.0 1e-06 
0.0 0.371 0 2.0 1e-06 
0.0 0.3711 0 2.0 1e-06 
0.0 0.3712 0 2.0 1e-06 
0.0 0.3713 0 2.0 1e-06 
0.0 0.3714 0 2.0 1e-06 
0.0 0.3715 0 2.0 1e-06 
0.0 0.3716 0 2.0 1e-06 
0.0 0.3717 0 2.0 1e-06 
0.0 0.3718 0 2.0 1e-06 
0.0 0.3719 0 2.0 1e-06 
0.0 0.372 0 2.0 1e-06 
0.0 0.3721 0 2.0 1e-06 
0.0 0.3722 0 2.0 1e-06 
0.0 0.3723 0 2.0 1e-06 
0.0 0.3724 0 2.0 1e-06 
0.0 0.3725 0 2.0 1e-06 
0.0 0.3726 0 2.0 1e-06 
0.0 0.3727 0 2.0 1e-06 
0.0 0.3728 0 2.0 1e-06 
0.0 0.3729 0 2.0 1e-06 
0.0 0.373 0 2.0 1e-06 
0.0 0.3731 0 2.0 1e-06 
0.0 0.3732 0 2.0 1e-06 
0.0 0.3733 0 2.0 1e-06 
0.0 0.3734 0 2.0 1e-06 
0.0 0.3735 0 2.0 1e-06 
0.0 0.3736 0 2.0 1e-06 
0.0 0.3737 0 2.0 1e-06 
0.0 0.3738 0 2.0 1e-06 
0.0 0.3739 0 2.0 1e-06 
0.0 0.374 0 2.0 1e-06 
0.0 0.3741 0 2.0 1e-06 
0.0 0.3742 0 2.0 1e-06 
0.0 0.3743 0 2.0 1e-06 
0.0 0.3744 0 2.0 1e-06 
0.0 0.3745 0 2.0 1e-06 
0.0 0.3746 0 2.0 1e-06 
0.0 0.3747 0 2.0 1e-06 
0.0 0.3748 0 2.0 1e-06 
0.0 0.3749 0 2.0 1e-06 
0.0 0.375 0 2.0 1e-06 
0.0 0.3751 0 2.0 1e-06 
0.0 0.3752 0 2.0 1e-06 
0.0 0.3753 0 2.0 1e-06 
0.0 0.3754 0 2.0 1e-06 
0.0 0.3755 0 2.0 1e-06 
0.0 0.3756 0 2.0 1e-06 
0.0 0.3757 0 2.0 1e-06 
0.0 0.3758 0 2.0 1e-06 
0.0 0.3759 0 2.0 1e-06 
0.0 0.376 0 2.0 1e-06 
0.0 0.3761 0 2.0 1e-06 
0.0 0.3762 0 2.0 1e-06 
0.0 0.3763 0 2.0 1e-06 
0.0 0.3764 0 2.0 1e-06 
0.0 0.3765 0 2.0 1e-06 
0.0 0.3766 0 2.0 1e-06 
0.0 0.3767 0 2.0 1e-06 
0.0 0.3768 0 2.0 1e-06 
0.0 0.3769 0 2.0 1e-06 
0.0 0.377 0 2.0 1e-06 
0.0 0.3771 0 2.0 1e-06 
0.0 0.3772 0 2.0 1e-06 
0.0 0.3773 0 2.0 1e-06 
0.0 0.3774 0 2.0 1e-06 
0.0 0.3775 0 2.0 1e-06 
0.0 0.3776 0 2.0 1e-06 
0.0 0.3777 0 2.0 1e-06 
0.0 0.3778 0 2.0 1e-06 
0.0 0.3779 0 2.0 1e-06 
0.0 0.378 0 2.0 1e-06 
0.0 0.3781 0 2.0 1e-06 
0.0 0.3782 0 2.0 1e-06 
0.0 0.3783 0 2.0 1e-06 
0.0 0.3784 0 2.0 1e-06 
0.0 0.3785 0 2.0 1e-06 
0.0 0.3786 0 2.0 1e-06 
0.0 0.3787 0 2.0 1e-06 
0.0 0.3788 0 2.0 1e-06 
0.0 0.3789 0 2.0 1e-06 
0.0 0.379 0 2.0 1e-06 
0.0 0.3791 0 2.0 1e-06 
0.0 0.3792 0 2.0 1e-06 
0.0 0.3793 0 2.0 1e-06 
0.0 0.3794 0 2.0 1e-06 
0.0 0.3795 0 2.0 1e-06 
0.0 0.3796 0 2.0 1e-06 
0.0 0.3797 0 2.0 1e-06 
0.0 0.3798 0 2.0 1e-06 
0.0 0.3799 0 2.0 1e-06 
0.0 0.38 0 2.0 1e-06 
0.0 0.3801 0 2.0 1e-06 
0.0 0.3802 0 2.0 1e-06 
0.0 0.3803 0 2.0 1e-06 
0.0 0.3804 0 2.0 1e-06 
0.0 0.3805 0 2.0 1e-06 
0.0 0.3806 0 2.0 1e-06 
0.0 0.3807 0 2.0 1e-06 
0.0 0.3808 0 2.0 1e-06 
0.0 0.3809 0 2.0 1e-06 
0.0 0.381 0 2.0 1e-06 
0.0 0.3811 0 2.0 1e-06 
0.0 0.3812 0 2.0 1e-06 
0.0 0.3813 0 2.0 1e-06 
0.0 0.3814 0 2.0 1e-06 
0.0 0.3815 0 2.0 1e-06 
0.0 0.3816 0 2.0 1e-06 
0.0 0.3817 0 2.0 1e-06 
0.0 0.3818 0 2.0 1e-06 
0.0 0.3819 0 2.0 1e-06 
0.0 0.382 0 2.0 1e-06 
0.0 0.3821 0 2.0 1e-06 
0.0 0.3822 0 2.0 1e-06 
0.0 0.3823 0 2.0 1e-06 
0.0 0.3824 0 2.0 1e-06 
0.0 0.3825 0 2.0 1e-06 
0.0 0.3826 0 2.0 1e-06 
0.0 0.3827 0 2.0 1e-06 
0.0 0.3828 0 2.0 1e-06 
0.0 0.3829 0 2.0 1e-06 
0.0 0.383 0 2.0 1e-06 
0.0 0.3831 0 2.0 1e-06 
0.0 0.3832 0 2.0 1e-06 
0.0 0.3833 0 2.0 1e-06 
0.0 0.3834 0 2.0 1e-06 
0.0 0.3835 0 2.0 1e-06 
0.0 0.3836 0 2.0 1e-06 
0.0 0.3837 0 2.0 1e-06 
0.0 0.3838 0 2.0 1e-06 
0.0 0.3839 0 2.0 1e-06 
0.0 0.384 0 2.0 1e-06 
0.0 0.3841 0 2.0 1e-06 
0.0 0.3842 0 2.0 1e-06 
0.0 0.3843 0 2.0 1e-06 
0.0 0.3844 0 2.0 1e-06 
0.0 0.3845 0 2.0 1e-06 
0.0 0.3846 0 2.0 1e-06 
0.0 0.3847 0 2.0 1e-06 
0.0 0.3848 0 2.0 1e-06 
0.0 0.3849 0 2.0 1e-06 
0.0 0.385 0 2.0 1e-06 
0.0 0.3851 0 2.0 1e-06 
0.0 0.3852 0 2.0 1e-06 
0.0 0.3853 0 2.0 1e-06 
0.0 0.3854 0 2.0 1e-06 
0.0 0.3855 0 2.0 1e-06 
0.0 0.3856 0 2.0 1e-06 
0.0 0.3857 0 2.0 1e-06 
0.0 0.3858 0 2.0 1e-06 
0.0 0.3859 0 2.0 1e-06 
0.0 0.386 0 2.0 1e-06 
0.0 0.3861 0 2.0 1e-06 
0.0 0.3862 0 2.0 1e-06 
0.0 0.3863 0 2.0 1e-06 
0.0 0.3864 0 2.0 1e-06 
0.0 0.3865 0 2.0 1e-06 
0.0 0.3866 0 2.0 1e-06 
0.0 0.3867 0 2.0 1e-06 
0.0 0.3868 0 2.0 1e-06 
0.0 0.3869 0 2.0 1e-06 
0.0 0.387 0 2.0 1e-06 
0.0 0.3871 0 2.0 1e-06 
0.0 0.3872 0 2.0 1e-06 
0.0 0.3873 0 2.0 1e-06 
0.0 0.3874 0 2.0 1e-06 
0.0 0.3875 0 2.0 1e-06 
0.0 0.3876 0 2.0 1e-06 
0.0 0.3877 0 2.0 1e-06 
0.0 0.3878 0 2.0 1e-06 
0.0 0.3879 0 2.0 1e-06 
0.0 0.388 0 2.0 1e-06 
0.0 0.3881 0 2.0 1e-06 
0.0 0.3882 0 2.0 1e-06 
0.0 0.3883 0 2.0 1e-06 
0.0 0.3884 0 2.0 1e-06 
0.0 0.3885 0 2.0 1e-06 
0.0 0.3886 0 2.0 1e-06 
0.0 0.3887 0 2.0 1e-06 
0.0 0.3888 0 2.0 1e-06 
0.0 0.3889 0 2.0 1e-06 
0.0 0.389 0 2.0 1e-06 
0.0 0.3891 0 2.0 1e-06 
0.0 0.3892 0 2.0 1e-06 
0.0 0.3893 0 2.0 1e-06 
0.0 0.3894 0 2.0 1e-06 
0.0 0.3895 0 2.0 1e-06 
0.0 0.3896 0 2.0 1e-06 
0.0 0.3897 0 2.0 1e-06 
0.0 0.3898 0 2.0 1e-06 
0.0 0.3899 0 2.0 1e-06 
0.0 0.39 0 2.0 1e-06 
0.0 0.3901 0 2.0 1e-06 
0.0 0.3902 0 2.0 1e-06 
0.0 0.3903 0 2.0 1e-06 
0.0 0.3904 0 2.0 1e-06 
0.0 0.3905 0 2.0 1e-06 
0.0 0.3906 0 2.0 1e-06 
0.0 0.3907 0 2.0 1e-06 
0.0 0.3908 0 2.0 1e-06 
0.0 0.3909 0 2.0 1e-06 
0.0 0.391 0 2.0 1e-06 
0.0 0.3911 0 2.0 1e-06 
0.0 0.3912 0 2.0 1e-06 
0.0 0.3913 0 2.0 1e-06 
0.0 0.3914 0 2.0 1e-06 
0.0 0.3915 0 2.0 1e-06 
0.0 0.3916 0 2.0 1e-06 
0.0 0.3917 0 2.0 1e-06 
0.0 0.3918 0 2.0 1e-06 
0.0 0.3919 0 2.0 1e-06 
0.0 0.392 0 2.0 1e-06 
0.0 0.3921 0 2.0 1e-06 
0.0 0.3922 0 2.0 1e-06 
0.0 0.3923 0 2.0 1e-06 
0.0 0.3924 0 2.0 1e-06 
0.0 0.3925 0 2.0 1e-06 
0.0 0.3926 0 2.0 1e-06 
0.0 0.3927 0 2.0 1e-06 
0.0 0.3928 0 2.0 1e-06 
0.0 0.3929 0 2.0 1e-06 
0.0 0.393 0 2.0 1e-06 
0.0 0.3931 0 2.0 1e-06 
0.0 0.3932 0 2.0 1e-06 
0.0 0.3933 0 2.0 1e-06 
0.0 0.3934 0 2.0 1e-06 
0.0 0.3935 0 2.0 1e-06 
0.0 0.3936 0 2.0 1e-06 
0.0 0.3937 0 2.0 1e-06 
0.0 0.3938 0 2.0 1e-06 
0.0 0.3939 0 2.0 1e-06 
0.0 0.394 0 2.0 1e-06 
0.0 0.3941 0 2.0 1e-06 
0.0 0.3942 0 2.0 1e-06 
0.0 0.3943 0 2.0 1e-06 
0.0 0.3944 0 2.0 1e-06 
0.0 0.3945 0 2.0 1e-06 
0.0 0.3946 0 2.0 1e-06 
0.0 0.3947 0 2.0 1e-06 
0.0 0.3948 0 2.0 1e-06 
0.0 0.3949 0 2.0 1e-06 
0.0 0.395 0 2.0 1e-06 
0.0 0.3951 0 2.0 1e-06 
0.0 0.3952 0 2.0 1e-06 
0.0 0.3953 0 2.0 1e-06 
0.0 0.3954 0 2.0 1e-06 
0.0 0.3955 0 2.0 1e-06 
0.0 0.3956 0 2.0 1e-06 
0.0 0.3957 0 2.0 1e-06 
0.0 0.3958 0 2.0 1e-06 
0.0 0.3959 0 2.0 1e-06 
0.0 0.396 0 2.0 1e-06 
0.0 0.3961 0 2.0 1e-06 
0.0 0.3962 0 2.0 1e-06 
0.0 0.3963 0 2.0 1e-06 
0.0 0.3964 0 2.0 1e-06 
0.0 0.3965 0 2.0 1e-06 
0.0 0.3966 0 2.0 1e-06 
0.0 0.3967 0 2.0 1e-06 
0.0 0.3968 0 2.0 1e-06 
0.0 0.3969 0 2.0 1e-06 
0.0 0.397 0 2.0 1e-06 
0.0 0.3971 0 2.0 1e-06 
0.0 0.3972 0 2.0 1e-06 
0.0 0.3973 0 2.0 1e-06 
0.0 0.3974 0 2.0 1e-06 
0.0 0.3975 0 2.0 1e-06 
0.0 0.3976 0 2.0 1e-06 
0.0 0.3977 0 2.0 1e-06 
0.0 0.3978 0 2.0 1e-06 
0.0 0.3979 0 2.0 1e-06 
0.0 0.398 0 2.0 1e-06 
0.0 0.3981 0 2.0 1e-06 
0.0 0.3982 0 2.0 1e-06 
0.0 0.3983 0 2.0 1e-06 
0.0 0.3984 0 2.0 1e-06 
0.0 0.3985 0 2.0 1e-06 
0.0 0.3986 0 2.0 1e-06 
0.0 0.3987 0 2.0 1e-06 
0.0 0.3988 0 2.0 1e-06 
0.0 0.3989 0 2.0 1e-06 
0.0 0.399 0 2.0 1e-06 
0.0 0.3991 0 2.0 1e-06 
0.0 0.3992 0 2.0 1e-06 
0.0 0.3993 0 2.0 1e-06 
0.0 0.3994 0 2.0 1e-06 
0.0 0.3995 0 2.0 1e-06 
0.0 0.3996 0 2.0 1e-06 
0.0 0.3997 0 2.0 1e-06 
0.0 0.3998 0 2.0 1e-06 
0.0 0.3999 0 2.0 1e-06 
0.0 0.4 0 2.0 1e-06 
0.0 0.4001 0 2.0 1e-06 
0.0 0.4002 0 2.0 1e-06 
0.0 0.4003 0 2.0 1e-06 
0.0 0.4004 0 2.0 1e-06 
0.0 0.4005 0 2.0 1e-06 
0.0 0.4006 0 2.0 1e-06 
0.0 0.4007 0 2.0 1e-06 
0.0 0.4008 0 2.0 1e-06 
0.0 0.4009 0 2.0 1e-06 
0.0 0.401 0 2.0 1e-06 
0.0 0.4011 0 2.0 1e-06 
0.0 0.4012 0 2.0 1e-06 
0.0 0.4013 0 2.0 1e-06 
0.0 0.4014 0 2.0 1e-06 
0.0 0.4015 0 2.0 1e-06 
0.0 0.4016 0 2.0 1e-06 
0.0 0.4017 0 2.0 1e-06 
0.0 0.4018 0 2.0 1e-06 
0.0 0.4019 0 2.0 1e-06 
0.0 0.402 0 2.0 1e-06 
0.0 0.4021 0 2.0 1e-06 
0.0 0.4022 0 2.0 1e-06 
0.0 0.4023 0 2.0 1e-06 
0.0 0.4024 0 2.0 1e-06 
0.0 0.4025 0 2.0 1e-06 
0.0 0.4026 0 2.0 1e-06 
0.0 0.4027 0 2.0 1e-06 
0.0 0.4028 0 2.0 1e-06 
0.0 0.4029 0 2.0 1e-06 
0.0 0.403 0 2.0 1e-06 
0.0 0.4031 0 2.0 1e-06 
0.0 0.4032 0 2.0 1e-06 
0.0 0.4033 0 2.0 1e-06 
0.0 0.4034 0 2.0 1e-06 
0.0 0.4035 0 2.0 1e-06 
0.0 0.4036 0 2.0 1e-06 
0.0 0.4037 0 2.0 1e-06 
0.0 0.4038 0 2.0 1e-06 
0.0 0.4039 0 2.0 1e-06 
0.0 0.404 0 2.0 1e-06 
0.0 0.4041 0 2.0 1e-06 
0.0 0.4042 0 2.0 1e-06 
0.0 0.4043 0 2.0 1e-06 
0.0 0.4044 0 2.0 1e-06 
0.0 0.4045 0 2.0 1e-06 
0.0 0.4046 0 2.0 1e-06 
0.0 0.4047 0 2.0 1e-06 
0.0 0.4048 0 2.0 1e-06 
0.0 0.4049 0 2.0 1e-06 
0.0 0.405 0 2.0 1e-06 
0.0 0.4051 0 2.0 1e-06 
0.0 0.4052 0 2.0 1e-06 
0.0 0.4053 0 2.0 1e-06 
0.0 0.4054 0 2.0 1e-06 
0.0 0.4055 0 2.0 1e-06 
0.0 0.4056 0 2.0 1e-06 
0.0 0.4057 0 2.0 1e-06 
0.0 0.4058 0 2.0 1e-06 
0.0 0.4059 0 2.0 1e-06 
0.0 0.406 0 2.0 1e-06 
0.0 0.4061 0 2.0 1e-06 
0.0 0.4062 0 2.0 1e-06 
0.0 0.4063 0 2.0 1e-06 
0.0 0.4064 0 2.0 1e-06 
0.0 0.4065 0 2.0 1e-06 
0.0 0.4066 0 2.0 1e-06 
0.0 0.4067 0 2.0 1e-06 
0.0 0.4068 0 2.0 1e-06 
0.0 0.4069 0 2.0 1e-06 
0.0 0.407 0 2.0 1e-06 
0.0 0.4071 0 2.0 1e-06 
0.0 0.4072 0 2.0 1e-06 
0.0 0.4073 0 2.0 1e-06 
0.0 0.4074 0 2.0 1e-06 
0.0 0.4075 0 2.0 1e-06 
0.0 0.4076 0 2.0 1e-06 
0.0 0.4077 0 2.0 1e-06 
0.0 0.4078 0 2.0 1e-06 
0.0 0.4079 0 2.0 1e-06 
0.0 0.408 0 2.0 1e-06 
0.0 0.4081 0 2.0 1e-06 
0.0 0.4082 0 2.0 1e-06 
0.0 0.4083 0 2.0 1e-06 
0.0 0.4084 0 2.0 1e-06 
0.0 0.4085 0 2.0 1e-06 
0.0 0.4086 0 2.0 1e-06 
0.0 0.4087 0 2.0 1e-06 
0.0 0.4088 0 2.0 1e-06 
0.0 0.4089 0 2.0 1e-06 
0.0 0.409 0 2.0 1e-06 
0.0 0.4091 0 2.0 1e-06 
0.0 0.4092 0 2.0 1e-06 
0.0 0.4093 0 2.0 1e-06 
0.0 0.4094 0 2.0 1e-06 
0.0 0.4095 0 2.0 1e-06 
0.0 0.4096 0 2.0 1e-06 
0.0 0.4097 0 2.0 1e-06 
0.0 0.4098 0 2.0 1e-06 
0.0 0.4099 0 2.0 1e-06 
0.0 0.41 0 2.0 1e-06 
0.0 0.4101 0 2.0 1e-06 
0.0 0.4102 0 2.0 1e-06 
0.0 0.4103 0 2.0 1e-06 
0.0 0.4104 0 2.0 1e-06 
0.0 0.4105 0 2.0 1e-06 
0.0 0.4106 0 2.0 1e-06 
0.0 0.4107 0 2.0 1e-06 
0.0 0.4108 0 2.0 1e-06 
0.0 0.4109 0 2.0 1e-06 
0.0 0.411 0 2.0 1e-06 
0.0 0.4111 0 2.0 1e-06 
0.0 0.4112 0 2.0 1e-06 
0.0 0.4113 0 2.0 1e-06 
0.0 0.4114 0 2.0 1e-06 
0.0 0.4115 0 2.0 1e-06 
0.0 0.4116 0 2.0 1e-06 
0.0 0.4117 0 2.0 1e-06 
0.0 0.4118 0 2.0 1e-06 
0.0 0.4119 0 2.0 1e-06 
0.0 0.412 0 2.0 1e-06 
0.0 0.4121 0 2.0 1e-06 
0.0 0.4122 0 2.0 1e-06 
0.0 0.4123 0 2.0 1e-06 
0.0 0.4124 0 2.0 1e-06 
0.0 0.4125 0 2.0 1e-06 
0.0 0.4126 0 2.0 1e-06 
0.0 0.4127 0 2.0 1e-06 
0.0 0.4128 0 2.0 1e-06 
0.0 0.4129 0 2.0 1e-06 
0.0 0.413 0 2.0 1e-06 
0.0 0.4131 0 2.0 1e-06 
0.0 0.4132 0 2.0 1e-06 
0.0 0.4133 0 2.0 1e-06 
0.0 0.4134 0 2.0 1e-06 
0.0 0.4135 0 2.0 1e-06 
0.0 0.4136 0 2.0 1e-06 
0.0 0.4137 0 2.0 1e-06 
0.0 0.4138 0 2.0 1e-06 
0.0 0.4139 0 2.0 1e-06 
0.0 0.414 0 2.0 1e-06 
0.0 0.4141 0 2.0 1e-06 
0.0 0.4142 0 2.0 1e-06 
0.0 0.4143 0 2.0 1e-06 
0.0 0.4144 0 2.0 1e-06 
0.0 0.4145 0 2.0 1e-06 
0.0 0.4146 0 2.0 1e-06 
0.0 0.4147 0 2.0 1e-06 
0.0 0.4148 0 2.0 1e-06 
0.0 0.4149 0 2.0 1e-06 
0.0 0.415 0 2.0 1e-06 
0.0 0.4151 0 2.0 1e-06 
0.0 0.4152 0 2.0 1e-06 
0.0 0.4153 0 2.0 1e-06 
0.0 0.4154 0 2.0 1e-06 
0.0 0.4155 0 2.0 1e-06 
0.0 0.4156 0 2.0 1e-06 
0.0 0.4157 0 2.0 1e-06 
0.0 0.4158 0 2.0 1e-06 
0.0 0.4159 0 2.0 1e-06 
0.0 0.416 0 2.0 1e-06 
0.0 0.4161 0 2.0 1e-06 
0.0 0.4162 0 2.0 1e-06 
0.0 0.4163 0 2.0 1e-06 
0.0 0.4164 0 2.0 1e-06 
0.0 0.4165 0 2.0 1e-06 
0.0 0.4166 0 2.0 1e-06 
0.0 0.4167 0 2.0 1e-06 
0.0 0.4168 0 2.0 1e-06 
0.0 0.4169 0 2.0 1e-06 
0.0 0.417 0 2.0 1e-06 
0.0 0.4171 0 2.0 1e-06 
0.0 0.4172 0 2.0 1e-06 
0.0 0.4173 0 2.0 1e-06 
0.0 0.4174 0 2.0 1e-06 
0.0 0.4175 0 2.0 1e-06 
0.0 0.4176 0 2.0 1e-06 
0.0 0.4177 0 2.0 1e-06 
0.0 0.4178 0 2.0 1e-06 
0.0 0.4179 0 2.0 1e-06 
0.0 0.418 0 2.0 1e-06 
0.0 0.4181 0 2.0 1e-06 
0.0 0.4182 0 2.0 1e-06 
0.0 0.4183 0 2.0 1e-06 
0.0 0.4184 0 2.0 1e-06 
0.0 0.4185 0 2.0 1e-06 
0.0 0.4186 0 2.0 1e-06 
0.0 0.4187 0 2.0 1e-06 
0.0 0.4188 0 2.0 1e-06 
0.0 0.4189 0 2.0 1e-06 
0.0 0.419 0 2.0 1e-06 
0.0 0.4191 0 2.0 1e-06 
0.0 0.4192 0 2.0 1e-06 
0.0 0.4193 0 2.0 1e-06 
0.0 0.4194 0 2.0 1e-06 
0.0 0.4195 0 2.0 1e-06 
0.0 0.4196 0 2.0 1e-06 
0.0 0.4197 0 2.0 1e-06 
0.0 0.4198 0 2.0 1e-06 
0.0 0.4199 0 2.0 1e-06 
0.0 0.42 0 2.0 1e-06 
0.0 0.4201 0 2.0 1e-06 
0.0 0.4202 0 2.0 1e-06 
0.0 0.4203 0 2.0 1e-06 
0.0 0.4204 0 2.0 1e-06 
0.0 0.4205 0 2.0 1e-06 
0.0 0.4206 0 2.0 1e-06 
0.0 0.4207 0 2.0 1e-06 
0.0 0.4208 0 2.0 1e-06 
0.0 0.4209 0 2.0 1e-06 
0.0 0.421 0 2.0 1e-06 
0.0 0.4211 0 2.0 1e-06 
0.0 0.4212 0 2.0 1e-06 
0.0 0.4213 0 2.0 1e-06 
0.0 0.4214 0 2.0 1e-06 
0.0 0.4215 0 2.0 1e-06 
0.0 0.4216 0 2.0 1e-06 
0.0 0.4217 0 2.0 1e-06 
0.0 0.4218 0 2.0 1e-06 
0.0 0.4219 0 2.0 1e-06 
0.0 0.422 0 2.0 1e-06 
0.0 0.4221 0 2.0 1e-06 
0.0 0.4222 0 2.0 1e-06 
0.0 0.4223 0 2.0 1e-06 
0.0 0.4224 0 2.0 1e-06 
0.0 0.4225 0 2.0 1e-06 
0.0 0.4226 0 2.0 1e-06 
0.0 0.4227 0 2.0 1e-06 
0.0 0.4228 0 2.0 1e-06 
0.0 0.4229 0 2.0 1e-06 
0.0 0.423 0 2.0 1e-06 
0.0 0.4231 0 2.0 1e-06 
0.0 0.4232 0 2.0 1e-06 
0.0 0.4233 0 2.0 1e-06 
0.0 0.4234 0 2.0 1e-06 
0.0 0.4235 0 2.0 1e-06 
0.0 0.4236 0 2.0 1e-06 
0.0 0.4237 0 2.0 1e-06 
0.0 0.4238 0 2.0 1e-06 
0.0 0.4239 0 2.0 1e-06 
0.0 0.424 0 2.0 1e-06 
0.0 0.4241 0 2.0 1e-06 
0.0 0.4242 0 2.0 1e-06 
0.0 0.4243 0 2.0 1e-06 
0.0 0.4244 0 2.0 1e-06 
0.0 0.4245 0 2.0 1e-06 
0.0 0.4246 0 2.0 1e-06 
0.0 0.4247 0 2.0 1e-06 
0.0 0.4248 0 2.0 1e-06 
0.0 0.4249 0 2.0 1e-06 
0.0 0.425 0 2.0 1e-06 
0.0 0.4251 0 2.0 1e-06 
0.0 0.4252 0 2.0 1e-06 
0.0 0.4253 0 2.0 1e-06 
0.0 0.4254 0 2.0 1e-06 
0.0 0.4255 0 2.0 1e-06 
0.0 0.4256 0 2.0 1e-06 
0.0 0.4257 0 2.0 1e-06 
0.0 0.4258 0 2.0 1e-06 
0.0 0.4259 0 2.0 1e-06 
0.0 0.426 0 2.0 1e-06 
0.0 0.4261 0 2.0 1e-06 
0.0 0.4262 0 2.0 1e-06 
0.0 0.4263 0 2.0 1e-06 
0.0 0.4264 0 2.0 1e-06 
0.0 0.4265 0 2.0 1e-06 
0.0 0.4266 0 2.0 1e-06 
0.0 0.4267 0 2.0 1e-06 
0.0 0.4268 0 2.0 1e-06 
0.0 0.4269 0 2.0 1e-06 
0.0 0.427 0 2.0 1e-06 
0.0 0.4271 0 2.0 1e-06 
0.0 0.4272 0 2.0 1e-06 
0.0 0.4273 0 2.0 1e-06 
0.0 0.4274 0 2.0 1e-06 
0.0 0.4275 0 2.0 1e-06 
0.0 0.4276 0 2.0 1e-06 
0.0 0.4277 0 2.0 1e-06 
0.0 0.4278 0 2.0 1e-06 
0.0 0.4279 0 2.0 1e-06 
0.0 0.428 0 2.0 1e-06 
0.0 0.4281 0 2.0 1e-06 
0.0 0.4282 0 2.0 1e-06 
0.0 0.4283 0 2.0 1e-06 
0.0 0.4284 0 2.0 1e-06 
0.0 0.4285 0 2.0 1e-06 
0.0 0.4286 0 2.0 1e-06 
0.0 0.4287 0 2.0 1e-06 
0.0 0.4288 0 2.0 1e-06 
0.0 0.4289 0 2.0 1e-06 
0.0 0.429 0 2.0 1e-06 
0.0 0.4291 0 2.0 1e-06 
0.0 0.4292 0 2.0 1e-06 
0.0 0.4293 0 2.0 1e-06 
0.0 0.4294 0 2.0 1e-06 
0.0 0.4295 0 2.0 1e-06 
0.0 0.4296 0 2.0 1e-06 
0.0 0.4297 0 2.0 1e-06 
0.0 0.4298 0 2.0 1e-06 
0.0 0.4299 0 2.0 1e-06 
0.0 0.43 0 2.0 1e-06 
0.0 0.4301 0 2.0 1e-06 
0.0 0.4302 0 2.0 1e-06 
0.0 0.4303 0 2.0 1e-06 
0.0 0.4304 0 2.0 1e-06 
0.0 0.4305 0 2.0 1e-06 
0.0 0.4306 0 2.0 1e-06 
0.0 0.4307 0 2.0 1e-06 
0.0 0.4308 0 2.0 1e-06 
0.0 0.4309 0 2.0 1e-06 
0.0 0.431 0 2.0 1e-06 
0.0 0.4311 0 2.0 1e-06 
0.0 0.4312 0 2.0 1e-06 
0.0 0.4313 0 2.0 1e-06 
0.0 0.4314 0 2.0 1e-06 
0.0 0.4315 0 2.0 1e-06 
0.0 0.4316 0 2.0 1e-06 
0.0 0.4317 0 2.0 1e-06 
0.0 0.4318 0 2.0 1e-06 
0.0 0.4319 0 2.0 1e-06 
0.0 0.432 0 2.0 1e-06 
0.0 0.4321 0 2.0 1e-06 
0.0 0.4322 0 2.0 1e-06 
0.0 0.4323 0 2.0 1e-06 
0.0 0.4324 0 2.0 1e-06 
0.0 0.4325 0 2.0 1e-06 
0.0 0.4326 0 2.0 1e-06 
0.0 0.4327 0 2.0 1e-06 
0.0 0.4328 0 2.0 1e-06 
0.0 0.4329 0 2.0 1e-06 
0.0 0.433 0 2.0 1e-06 
0.0 0.4331 0 2.0 1e-06 
0.0 0.4332 0 2.0 1e-06 
0.0 0.4333 0 2.0 1e-06 
0.0 0.4334 0 2.0 1e-06 
0.0 0.4335 0 2.0 1e-06 
0.0 0.4336 0 2.0 1e-06 
0.0 0.4337 0 2.0 1e-06 
0.0 0.4338 0 2.0 1e-06 
0.0 0.4339 0 2.0 1e-06 
0.0 0.434 0 2.0 1e-06 
0.0 0.4341 0 2.0 1e-06 
0.0 0.4342 0 2.0 1e-06 
0.0 0.4343 0 2.0 1e-06 
0.0 0.4344 0 2.0 1e-06 
0.0 0.4345 0 2.0 1e-06 
0.0 0.4346 0 2.0 1e-06 
0.0 0.4347 0 2.0 1e-06 
0.0 0.4348 0 2.0 1e-06 
0.0 0.4349 0 2.0 1e-06 
0.0 0.435 0 2.0 1e-06 
0.0 0.4351 0 2.0 1e-06 
0.0 0.4352 0 2.0 1e-06 
0.0 0.4353 0 2.0 1e-06 
0.0 0.4354 0 2.0 1e-06 
0.0 0.4355 0 2.0 1e-06 
0.0 0.4356 0 2.0 1e-06 
0.0 0.4357 0 2.0 1e-06 
0.0 0.4358 0 2.0 1e-06 
0.0 0.4359 0 2.0 1e-06 
0.0 0.436 0 2.0 1e-06 
0.0 0.4361 0 2.0 1e-06 
0.0 0.4362 0 2.0 1e-06 
0.0 0.4363 0 2.0 1e-06 
0.0 0.4364 0 2.0 1e-06 
0.0 0.4365 0 2.0 1e-06 
0.0 0.4366 0 2.0 1e-06 
0.0 0.4367 0 2.0 1e-06 
0.0 0.4368 0 2.0 1e-06 
0.0 0.4369 0 2.0 1e-06 
0.0 0.437 0 2.0 1e-06 
0.0 0.4371 0 2.0 1e-06 
0.0 0.4372 0 2.0 1e-06 
0.0 0.4373 0 2.0 1e-06 
0.0 0.4374 0 2.0 1e-06 
0.0 0.4375 0 2.0 1e-06 
0.0 0.4376 0 2.0 1e-06 
0.0 0.4377 0 2.0 1e-06 
0.0 0.4378 0 2.0 1e-06 
0.0 0.4379 0 2.0 1e-06 
0.0 0.438 0 2.0 1e-06 
0.0 0.4381 0 2.0 1e-06 
0.0 0.4382 0 2.0 1e-06 
0.0 0.4383 0 2.0 1e-06 
0.0 0.4384 0 2.0 1e-06 
0.0 0.4385 0 2.0 1e-06 
0.0 0.4386 0 2.0 1e-06 
0.0 0.4387 0 2.0 1e-06 
0.0 0.4388 0 2.0 1e-06 
0.0 0.4389 0 2.0 1e-06 
0.0 0.439 0 2.0 1e-06 
0.0 0.4391 0 2.0 1e-06 
0.0 0.4392 0 2.0 1e-06 
0.0 0.4393 0 2.0 1e-06 
0.0 0.4394 0 2.0 1e-06 
0.0 0.4395 0 2.0 1e-06 
0.0 0.4396 0 2.0 1e-06 
0.0 0.4397 0 2.0 1e-06 
0.0 0.4398 0 2.0 1e-06 
0.0 0.4399 0 2.0 1e-06 
0.0 0.44 0 2.0 1e-06 
0.0 0.4401 0 2.0 1e-06 
0.0 0.4402 0 2.0 1e-06 
0.0 0.4403 0 2.0 1e-06 
0.0 0.4404 0 2.0 1e-06 
0.0 0.4405 0 2.0 1e-06 
0.0 0.4406 0 2.0 1e-06 
0.0 0.4407 0 2.0 1e-06 
0.0 0.4408 0 2.0 1e-06 
0.0 0.4409 0 2.0 1e-06 
0.0 0.441 0 2.0 1e-06 
0.0 0.4411 0 2.0 1e-06 
0.0 0.4412 0 2.0 1e-06 
0.0 0.4413 0 2.0 1e-06 
0.0 0.4414 0 2.0 1e-06 
0.0 0.4415 0 2.0 1e-06 
0.0 0.4416 0 2.0 1e-06 
0.0 0.4417 0 2.0 1e-06 
0.0 0.4418 0 2.0 1e-06 
0.0 0.4419 0 2.0 1e-06 
0.0 0.442 0 2.0 1e-06 
0.0 0.4421 0 2.0 1e-06 
0.0 0.4422 0 2.0 1e-06 
0.0 0.4423 0 2.0 1e-06 
0.0 0.4424 0 2.0 1e-06 
0.0 0.4425 0 2.0 1e-06 
0.0 0.4426 0 2.0 1e-06 
0.0 0.4427 0 2.0 1e-06 
0.0 0.4428 0 2.0 1e-06 
0.0 0.4429 0 2.0 1e-06 
0.0 0.443 0 2.0 1e-06 
0.0 0.4431 0 2.0 1e-06 
0.0 0.4432 0 2.0 1e-06 
0.0 0.4433 0 2.0 1e-06 
0.0 0.4434 0 2.0 1e-06 
0.0 0.4435 0 2.0 1e-06 
0.0 0.4436 0 2.0 1e-06 
0.0 0.4437 0 2.0 1e-06 
0.0 0.4438 0 2.0 1e-06 
0.0 0.4439 0 2.0 1e-06 
0.0 0.444 0 2.0 1e-06 
0.0 0.4441 0 2.0 1e-06 
0.0 0.4442 0 2.0 1e-06 
0.0 0.4443 0 2.0 1e-06 
0.0 0.4444 0 2.0 1e-06 
0.0 0.4445 0 2.0 1e-06 
0.0 0.4446 0 2.0 1e-06 
0.0 0.4447 0 2.0 1e-06 
0.0 0.4448 0 2.0 1e-06 
0.0 0.4449 0 2.0 1e-06 
0.0 0.445 0 2.0 1e-06 
0.0 0.4451 0 2.0 1e-06 
0.0 0.4452 0 2.0 1e-06 
0.0 0.4453 0 2.0 1e-06 
0.0 0.4454 0 2.0 1e-06 
0.0 0.4455 0 2.0 1e-06 
0.0 0.4456 0 2.0 1e-06 
0.0 0.4457 0 2.0 1e-06 
0.0 0.4458 0 2.0 1e-06 
0.0 0.4459 0 2.0 1e-06 
0.0 0.446 0 2.0 1e-06 
0.0 0.4461 0 2.0 1e-06 
0.0 0.4462 0 2.0 1e-06 
0.0 0.4463 0 2.0 1e-06 
0.0 0.4464 0 2.0 1e-06 
0.0 0.4465 0 2.0 1e-06 
0.0 0.4466 0 2.0 1e-06 
0.0 0.4467 0 2.0 1e-06 
0.0 0.4468 0 2.0 1e-06 
0.0 0.4469 0 2.0 1e-06 
0.0 0.447 0 2.0 1e-06 
0.0 0.4471 0 2.0 1e-06 
0.0 0.4472 0 2.0 1e-06 
0.0 0.4473 0 2.0 1e-06 
0.0 0.4474 0 2.0 1e-06 
0.0 0.4475 0 2.0 1e-06 
0.0 0.4476 0 2.0 1e-06 
0.0 0.4477 0 2.0 1e-06 
0.0 0.4478 0 2.0 1e-06 
0.0 0.4479 0 2.0 1e-06 
0.0 0.448 0 2.0 1e-06 
0.0 0.4481 0 2.0 1e-06 
0.0 0.4482 0 2.0 1e-06 
0.0 0.4483 0 2.0 1e-06 
0.0 0.4484 0 2.0 1e-06 
0.0 0.4485 0 2.0 1e-06 
0.0 0.4486 0 2.0 1e-06 
0.0 0.4487 0 2.0 1e-06 
0.0 0.4488 0 2.0 1e-06 
0.0 0.4489 0 2.0 1e-06 
0.0 0.449 0 2.0 1e-06 
0.0 0.4491 0 2.0 1e-06 
0.0 0.4492 0 2.0 1e-06 
0.0 0.4493 0 2.0 1e-06 
0.0 0.4494 0 2.0 1e-06 
0.0 0.4495 0 2.0 1e-06 
0.0 0.4496 0 2.0 1e-06 
0.0 0.4497 0 2.0 1e-06 
0.0 0.4498 0 2.0 1e-06 
0.0 0.4499 0 2.0 1e-06 
0.0 0.45 0 2.0 1e-06 
0.0 0.4501 0 2.0 1e-06 
0.0 0.4502 0 2.0 1e-06 
0.0 0.4503 0 2.0 1e-06 
0.0 0.4504 0 2.0 1e-06 
0.0 0.4505 0 2.0 1e-06 
0.0 0.4506 0 2.0 1e-06 
0.0 0.4507 0 2.0 1e-06 
0.0 0.4508 0 2.0 1e-06 
0.0 0.4509 0 2.0 1e-06 
0.0 0.451 0 2.0 1e-06 
0.0 0.4511 0 2.0 1e-06 
0.0 0.4512 0 2.0 1e-06 
0.0 0.4513 0 2.0 1e-06 
0.0 0.4514 0 2.0 1e-06 
0.0 0.4515 0 2.0 1e-06 
0.0 0.4516 0 2.0 1e-06 
0.0 0.4517 0 2.0 1e-06 
0.0 0.4518 0 2.0 1e-06 
0.0 0.4519 0 2.0 1e-06 
0.0 0.452 0 2.0 1e-06 
0.0 0.4521 0 2.0 1e-06 
0.0 0.4522 0 2.0 1e-06 
0.0 0.4523 0 2.0 1e-06 
0.0 0.4524 0 2.0 1e-06 
0.0 0.4525 0 2.0 1e-06 
0.0 0.4526 0 2.0 1e-06 
0.0 0.4527 0 2.0 1e-06 
0.0 0.4528 0 2.0 1e-06 
0.0 0.4529 0 2.0 1e-06 
0.0 0.453 0 2.0 1e-06 
0.0 0.4531 0 2.0 1e-06 
0.0 0.4532 0 2.0 1e-06 
0.0 0.4533 0 2.0 1e-06 
0.0 0.4534 0 2.0 1e-06 
0.0 0.4535 0 2.0 1e-06 
0.0 0.4536 0 2.0 1e-06 
0.0 0.4537 0 2.0 1e-06 
0.0 0.4538 0 2.0 1e-06 
0.0 0.4539 0 2.0 1e-06 
0.0 0.454 0 2.0 1e-06 
0.0 0.4541 0 2.0 1e-06 
0.0 0.4542 0 2.0 1e-06 
0.0 0.4543 0 2.0 1e-06 
0.0 0.4544 0 2.0 1e-06 
0.0 0.4545 0 2.0 1e-06 
0.0 0.4546 0 2.0 1e-06 
0.0 0.4547 0 2.0 1e-06 
0.0 0.4548 0 2.0 1e-06 
0.0 0.4549 0 2.0 1e-06 
0.0 0.455 0 2.0 1e-06 
0.0 0.4551 0 2.0 1e-06 
0.0 0.4552 0 2.0 1e-06 
0.0 0.4553 0 2.0 1e-06 
0.0 0.4554 0 2.0 1e-06 
0.0 0.4555 0 2.0 1e-06 
0.0 0.4556 0 2.0 1e-06 
0.0 0.4557 0 2.0 1e-06 
0.0 0.4558 0 2.0 1e-06 
0.0 0.4559 0 2.0 1e-06 
0.0 0.456 0 2.0 1e-06 
0.0 0.4561 0 2.0 1e-06 
0.0 0.4562 0 2.0 1e-06 
0.0 0.4563 0 2.0 1e-06 
0.0 0.4564 0 2.0 1e-06 
0.0 0.4565 0 2.0 1e-06 
0.0 0.4566 0 2.0 1e-06 
0.0 0.4567 0 2.0 1e-06 
0.0 0.4568 0 2.0 1e-06 
0.0 0.4569 0 2.0 1e-06 
0.0 0.457 0 2.0 1e-06 
0.0 0.4571 0 2.0 1e-06 
0.0 0.4572 0 2.0 1e-06 
0.0 0.4573 0 2.0 1e-06 
0.0 0.4574 0 2.0 1e-06 
0.0 0.4575 0 2.0 1e-06 
0.0 0.4576 0 2.0 1e-06 
0.0 0.4577 0 2.0 1e-06 
0.0 0.4578 0 2.0 1e-06 
0.0 0.4579 0 2.0 1e-06 
0.0 0.458 0 2.0 1e-06 
0.0 0.4581 0 2.0 1e-06 
0.0 0.4582 0 2.0 1e-06 
0.0 0.4583 0 2.0 1e-06 
0.0 0.4584 0 2.0 1e-06 
0.0 0.4585 0 2.0 1e-06 
0.0 0.4586 0 2.0 1e-06 
0.0 0.4587 0 2.0 1e-06 
0.0 0.4588 0 2.0 1e-06 
0.0 0.4589 0 2.0 1e-06 
0.0 0.459 0 2.0 1e-06 
0.0 0.4591 0 2.0 1e-06 
0.0 0.4592 0 2.0 1e-06 
0.0 0.4593 0 2.0 1e-06 
0.0 0.4594 0 2.0 1e-06 
0.0 0.4595 0 2.0 1e-06 
0.0 0.4596 0 2.0 1e-06 
0.0 0.4597 0 2.0 1e-06 
0.0 0.4598 0 2.0 1e-06 
0.0 0.4599 0 2.0 1e-06 
0.0 0.46 0 2.0 1e-06 
0.0 0.4601 0 2.0 1e-06 
0.0 0.4602 0 2.0 1e-06 
0.0 0.4603 0 2.0 1e-06 
0.0 0.4604 0 2.0 1e-06 
0.0 0.4605 0 2.0 1e-06 
0.0 0.4606 0 2.0 1e-06 
0.0 0.4607 0 2.0 1e-06 
0.0 0.4608 0 2.0 1e-06 
0.0 0.4609 0 2.0 1e-06 
0.0 0.461 0 2.0 1e-06 
0.0 0.4611 0 2.0 1e-06 
0.0 0.4612 0 2.0 1e-06 
0.0 0.4613 0 2.0 1e-06 
0.0 0.4614 0 2.0 1e-06 
0.0 0.4615 0 2.0 1e-06 
0.0 0.4616 0 2.0 1e-06 
0.0 0.4617 0 2.0 1e-06 
0.0 0.4618 0 2.0 1e-06 
0.0 0.4619 0 2.0 1e-06 
0.0 0.462 0 2.0 1e-06 
0.0 0.4621 0 2.0 1e-06 
0.0 0.4622 0 2.0 1e-06 
0.0 0.4623 0 2.0 1e-06 
0.0 0.4624 0 2.0 1e-06 
0.0 0.4625 0 2.0 1e-06 
0.0 0.4626 0 2.0 1e-06 
0.0 0.4627 0 2.0 1e-06 
0.0 0.4628 0 2.0 1e-06 
0.0 0.4629 0 2.0 1e-06 
0.0 0.463 0 2.0 1e-06 
0.0 0.4631 0 2.0 1e-06 
0.0 0.4632 0 2.0 1e-06 
0.0 0.4633 0 2.0 1e-06 
0.0 0.4634 0 2.0 1e-06 
0.0 0.4635 0 2.0 1e-06 
0.0 0.4636 0 2.0 1e-06 
0.0 0.4637 0 2.0 1e-06 
0.0 0.4638 0 2.0 1e-06 
0.0 0.4639 0 2.0 1e-06 
0.0 0.464 0 2.0 1e-06 
0.0 0.4641 0 2.0 1e-06 
0.0 0.4642 0 2.0 1e-06 
0.0 0.4643 0 2.0 1e-06 
0.0 0.4644 0 2.0 1e-06 
0.0 0.4645 0 2.0 1e-06 
0.0 0.4646 0 2.0 1e-06 
0.0 0.4647 0 2.0 1e-06 
0.0 0.4648 0 2.0 1e-06 
0.0 0.4649 0 2.0 1e-06 
0.0 0.465 0 2.0 1e-06 
0.0 0.4651 0 2.0 1e-06 
0.0 0.4652 0 2.0 1e-06 
0.0 0.4653 0 2.0 1e-06 
0.0 0.4654 0 2.0 1e-06 
0.0 0.4655 0 2.0 1e-06 
0.0 0.4656 0 2.0 1e-06 
0.0 0.4657 0 2.0 1e-06 
0.0 0.4658 0 2.0 1e-06 
0.0 0.4659 0 2.0 1e-06 
0.0 0.466 0 2.0 1e-06 
0.0 0.4661 0 2.0 1e-06 
0.0 0.4662 0 2.0 1e-06 
0.0 0.4663 0 2.0 1e-06 
0.0 0.4664 0 2.0 1e-06 
0.0 0.4665 0 2.0 1e-06 
0.0 0.4666 0 2.0 1e-06 
0.0 0.4667 0 2.0 1e-06 
0.0 0.4668 0 2.0 1e-06 
0.0 0.4669 0 2.0 1e-06 
0.0 0.467 0 2.0 1e-06 
0.0 0.4671 0 2.0 1e-06 
0.0 0.4672 0 2.0 1e-06 
0.0 0.4673 0 2.0 1e-06 
0.0 0.4674 0 2.0 1e-06 
0.0 0.4675 0 2.0 1e-06 
0.0 0.4676 0 2.0 1e-06 
0.0 0.4677 0 2.0 1e-06 
0.0 0.4678 0 2.0 1e-06 
0.0 0.4679 0 2.0 1e-06 
0.0 0.468 0 2.0 1e-06 
0.0 0.4681 0 2.0 1e-06 
0.0 0.4682 0 2.0 1e-06 
0.0 0.4683 0 2.0 1e-06 
0.0 0.4684 0 2.0 1e-06 
0.0 0.4685 0 2.0 1e-06 
0.0 0.4686 0 2.0 1e-06 
0.0 0.4687 0 2.0 1e-06 
0.0 0.4688 0 2.0 1e-06 
0.0 0.4689 0 2.0 1e-06 
0.0 0.469 0 2.0 1e-06 
0.0 0.4691 0 2.0 1e-06 
0.0 0.4692 0 2.0 1e-06 
0.0 0.4693 0 2.0 1e-06 
0.0 0.4694 0 2.0 1e-06 
0.0 0.4695 0 2.0 1e-06 
0.0 0.4696 0 2.0 1e-06 
0.0 0.4697 0 2.0 1e-06 
0.0 0.4698 0 2.0 1e-06 
0.0 0.4699 0 2.0 1e-06 
0.0 0.47 0 2.0 1e-06 
0.0 0.4701 0 2.0 1e-06 
0.0 0.4702 0 2.0 1e-06 
0.0 0.4703 0 2.0 1e-06 
0.0 0.4704 0 2.0 1e-06 
0.0 0.4705 0 2.0 1e-06 
0.0 0.4706 0 2.0 1e-06 
0.0 0.4707 0 2.0 1e-06 
0.0 0.4708 0 2.0 1e-06 
0.0 0.4709 0 2.0 1e-06 
0.0 0.471 0 2.0 1e-06 
0.0 0.4711 0 2.0 1e-06 
0.0 0.4712 0 2.0 1e-06 
0.0 0.4713 0 2.0 1e-06 
0.0 0.4714 0 2.0 1e-06 
0.0 0.4715 0 2.0 1e-06 
0.0 0.4716 0 2.0 1e-06 
0.0 0.4717 0 2.0 1e-06 
0.0 0.4718 0 2.0 1e-06 
0.0 0.4719 0 2.0 1e-06 
0.0 0.472 0 2.0 1e-06 
0.0 0.4721 0 2.0 1e-06 
0.0 0.4722 0 2.0 1e-06 
0.0 0.4723 0 2.0 1e-06 
0.0 0.4724 0 2.0 1e-06 
0.0 0.4725 0 2.0 1e-06 
0.0 0.4726 0 2.0 1e-06 
0.0 0.4727 0 2.0 1e-06 
0.0 0.4728 0 2.0 1e-06 
0.0 0.4729 0 2.0 1e-06 
0.0 0.473 0 2.0 1e-06 
0.0 0.4731 0 2.0 1e-06 
0.0 0.4732 0 2.0 1e-06 
0.0 0.4733 0 2.0 1e-06 
0.0 0.4734 0 2.0 1e-06 
0.0 0.4735 0 2.0 1e-06 
0.0 0.4736 0 2.0 1e-06 
0.0 0.4737 0 2.0 1e-06 
0.0 0.4738 0 2.0 1e-06 
0.0 0.4739 0 2.0 1e-06 
0.0 0.474 0 2.0 1e-06 
0.0 0.4741 0 2.0 1e-06 
0.0 0.4742 0 2.0 1e-06 
0.0 0.4743 0 2.0 1e-06 
0.0 0.4744 0 2.0 1e-06 
0.0 0.4745 0 2.0 1e-06 
0.0 0.4746 0 2.0 1e-06 
0.0 0.4747 0 2.0 1e-06 
0.0 0.4748 0 2.0 1e-06 
0.0 0.4749 0 2.0 1e-06 
0.0 0.475 0 2.0 1e-06 
0.0 0.4751 0 2.0 1e-06 
0.0 0.4752 0 2.0 1e-06 
0.0 0.4753 0 2.0 1e-06 
0.0 0.4754 0 2.0 1e-06 
0.0 0.4755 0 2.0 1e-06 
0.0 0.4756 0 2.0 1e-06 
0.0 0.4757 0 2.0 1e-06 
0.0 0.4758 0 2.0 1e-06 
0.0 0.4759 0 2.0 1e-06 
0.0 0.476 0 2.0 1e-06 
0.0 0.4761 0 2.0 1e-06 
0.0 0.4762 0 2.0 1e-06 
0.0 0.4763 0 2.0 1e-06 
0.0 0.4764 0 2.0 1e-06 
0.0 0.4765 0 2.0 1e-06 
0.0 0.4766 0 2.0 1e-06 
0.0 0.4767 0 2.0 1e-06 
0.0 0.4768 0 2.0 1e-06 
0.0 0.4769 0 2.0 1e-06 
0.0 0.477 0 2.0 1e-06 
0.0 0.4771 0 2.0 1e-06 
0.0 0.4772 0 2.0 1e-06 
0.0 0.4773 0 2.0 1e-06 
0.0 0.4774 0 2.0 1e-06 
0.0 0.4775 0 2.0 1e-06 
0.0 0.4776 0 2.0 1e-06 
0.0 0.4777 0 2.0 1e-06 
0.0 0.4778 0 2.0 1e-06 
0.0 0.4779 0 2.0 1e-06 
0.0 0.478 0 2.0 1e-06 
0.0 0.4781 0 2.0 1e-06 
0.0 0.4782 0 2.0 1e-06 
0.0 0.4783 0 2.0 1e-06 
0.0 0.4784 0 2.0 1e-06 
0.0 0.4785 0 2.0 1e-06 
0.0 0.4786 0 2.0 1e-06 
0.0 0.4787 0 2.0 1e-06 
0.0 0.4788 0 2.0 1e-06 
0.0 0.4789 0 2.0 1e-06 
0.0 0.479 0 2.0 1e-06 
0.0 0.4791 0 2.0 1e-06 
0.0 0.4792 0 2.0 1e-06 
0.0 0.4793 0 2.0 1e-06 
0.0 0.4794 0 2.0 1e-06 
0.0 0.4795 0 2.0 1e-06 
0.0 0.4796 0 2.0 1e-06 
0.0 0.4797 0 2.0 1e-06 
0.0 0.4798 0 2.0 1e-06 
0.0 0.4799 0 2.0 1e-06 
0.0 0.48 0 2.0 1e-06 
0.0 0.4801 0 2.0 1e-06 
0.0 0.4802 0 2.0 1e-06 
0.0 0.4803 0 2.0 1e-06 
0.0 0.4804 0 2.0 1e-06 
0.0 0.4805 0 2.0 1e-06 
0.0 0.4806 0 2.0 1e-06 
0.0 0.4807 0 2.0 1e-06 
0.0 0.4808 0 2.0 1e-06 
0.0 0.4809 0 2.0 1e-06 
0.0 0.481 0 2.0 1e-06 
0.0 0.4811 0 2.0 1e-06 
0.0 0.4812 0 2.0 1e-06 
0.0 0.4813 0 2.0 1e-06 
0.0 0.4814 0 2.0 1e-06 
0.0 0.4815 0 2.0 1e-06 
0.0 0.4816 0 2.0 1e-06 
0.0 0.4817 0 2.0 1e-06 
0.0 0.4818 0 2.0 1e-06 
0.0 0.4819 0 2.0 1e-06 
0.0 0.482 0 2.0 1e-06 
0.0 0.4821 0 2.0 1e-06 
0.0 0.4822 0 2.0 1e-06 
0.0 0.4823 0 2.0 1e-06 
0.0 0.4824 0 2.0 1e-06 
0.0 0.4825 0 2.0 1e-06 
0.0 0.4826 0 2.0 1e-06 
0.0 0.4827 0 2.0 1e-06 
0.0 0.4828 0 2.0 1e-06 
0.0 0.4829 0 2.0 1e-06 
0.0 0.483 0 2.0 1e-06 
0.0 0.4831 0 2.0 1e-06 
0.0 0.4832 0 2.0 1e-06 
0.0 0.4833 0 2.0 1e-06 
0.0 0.4834 0 2.0 1e-06 
0.0 0.4835 0 2.0 1e-06 
0.0 0.4836 0 2.0 1e-06 
0.0 0.4837 0 2.0 1e-06 
0.0 0.4838 0 2.0 1e-06 
0.0 0.4839 0 2.0 1e-06 
0.0 0.484 0 2.0 1e-06 
0.0 0.4841 0 2.0 1e-06 
0.0 0.4842 0 2.0 1e-06 
0.0 0.4843 0 2.0 1e-06 
0.0 0.4844 0 2.0 1e-06 
0.0 0.4845 0 2.0 1e-06 
0.0 0.4846 0 2.0 1e-06 
0.0 0.4847 0 2.0 1e-06 
0.0 0.4848 0 2.0 1e-06 
0.0 0.4849 0 2.0 1e-06 
0.0 0.485 0 2.0 1e-06 
0.0 0.4851 0 2.0 1e-06 
0.0 0.4852 0 2.0 1e-06 
0.0 0.4853 0 2.0 1e-06 
0.0 0.4854 0 2.0 1e-06 
0.0 0.4855 0 2.0 1e-06 
0.0 0.4856 0 2.0 1e-06 
0.0 0.4857 0 2.0 1e-06 
0.0 0.4858 0 2.0 1e-06 
0.0 0.4859 0 2.0 1e-06 
0.0 0.486 0 2.0 1e-06 
0.0 0.4861 0 2.0 1e-06 
0.0 0.4862 0 2.0 1e-06 
0.0 0.4863 0 2.0 1e-06 
0.0 0.4864 0 2.0 1e-06 
0.0 0.4865 0 2.0 1e-06 
0.0 0.4866 0 2.0 1e-06 
0.0 0.4867 0 2.0 1e-06 
0.0 0.4868 0 2.0 1e-06 
0.0 0.4869 0 2.0 1e-06 
0.0 0.487 0 2.0 1e-06 
0.0 0.4871 0 2.0 1e-06 
0.0 0.4872 0 2.0 1e-06 
0.0 0.4873 0 2.0 1e-06 
0.0 0.4874 0 2.0 1e-06 
0.0 0.4875 0 2.0 1e-06 
0.0 0.4876 0 2.0 1e-06 
0.0 0.4877 0 2.0 1e-06 
0.0 0.4878 0 2.0 1e-06 
0.0 0.4879 0 2.0 1e-06 
0.0 0.488 0 2.0 1e-06 
0.0 0.4881 0 2.0 1e-06 
0.0 0.4882 0 2.0 1e-06 
0.0 0.4883 0 2.0 1e-06 
0.0 0.4884 0 2.0 1e-06 
0.0 0.4885 0 2.0 1e-06 
0.0 0.4886 0 2.0 1e-06 
0.0 0.4887 0 2.0 1e-06 
0.0 0.4888 0 2.0 1e-06 
0.0 0.4889 0 2.0 1e-06 
0.0 0.489 0 2.0 1e-06 
0.0 0.4891 0 2.0 1e-06 
0.0 0.4892 0 2.0 1e-06 
0.0 0.4893 0 2.0 1e-06 
0.0 0.4894 0 2.0 1e-06 
0.0 0.4895 0 2.0 1e-06 
0.0 0.4896 0 2.0 1e-06 
0.0 0.4897 0 2.0 1e-06 
0.0 0.4898 0 2.0 1e-06 
0.0 0.4899 0 2.0 1e-06 
0.0 0.49 0 2.0 1e-06 
0.0 0.4901 0 2.0 1e-06 
0.0 0.4902 0 2.0 1e-06 
0.0 0.4903 0 2.0 1e-06 
0.0 0.4904 0 2.0 1e-06 
0.0 0.4905 0 2.0 1e-06 
0.0 0.4906 0 2.0 1e-06 
0.0 0.4907 0 2.0 1e-06 
0.0 0.4908 0 2.0 1e-06 
0.0 0.4909 0 2.0 1e-06 
0.0 0.491 0 2.0 1e-06 
0.0 0.4911 0 2.0 1e-06 
0.0 0.4912 0 2.0 1e-06 
0.0 0.4913 0 2.0 1e-06 
0.0 0.4914 0 2.0 1e-06 
0.0 0.4915 0 2.0 1e-06 
0.0 0.4916 0 2.0 1e-06 
0.0 0.4917 0 2.0 1e-06 
0.0 0.4918 0 2.0 1e-06 
0.0 0.4919 0 2.0 1e-06 
0.0 0.492 0 2.0 1e-06 
0.0 0.4921 0 2.0 1e-06 
0.0 0.4922 0 2.0 1e-06 
0.0 0.4923 0 2.0 1e-06 
0.0 0.4924 0 2.0 1e-06 
0.0 0.4925 0 2.0 1e-06 
0.0 0.4926 0 2.0 1e-06 
0.0 0.4927 0 2.0 1e-06 
0.0 0.4928 0 2.0 1e-06 
0.0 0.4929 0 2.0 1e-06 
0.0 0.493 0 2.0 1e-06 
0.0 0.4931 0 2.0 1e-06 
0.0 0.4932 0 2.0 1e-06 
0.0 0.4933 0 2.0 1e-06 
0.0 0.4934 0 2.0 1e-06 
0.0 0.4935 0 2.0 1e-06 
0.0 0.4936 0 2.0 1e-06 
0.0 0.4937 0 2.0 1e-06 
0.0 0.4938 0 2.0 1e-06 
0.0 0.4939 0 2.0 1e-06 
0.0 0.494 0 2.0 1e-06 
0.0 0.4941 0 2.0 1e-06 
0.0 0.4942 0 2.0 1e-06 
0.0 0.4943 0 2.0 1e-06 
0.0 0.4944 0 2.0 1e-06 
0.0 0.4945 0 2.0 1e-06 
0.0 0.4946 0 2.0 1e-06 
0.0 0.4947 0 2.0 1e-06 
0.0 0.4948 0 2.0 1e-06 
0.0 0.4949 0 2.0 1e-06 
0.0 0.495 0 2.0 1e-06 
0.0 0.4951 0 2.0 1e-06 
0.0 0.4952 0 2.0 1e-06 
0.0 0.4953 0 2.0 1e-06 
0.0 0.4954 0 2.0 1e-06 
0.0 0.4955 0 2.0 1e-06 
0.0 0.4956 0 2.0 1e-06 
0.0 0.4957 0 2.0 1e-06 
0.0 0.4958 0 2.0 1e-06 
0.0 0.4959 0 2.0 1e-06 
0.0 0.496 0 2.0 1e-06 
0.0 0.4961 0 2.0 1e-06 
0.0 0.4962 0 2.0 1e-06 
0.0 0.4963 0 2.0 1e-06 
0.0 0.4964 0 2.0 1e-06 
0.0 0.4965 0 2.0 1e-06 
0.0 0.4966 0 2.0 1e-06 
0.0 0.4967 0 2.0 1e-06 
0.0 0.4968 0 2.0 1e-06 
0.0 0.4969 0 2.0 1e-06 
0.0 0.497 0 2.0 1e-06 
0.0 0.4971 0 2.0 1e-06 
0.0 0.4972 0 2.0 1e-06 
0.0 0.4973 0 2.0 1e-06 
0.0 0.4974 0 2.0 1e-06 
0.0 0.4975 0 2.0 1e-06 
0.0 0.4976 0 2.0 1e-06 
0.0 0.4977 0 2.0 1e-06 
0.0 0.4978 0 2.0 1e-06 
0.0 0.4979 0 2.0 1e-06 
0.0 0.498 0 2.0 1e-06 
0.0 0.4981 0 2.0 1e-06 
0.0 0.4982 0 2.0 1e-06 
0.0 0.4983 0 2.0 1e-06 
0.0 0.4984 0 2.0 1e-06 
0.0 0.4985 0 2.0 1e-06 
0.0 0.4986 0 2.0 1e-06 
0.0 0.4987 0 2.0 1e-06 
0.0 0.4988 0 2.0 1e-06 
0.0 0.4989 0 2.0 1e-06 
0.0 0.499 0 2.0 1e-06 
0.0 0.4991 0 2.0 1e-06 
0.0 0.4992 0 2.0 1e-06 
0.0 0.4993 0 2.0 1e-06 
0.0 0.4994 0 2.0 1e-06 
0.0 0.4995 0 2.0 1e-06 
0.0 0.4996 0 2.0 1e-06 
0.0 0.4997 0 2.0 1e-06 
0.0 0.4998 0 2.0 1e-06 
0.0 0.4999 0 2.0 1e-06 
0.0 0.5 0 2.0 1e-06 
0.0 0.5001 0 2.0 1e-06 
0.0 0.5002 0 2.0 1e-06 
0.0 0.5003 0 2.0 1e-06 
0.0 0.5004 0 2.0 1e-06 
0.0 0.5005 0 2.0 1e-06 
0.0 0.5006 0 2.0 1e-06 
0.0 0.5007 0 2.0 1e-06 
0.0 0.5008 0 2.0 1e-06 
0.0 0.5009 0 2.0 1e-06 
0.0 0.501 0 2.0 1e-06 
0.0 0.5011 0 2.0 1e-06 
0.0 0.5012 0 2.0 1e-06 
0.0 0.5013 0 2.0 1e-06 
0.0 0.5014 0 2.0 1e-06 
0.0 0.5015 0 2.0 1e-06 
0.0 0.5016 0 2.0 1e-06 
0.0 0.5017 0 2.0 1e-06 
0.0 0.5018 0 2.0 1e-06 
0.0 0.5019 0 2.0 1e-06 
0.0 0.502 0 2.0 1e-06 
0.0 0.5021 0 2.0 1e-06 
0.0 0.5022 0 2.0 1e-06 
0.0 0.5023 0 2.0 1e-06 
0.0 0.5024 0 2.0 1e-06 
0.0 0.5025 0 2.0 1e-06 
0.0 0.5026 0 2.0 1e-06 
0.0 0.5027 0 2.0 1e-06 
0.0 0.5028 0 2.0 1e-06 
0.0 0.5029 0 2.0 1e-06 
0.0 0.503 0 2.0 1e-06 
0.0 0.5031 0 2.0 1e-06 
0.0 0.5032 0 2.0 1e-06 
0.0 0.5033 0 2.0 1e-06 
0.0 0.5034 0 2.0 1e-06 
0.0 0.5035 0 2.0 1e-06 
0.0 0.5036 0 2.0 1e-06 
0.0 0.5037 0 2.0 1e-06 
0.0 0.5038 0 2.0 1e-06 
0.0 0.5039 0 2.0 1e-06 
0.0 0.504 0 2.0 1e-06 
0.0 0.5041 0 2.0 1e-06 
0.0 0.5042 0 2.0 1e-06 
0.0 0.5043 0 2.0 1e-06 
0.0 0.5044 0 2.0 1e-06 
0.0 0.5045 0 2.0 1e-06 
0.0 0.5046 0 2.0 1e-06 
0.0 0.5047 0 2.0 1e-06 
0.0 0.5048 0 2.0 1e-06 
0.0 0.5049 0 2.0 1e-06 
0.0 0.505 0 2.0 1e-06 
0.0 0.5051 0 2.0 1e-06 
0.0 0.5052 0 2.0 1e-06 
0.0 0.5053 0 2.0 1e-06 
0.0 0.5054 0 2.0 1e-06 
0.0 0.5055 0 2.0 1e-06 
0.0 0.5056 0 2.0 1e-06 
0.0 0.5057 0 2.0 1e-06 
0.0 0.5058 0 2.0 1e-06 
0.0 0.5059 0 2.0 1e-06 
0.0 0.506 0 2.0 1e-06 
0.0 0.5061 0 2.0 1e-06 
0.0 0.5062 0 2.0 1e-06 
0.0 0.5063 0 2.0 1e-06 
0.0 0.5064 0 2.0 1e-06 
0.0 0.5065 0 2.0 1e-06 
0.0 0.5066 0 2.0 1e-06 
0.0 0.5067 0 2.0 1e-06 
0.0 0.5068 0 2.0 1e-06 
0.0 0.5069 0 2.0 1e-06 
0.0 0.507 0 2.0 1e-06 
0.0 0.5071 0 2.0 1e-06 
0.0 0.5072 0 2.0 1e-06 
0.0 0.5073 0 2.0 1e-06 
0.0 0.5074 0 2.0 1e-06 
0.0 0.5075 0 2.0 1e-06 
0.0 0.5076 0 2.0 1e-06 
0.0 0.5077 0 2.0 1e-06 
0.0 0.5078 0 2.0 1e-06 
0.0 0.5079 0 2.0 1e-06 
0.0 0.508 0 2.0 1e-06 
0.0 0.5081 0 2.0 1e-06 
0.0 0.5082 0 2.0 1e-06 
0.0 0.5083 0 2.0 1e-06 
0.0 0.5084 0 2.0 1e-06 
0.0 0.5085 0 2.0 1e-06 
0.0 0.5086 0 2.0 1e-06 
0.0 0.5087 0 2.0 1e-06 
0.0 0.5088 0 2.0 1e-06 
0.0 0.5089 0 2.0 1e-06 
0.0 0.509 0 2.0 1e-06 
0.0 0.5091 0 2.0 1e-06 
0.0 0.5092 0 2.0 1e-06 
0.0 0.5093 0 2.0 1e-06 
0.0 0.5094 0 2.0 1e-06 
0.0 0.5095 0 2.0 1e-06 
0.0 0.5096 0 2.0 1e-06 
0.0 0.5097 0 2.0 1e-06 
0.0 0.5098 0 2.0 1e-06 
0.0 0.5099 0 2.0 1e-06 
0.0 0.51 0 2.0 1e-06 
0.0 0.5101 0 2.0 1e-06 
0.0 0.5102 0 2.0 1e-06 
0.0 0.5103 0 2.0 1e-06 
0.0 0.5104 0 2.0 1e-06 
0.0 0.5105 0 2.0 1e-06 
0.0 0.5106 0 2.0 1e-06 
0.0 0.5107 0 2.0 1e-06 
0.0 0.5108 0 2.0 1e-06 
0.0 0.5109 0 2.0 1e-06 
0.0 0.511 0 2.0 1e-06 
0.0 0.5111 0 2.0 1e-06 
0.0 0.5112 0 2.0 1e-06 
0.0 0.5113 0 2.0 1e-06 
0.0 0.5114 0 2.0 1e-06 
0.0 0.5115 0 2.0 1e-06 
0.0 0.5116 0 2.0 1e-06 
0.0 0.5117 0 2.0 1e-06 
0.0 0.5118 0 2.0 1e-06 
0.0 0.5119 0 2.0 1e-06 
0.0 0.512 0 2.0 1e-06 
0.0 0.5121 0 2.0 1e-06 
0.0 0.5122 0 2.0 1e-06 
0.0 0.5123 0 2.0 1e-06 
0.0 0.5124 0 2.0 1e-06 
0.0 0.5125 0 2.0 1e-06 
0.0 0.5126 0 2.0 1e-06 
0.0 0.5127 0 2.0 1e-06 
0.0 0.5128 0 2.0 1e-06 
0.0 0.5129 0 2.0 1e-06 
0.0 0.513 0 2.0 1e-06 
0.0 0.5131 0 2.0 1e-06 
0.0 0.5132 0 2.0 1e-06 
0.0 0.5133 0 2.0 1e-06 
0.0 0.5134 0 2.0 1e-06 
0.0 0.5135 0 2.0 1e-06 
0.0 0.5136 0 2.0 1e-06 
0.0 0.5137 0 2.0 1e-06 
0.0 0.5138 0 2.0 1e-06 
0.0 0.5139 0 2.0 1e-06 
0.0 0.514 0 2.0 1e-06 
0.0 0.5141 0 2.0 1e-06 
0.0 0.5142 0 2.0 1e-06 
0.0 0.5143 0 2.0 1e-06 
0.0 0.5144 0 2.0 1e-06 
0.0 0.5145 0 2.0 1e-06 
0.0 0.5146 0 2.0 1e-06 
0.0 0.5147 0 2.0 1e-06 
0.0 0.5148 0 2.0 1e-06 
0.0 0.5149 0 2.0 1e-06 
0.0 0.515 0 2.0 1e-06 
0.0 0.5151 0 2.0 1e-06 
0.0 0.5152 0 2.0 1e-06 
0.0 0.5153 0 2.0 1e-06 
0.0 0.5154 0 2.0 1e-06 
0.0 0.5155 0 2.0 1e-06 
0.0 0.5156 0 2.0 1e-06 
0.0 0.5157 0 2.0 1e-06 
0.0 0.5158 0 2.0 1e-06 
0.0 0.5159 0 2.0 1e-06 
0.0 0.516 0 2.0 1e-06 
0.0 0.5161 0 2.0 1e-06 
0.0 0.5162 0 2.0 1e-06 
0.0 0.5163 0 2.0 1e-06 
0.0 0.5164 0 2.0 1e-06 
0.0 0.5165 0 2.0 1e-06 
0.0 0.5166 0 2.0 1e-06 
0.0 0.5167 0 2.0 1e-06 
0.0 0.5168 0 2.0 1e-06 
0.0 0.5169 0 2.0 1e-06 
0.0 0.517 0 2.0 1e-06 
0.0 0.5171 0 2.0 1e-06 
0.0 0.5172 0 2.0 1e-06 
0.0 0.5173 0 2.0 1e-06 
0.0 0.5174 0 2.0 1e-06 
0.0 0.5175 0 2.0 1e-06 
0.0 0.5176 0 2.0 1e-06 
0.0 0.5177 0 2.0 1e-06 
0.0 0.5178 0 2.0 1e-06 
0.0 0.5179 0 2.0 1e-06 
0.0 0.518 0 2.0 1e-06 
0.0 0.5181 0 2.0 1e-06 
0.0 0.5182 0 2.0 1e-06 
0.0 0.5183 0 2.0 1e-06 
0.0 0.5184 0 2.0 1e-06 
0.0 0.5185 0 2.0 1e-06 
0.0 0.5186 0 2.0 1e-06 
0.0 0.5187 0 2.0 1e-06 
0.0 0.5188 0 2.0 1e-06 
0.0 0.5189 0 2.0 1e-06 
0.0 0.519 0 2.0 1e-06 
0.0 0.5191 0 2.0 1e-06 
0.0 0.5192 0 2.0 1e-06 
0.0 0.5193 0 2.0 1e-06 
0.0 0.5194 0 2.0 1e-06 
0.0 0.5195 0 2.0 1e-06 
0.0 0.5196 0 2.0 1e-06 
0.0 0.5197 0 2.0 1e-06 
0.0 0.5198 0 2.0 1e-06 
0.0 0.5199 0 2.0 1e-06 
0.0 0.52 0 2.0 1e-06 
0.0 0.5201 0 2.0 1e-06 
0.0 0.5202 0 2.0 1e-06 
0.0 0.5203 0 2.0 1e-06 
0.0 0.5204 0 2.0 1e-06 
0.0 0.5205 0 2.0 1e-06 
0.0 0.5206 0 2.0 1e-06 
0.0 0.5207 0 2.0 1e-06 
0.0 0.5208 0 2.0 1e-06 
0.0 0.5209 0 2.0 1e-06 
0.0 0.521 0 2.0 1e-06 
0.0 0.5211 0 2.0 1e-06 
0.0 0.5212 0 2.0 1e-06 
0.0 0.5213 0 2.0 1e-06 
0.0 0.5214 0 2.0 1e-06 
0.0 0.5215 0 2.0 1e-06 
0.0 0.5216 0 2.0 1e-06 
0.0 0.5217 0 2.0 1e-06 
0.0 0.5218 0 2.0 1e-06 
0.0 0.5219 0 2.0 1e-06 
0.0 0.522 0 2.0 1e-06 
0.0 0.5221 0 2.0 1e-06 
0.0 0.5222 0 2.0 1e-06 
0.0 0.5223 0 2.0 1e-06 
0.0 0.5224 0 2.0 1e-06 
0.0 0.5225 0 2.0 1e-06 
0.0 0.5226 0 2.0 1e-06 
0.0 0.5227 0 2.0 1e-06 
0.0 0.5228 0 2.0 1e-06 
0.0 0.5229 0 2.0 1e-06 
0.0 0.523 0 2.0 1e-06 
0.0 0.5231 0 2.0 1e-06 
0.0 0.5232 0 2.0 1e-06 
0.0 0.5233 0 2.0 1e-06 
0.0 0.5234 0 2.0 1e-06 
0.0 0.5235 0 2.0 1e-06 
0.0 0.5236 0 2.0 1e-06 
0.0 0.5237 0 2.0 1e-06 
0.0 0.5238 0 2.0 1e-06 
0.0 0.5239 0 2.0 1e-06 
0.0 0.524 0 2.0 1e-06 
0.0 0.5241 0 2.0 1e-06 
0.0 0.5242 0 2.0 1e-06 
0.0 0.5243 0 2.0 1e-06 
0.0 0.5244 0 2.0 1e-06 
0.0 0.5245 0 2.0 1e-06 
0.0 0.5246 0 2.0 1e-06 
0.0 0.5247 0 2.0 1e-06 
0.0 0.5248 0 2.0 1e-06 
0.0 0.5249 0 2.0 1e-06 
0.0 0.525 0 2.0 1e-06 
0.0 0.5251 0 2.0 1e-06 
0.0 0.5252 0 2.0 1e-06 
0.0 0.5253 0 2.0 1e-06 
0.0 0.5254 0 2.0 1e-06 
0.0 0.5255 0 2.0 1e-06 
0.0 0.5256 0 2.0 1e-06 
0.0 0.5257 0 2.0 1e-06 
0.0 0.5258 0 2.0 1e-06 
0.0 0.5259 0 2.0 1e-06 
0.0 0.526 0 2.0 1e-06 
0.0 0.5261 0 2.0 1e-06 
0.0 0.5262 0 2.0 1e-06 
0.0 0.5263 0 2.0 1e-06 
0.0 0.5264 0 2.0 1e-06 
0.0 0.5265 0 2.0 1e-06 
0.0 0.5266 0 2.0 1e-06 
0.0 0.5267 0 2.0 1e-06 
0.0 0.5268 0 2.0 1e-06 
0.0 0.5269 0 2.0 1e-06 
0.0 0.527 0 2.0 1e-06 
0.0 0.5271 0 2.0 1e-06 
0.0 0.5272 0 2.0 1e-06 
0.0 0.5273 0 2.0 1e-06 
0.0 0.5274 0 2.0 1e-06 
0.0 0.5275 0 2.0 1e-06 
0.0 0.5276 0 2.0 1e-06 
0.0 0.5277 0 2.0 1e-06 
0.0 0.5278 0 2.0 1e-06 
0.0 0.5279 0 2.0 1e-06 
0.0 0.528 0 2.0 1e-06 
0.0 0.5281 0 2.0 1e-06 
0.0 0.5282 0 2.0 1e-06 
0.0 0.5283 0 2.0 1e-06 
0.0 0.5284 0 2.0 1e-06 
0.0 0.5285 0 2.0 1e-06 
0.0 0.5286 0 2.0 1e-06 
0.0 0.5287 0 2.0 1e-06 
0.0 0.5288 0 2.0 1e-06 
0.0 0.5289 0 2.0 1e-06 
0.0 0.529 0 2.0 1e-06 
0.0 0.5291 0 2.0 1e-06 
0.0 0.5292 0 2.0 1e-06 
0.0 0.5293 0 2.0 1e-06 
0.0 0.5294 0 2.0 1e-06 
0.0 0.5295 0 2.0 1e-06 
0.0 0.5296 0 2.0 1e-06 
0.0 0.5297 0 2.0 1e-06 
0.0 0.5298 0 2.0 1e-06 
0.0 0.5299 0 2.0 1e-06 
0.0 0.53 0 2.0 1e-06 
0.0 0.5301 0 2.0 1e-06 
0.0 0.5302 0 2.0 1e-06 
0.0 0.5303 0 2.0 1e-06 
0.0 0.5304 0 2.0 1e-06 
0.0 0.5305 0 2.0 1e-06 
0.0 0.5306 0 2.0 1e-06 
0.0 0.5307 0 2.0 1e-06 
0.0 0.5308 0 2.0 1e-06 
0.0 0.5309 0 2.0 1e-06 
0.0 0.531 0 2.0 1e-06 
0.0 0.5311 0 2.0 1e-06 
0.0 0.5312 0 2.0 1e-06 
0.0 0.5313 0 2.0 1e-06 
0.0 0.5314 0 2.0 1e-06 
0.0 0.5315 0 2.0 1e-06 
0.0 0.5316 0 2.0 1e-06 
0.0 0.5317 0 2.0 1e-06 
0.0 0.5318 0 2.0 1e-06 
0.0 0.5319 0 2.0 1e-06 
0.0 0.532 0 2.0 1e-06 
0.0 0.5321 0 2.0 1e-06 
0.0 0.5322 0 2.0 1e-06 
0.0 0.5323 0 2.0 1e-06 
0.0 0.5324 0 2.0 1e-06 
0.0 0.5325 0 2.0 1e-06 
0.0 0.5326 0 2.0 1e-06 
0.0 0.5327 0 2.0 1e-06 
0.0 0.5328 0 2.0 1e-06 
0.0 0.5329 0 2.0 1e-06 
0.0 0.533 0 2.0 1e-06 
0.0 0.5331 0 2.0 1e-06 
0.0 0.5332 0 2.0 1e-06 
0.0 0.5333 0 2.0 1e-06 
0.0 0.5334 0 2.0 1e-06 
0.0 0.5335 0 2.0 1e-06 
0.0 0.5336 0 2.0 1e-06 
0.0 0.5337 0 2.0 1e-06 
0.0 0.5338 0 2.0 1e-06 
0.0 0.5339 0 2.0 1e-06 
0.0 0.534 0 2.0 1e-06 
0.0 0.5341 0 2.0 1e-06 
0.0 0.5342 0 2.0 1e-06 
0.0 0.5343 0 2.0 1e-06 
0.0 0.5344 0 2.0 1e-06 
0.0 0.5345 0 2.0 1e-06 
0.0 0.5346 0 2.0 1e-06 
0.0 0.5347 0 2.0 1e-06 
0.0 0.5348 0 2.0 1e-06 
0.0 0.5349 0 2.0 1e-06 
0.0 0.535 0 2.0 1e-06 
0.0 0.5351 0 2.0 1e-06 
0.0 0.5352 0 2.0 1e-06 
0.0 0.5353 0 2.0 1e-06 
0.0 0.5354 0 2.0 1e-06 
0.0 0.5355 0 2.0 1e-06 
0.0 0.5356 0 2.0 1e-06 
0.0 0.5357 0 2.0 1e-06 
0.0 0.5358 0 2.0 1e-06 
0.0 0.5359 0 2.0 1e-06 
0.0 0.536 0 2.0 1e-06 
0.0 0.5361 0 2.0 1e-06 
0.0 0.5362 0 2.0 1e-06 
0.0 0.5363 0 2.0 1e-06 
0.0 0.5364 0 2.0 1e-06 
0.0 0.5365 0 2.0 1e-06 
0.0 0.5366 0 2.0 1e-06 
0.0 0.5367 0 2.0 1e-06 
0.0 0.5368 0 2.0 1e-06 
0.0 0.5369 0 2.0 1e-06 
0.0 0.537 0 2.0 1e-06 
0.0 0.5371 0 2.0 1e-06 
0.0 0.5372 0 2.0 1e-06 
0.0 0.5373 0 2.0 1e-06 
0.0 0.5374 0 2.0 1e-06 
0.0 0.5375 0 2.0 1e-06 
0.0 0.5376 0 2.0 1e-06 
0.0 0.5377 0 2.0 1e-06 
0.0 0.5378 0 2.0 1e-06 
0.0 0.5379 0 2.0 1e-06 
0.0 0.538 0 2.0 1e-06 
0.0 0.5381 0 2.0 1e-06 
0.0 0.5382 0 2.0 1e-06 
0.0 0.5383 0 2.0 1e-06 
0.0 0.5384 0 2.0 1e-06 
0.0 0.5385 0 2.0 1e-06 
0.0 0.5386 0 2.0 1e-06 
0.0 0.5387 0 2.0 1e-06 
0.0 0.5388 0 2.0 1e-06 
0.0 0.5389 0 2.0 1e-06 
0.0 0.539 0 2.0 1e-06 
0.0 0.5391 0 2.0 1e-06 
0.0 0.5392 0 2.0 1e-06 
0.0 0.5393 0 2.0 1e-06 
0.0 0.5394 0 2.0 1e-06 
0.0 0.5395 0 2.0 1e-06 
0.0 0.5396 0 2.0 1e-06 
0.0 0.5397 0 2.0 1e-06 
0.0 0.5398 0 2.0 1e-06 
0.0 0.5399 0 2.0 1e-06 
0.0 0.54 0 2.0 1e-06 
0.0 0.5401 0 2.0 1e-06 
0.0 0.5402 0 2.0 1e-06 
0.0 0.5403 0 2.0 1e-06 
0.0 0.5404 0 2.0 1e-06 
0.0 0.5405 0 2.0 1e-06 
0.0 0.5406 0 2.0 1e-06 
0.0 0.5407 0 2.0 1e-06 
0.0 0.5408 0 2.0 1e-06 
0.0 0.5409 0 2.0 1e-06 
0.0 0.541 0 2.0 1e-06 
0.0 0.5411 0 2.0 1e-06 
0.0 0.5412 0 2.0 1e-06 
0.0 0.5413 0 2.0 1e-06 
0.0 0.5414 0 2.0 1e-06 
0.0 0.5415 0 2.0 1e-06 
0.0 0.5416 0 2.0 1e-06 
0.0 0.5417 0 2.0 1e-06 
0.0 0.5418 0 2.0 1e-06 
0.0 0.5419 0 2.0 1e-06 
0.0 0.542 0 2.0 1e-06 
0.0 0.5421 0 2.0 1e-06 
0.0 0.5422 0 2.0 1e-06 
0.0 0.5423 0 2.0 1e-06 
0.0 0.5424 0 2.0 1e-06 
0.0 0.5425 0 2.0 1e-06 
0.0 0.5426 0 2.0 1e-06 
0.0 0.5427 0 2.0 1e-06 
0.0 0.5428 0 2.0 1e-06 
0.0 0.5429 0 2.0 1e-06 
0.0 0.543 0 2.0 1e-06 
0.0 0.5431 0 2.0 1e-06 
0.0 0.5432 0 2.0 1e-06 
0.0 0.5433 0 2.0 1e-06 
0.0 0.5434 0 2.0 1e-06 
0.0 0.5435 0 2.0 1e-06 
0.0 0.5436 0 2.0 1e-06 
0.0 0.5437 0 2.0 1e-06 
0.0 0.5438 0 2.0 1e-06 
0.0 0.5439 0 2.0 1e-06 
0.0 0.544 0 2.0 1e-06 
0.0 0.5441 0 2.0 1e-06 
0.0 0.5442 0 2.0 1e-06 
0.0 0.5443 0 2.0 1e-06 
0.0 0.5444 0 2.0 1e-06 
0.0 0.5445 0 2.0 1e-06 
0.0 0.5446 0 2.0 1e-06 
0.0 0.5447 0 2.0 1e-06 
0.0 0.5448 0 2.0 1e-06 
0.0 0.5449 0 2.0 1e-06 
0.0 0.545 0 2.0 1e-06 
0.0 0.5451 0 2.0 1e-06 
0.0 0.5452 0 2.0 1e-06 
0.0 0.5453 0 2.0 1e-06 
0.0 0.5454 0 2.0 1e-06 
0.0 0.5455 0 2.0 1e-06 
0.0 0.5456 0 2.0 1e-06 
0.0 0.5457 0 2.0 1e-06 
0.0 0.5458 0 2.0 1e-06 
0.0 0.5459 0 2.0 1e-06 
0.0 0.546 0 2.0 1e-06 
0.0 0.5461 0 2.0 1e-06 
0.0 0.5462 0 2.0 1e-06 
0.0 0.5463 0 2.0 1e-06 
0.0 0.5464 0 2.0 1e-06 
0.0 0.5465 0 2.0 1e-06 
0.0 0.5466 0 2.0 1e-06 
0.0 0.5467 0 2.0 1e-06 
0.0 0.5468 0 2.0 1e-06 
0.0 0.5469 0 2.0 1e-06 
0.0 0.547 0 2.0 1e-06 
0.0 0.5471 0 2.0 1e-06 
0.0 0.5472 0 2.0 1e-06 
0.0 0.5473 0 2.0 1e-06 
0.0 0.5474 0 2.0 1e-06 
0.0 0.5475 0 2.0 1e-06 
0.0 0.5476 0 2.0 1e-06 
0.0 0.5477 0 2.0 1e-06 
0.0 0.5478 0 2.0 1e-06 
0.0 0.5479 0 2.0 1e-06 
0.0 0.548 0 2.0 1e-06 
0.0 0.5481 0 2.0 1e-06 
0.0 0.5482 0 2.0 1e-06 
0.0 0.5483 0 2.0 1e-06 
0.0 0.5484 0 2.0 1e-06 
0.0 0.5485 0 2.0 1e-06 
0.0 0.5486 0 2.0 1e-06 
0.0 0.5487 0 2.0 1e-06 
0.0 0.5488 0 2.0 1e-06 
0.0 0.5489 0 2.0 1e-06 
0.0 0.549 0 2.0 1e-06 
0.0 0.5491 0 2.0 1e-06 
0.0 0.5492 0 2.0 1e-06 
0.0 0.5493 0 2.0 1e-06 
0.0 0.5494 0 2.0 1e-06 
0.0 0.5495 0 2.0 1e-06 
0.0 0.5496 0 2.0 1e-06 
0.0 0.5497 0 2.0 1e-06 
0.0 0.5498 0 2.0 1e-06 
0.0 0.5499 0 2.0 1e-06 
0.0 0.55 0 2.0 1e-06 
0.0 0.5501 0 2.0 1e-06 
0.0 0.5502 0 2.0 1e-06 
0.0 0.5503 0 2.0 1e-06 
0.0 0.5504 0 2.0 1e-06 
0.0 0.5505 0 2.0 1e-06 
0.0 0.5506 0 2.0 1e-06 
0.0 0.5507 0 2.0 1e-06 
0.0 0.5508 0 2.0 1e-06 
0.0 0.5509 0 2.0 1e-06 
0.0 0.551 0 2.0 1e-06 
0.0 0.5511 0 2.0 1e-06 
0.0 0.5512 0 2.0 1e-06 
0.0 0.5513 0 2.0 1e-06 
0.0 0.5514 0 2.0 1e-06 
0.0 0.5515 0 2.0 1e-06 
0.0 0.5516 0 2.0 1e-06 
0.0 0.5517 0 2.0 1e-06 
0.0 0.5518 0 2.0 1e-06 
0.0 0.5519 0 2.0 1e-06 
0.0 0.552 0 2.0 1e-06 
0.0 0.5521 0 2.0 1e-06 
0.0 0.5522 0 2.0 1e-06 
0.0 0.5523 0 2.0 1e-06 
0.0 0.5524 0 2.0 1e-06 
0.0 0.5525 0 2.0 1e-06 
0.0 0.5526 0 2.0 1e-06 
0.0 0.5527 0 2.0 1e-06 
0.0 0.5528 0 2.0 1e-06 
0.0 0.5529 0 2.0 1e-06 
0.0 0.553 0 2.0 1e-06 
0.0 0.5531 0 2.0 1e-06 
0.0 0.5532 0 2.0 1e-06 
0.0 0.5533 0 2.0 1e-06 
0.0 0.5534 0 2.0 1e-06 
0.0 0.5535 0 2.0 1e-06 
0.0 0.5536 0 2.0 1e-06 
0.0 0.5537 0 2.0 1e-06 
0.0 0.5538 0 2.0 1e-06 
0.0 0.5539 0 2.0 1e-06 
0.0 0.554 0 2.0 1e-06 
0.0 0.5541 0 2.0 1e-06 
0.0 0.5542 0 2.0 1e-06 
0.0 0.5543 0 2.0 1e-06 
0.0 0.5544 0 2.0 1e-06 
0.0 0.5545 0 2.0 1e-06 
0.0 0.5546 0 2.0 1e-06 
0.0 0.5547 0 2.0 1e-06 
0.0 0.5548 0 2.0 1e-06 
0.0 0.5549 0 2.0 1e-06 
0.0 0.555 0 2.0 1e-06 
0.0 0.5551 0 2.0 1e-06 
0.0 0.5552 0 2.0 1e-06 
0.0 0.5553 0 2.0 1e-06 
0.0 0.5554 0 2.0 1e-06 
0.0 0.5555 0 2.0 1e-06 
0.0 0.5556 0 2.0 1e-06 
0.0 0.5557 0 2.0 1e-06 
0.0 0.5558 0 2.0 1e-06 
0.0 0.5559 0 2.0 1e-06 
0.0 0.556 0 2.0 1e-06 
0.0 0.5561 0 2.0 1e-06 
0.0 0.5562 0 2.0 1e-06 
0.0 0.5563 0 2.0 1e-06 
0.0 0.5564 0 2.0 1e-06 
0.0 0.5565 0 2.0 1e-06 
0.0 0.5566 0 2.0 1e-06 
0.0 0.5567 0 2.0 1e-06 
0.0 0.5568 0 2.0 1e-06 
0.0 0.5569 0 2.0 1e-06 
0.0 0.557 0 2.0 1e-06 
0.0 0.5571 0 2.0 1e-06 
0.0 0.5572 0 2.0 1e-06 
0.0 0.5573 0 2.0 1e-06 
0.0 0.5574 0 2.0 1e-06 
0.0 0.5575 0 2.0 1e-06 
0.0 0.5576 0 2.0 1e-06 
0.0 0.5577 0 2.0 1e-06 
0.0 0.5578 0 2.0 1e-06 
0.0 0.5579 0 2.0 1e-06 
0.0 0.558 0 2.0 1e-06 
0.0 0.5581 0 2.0 1e-06 
0.0 0.5582 0 2.0 1e-06 
0.0 0.5583 0 2.0 1e-06 
0.0 0.5584 0 2.0 1e-06 
0.0 0.5585 0 2.0 1e-06 
0.0 0.5586 0 2.0 1e-06 
0.0 0.5587 0 2.0 1e-06 
0.0 0.5588 0 2.0 1e-06 
0.0 0.5589 0 2.0 1e-06 
0.0 0.559 0 2.0 1e-06 
0.0 0.5591 0 2.0 1e-06 
0.0 0.5592 0 2.0 1e-06 
0.0 0.5593 0 2.0 1e-06 
0.0 0.5594 0 2.0 1e-06 
0.0 0.5595 0 2.0 1e-06 
0.0 0.5596 0 2.0 1e-06 
0.0 0.5597 0 2.0 1e-06 
0.0 0.5598 0 2.0 1e-06 
0.0 0.5599 0 2.0 1e-06 
0.0 0.56 0 2.0 1e-06 
0.0 0.5601 0 2.0 1e-06 
0.0 0.5602 0 2.0 1e-06 
0.0 0.5603 0 2.0 1e-06 
0.0 0.5604 0 2.0 1e-06 
0.0 0.5605 0 2.0 1e-06 
0.0 0.5606 0 2.0 1e-06 
0.0 0.5607 0 2.0 1e-06 
0.0 0.5608 0 2.0 1e-06 
0.0 0.5609 0 2.0 1e-06 
0.0 0.561 0 2.0 1e-06 
0.0 0.5611 0 2.0 1e-06 
0.0 0.5612 0 2.0 1e-06 
0.0 0.5613 0 2.0 1e-06 
0.0 0.5614 0 2.0 1e-06 
0.0 0.5615 0 2.0 1e-06 
0.0 0.5616 0 2.0 1e-06 
0.0 0.5617 0 2.0 1e-06 
0.0 0.5618 0 2.0 1e-06 
0.0 0.5619 0 2.0 1e-06 
0.0 0.562 0 2.0 1e-06 
0.0 0.5621 0 2.0 1e-06 
0.0 0.5622 0 2.0 1e-06 
0.0 0.5623 0 2.0 1e-06 
0.0 0.5624 0 2.0 1e-06 
0.0 0.5625 0 2.0 1e-06 
0.0 0.5626 0 2.0 1e-06 
0.0 0.5627 0 2.0 1e-06 
0.0 0.5628 0 2.0 1e-06 
0.0 0.5629 0 2.0 1e-06 
0.0 0.563 0 2.0 1e-06 
0.0 0.5631 0 2.0 1e-06 
0.0 0.5632 0 2.0 1e-06 
0.0 0.5633 0 2.0 1e-06 
0.0 0.5634 0 2.0 1e-06 
0.0 0.5635 0 2.0 1e-06 
0.0 0.5636 0 2.0 1e-06 
0.0 0.5637 0 2.0 1e-06 
0.0 0.5638 0 2.0 1e-06 
0.0 0.5639 0 2.0 1e-06 
0.0 0.564 0 2.0 1e-06 
0.0 0.5641 0 2.0 1e-06 
0.0 0.5642 0 2.0 1e-06 
0.0 0.5643 0 2.0 1e-06 
0.0 0.5644 0 2.0 1e-06 
0.0 0.5645 0 2.0 1e-06 
0.0 0.5646 0 2.0 1e-06 
0.0 0.5647 0 2.0 1e-06 
0.0 0.5648 0 2.0 1e-06 
0.0 0.5649 0 2.0 1e-06 
0.0 0.565 0 2.0 1e-06 
0.0 0.5651 0 2.0 1e-06 
0.0 0.5652 0 2.0 1e-06 
0.0 0.5653 0 2.0 1e-06 
0.0 0.5654 0 2.0 1e-06 
0.0 0.5655 0 2.0 1e-06 
0.0 0.5656 0 2.0 1e-06 
0.0 0.5657 0 2.0 1e-06 
0.0 0.5658 0 2.0 1e-06 
0.0 0.5659 0 2.0 1e-06 
0.0 0.566 0 2.0 1e-06 
0.0 0.5661 0 2.0 1e-06 
0.0 0.5662 0 2.0 1e-06 
0.0 0.5663 0 2.0 1e-06 
0.0 0.5664 0 2.0 1e-06 
0.0 0.5665 0 2.0 1e-06 
0.0 0.5666 0 2.0 1e-06 
0.0 0.5667 0 2.0 1e-06 
0.0 0.5668 0 2.0 1e-06 
0.0 0.5669 0 2.0 1e-06 
0.0 0.567 0 2.0 1e-06 
0.0 0.5671 0 2.0 1e-06 
0.0 0.5672 0 2.0 1e-06 
0.0 0.5673 0 2.0 1e-06 
0.0 0.5674 0 2.0 1e-06 
0.0 0.5675 0 2.0 1e-06 
0.0 0.5676 0 2.0 1e-06 
0.0 0.5677 0 2.0 1e-06 
0.0 0.5678 0 2.0 1e-06 
0.0 0.5679 0 2.0 1e-06 
0.0 0.568 0 2.0 1e-06 
0.0 0.5681 0 2.0 1e-06 
0.0 0.5682 0 2.0 1e-06 
0.0 0.5683 0 2.0 1e-06 
0.0 0.5684 0 2.0 1e-06 
0.0 0.5685 0 2.0 1e-06 
0.0 0.5686 0 2.0 1e-06 
0.0 0.5687 0 2.0 1e-06 
0.0 0.5688 0 2.0 1e-06 
0.0 0.5689 0 2.0 1e-06 
0.0 0.569 0 2.0 1e-06 
0.0 0.5691 0 2.0 1e-06 
0.0 0.5692 0 2.0 1e-06 
0.0 0.5693 0 2.0 1e-06 
0.0 0.5694 0 2.0 1e-06 
0.0 0.5695 0 2.0 1e-06 
0.0 0.5696 0 2.0 1e-06 
0.0 0.5697 0 2.0 1e-06 
0.0 0.5698 0 2.0 1e-06 
0.0 0.5699 0 2.0 1e-06 
0.0 0.57 0 2.0 1e-06 
0.0 0.5701 0 2.0 1e-06 
0.0 0.5702 0 2.0 1e-06 
0.0 0.5703 0 2.0 1e-06 
0.0 0.5704 0 2.0 1e-06 
0.0 0.5705 0 2.0 1e-06 
0.0 0.5706 0 2.0 1e-06 
0.0 0.5707 0 2.0 1e-06 
0.0 0.5708 0 2.0 1e-06 
0.0 0.5709 0 2.0 1e-06 
0.0 0.571 0 2.0 1e-06 
0.0 0.5711 0 2.0 1e-06 
0.0 0.5712 0 2.0 1e-06 
0.0 0.5713 0 2.0 1e-06 
0.0 0.5714 0 2.0 1e-06 
0.0 0.5715 0 2.0 1e-06 
0.0 0.5716 0 2.0 1e-06 
0.0 0.5717 0 2.0 1e-06 
0.0 0.5718 0 2.0 1e-06 
0.0 0.5719 0 2.0 1e-06 
0.0 0.572 0 2.0 1e-06 
0.0 0.5721 0 2.0 1e-06 
0.0 0.5722 0 2.0 1e-06 
0.0 0.5723 0 2.0 1e-06 
0.0 0.5724 0 2.0 1e-06 
0.0 0.5725 0 2.0 1e-06 
0.0 0.5726 0 2.0 1e-06 
0.0 0.5727 0 2.0 1e-06 
0.0 0.5728 0 2.0 1e-06 
0.0 0.5729 0 2.0 1e-06 
0.0 0.573 0 2.0 1e-06 
0.0 0.5731 0 2.0 1e-06 
0.0 0.5732 0 2.0 1e-06 
0.0 0.5733 0 2.0 1e-06 
0.0 0.5734 0 2.0 1e-06 
0.0 0.5735 0 2.0 1e-06 
0.0 0.5736 0 2.0 1e-06 
0.0 0.5737 0 2.0 1e-06 
0.0 0.5738 0 2.0 1e-06 
0.0 0.5739 0 2.0 1e-06 
0.0 0.574 0 2.0 1e-06 
0.0 0.5741 0 2.0 1e-06 
0.0 0.5742 0 2.0 1e-06 
0.0 0.5743 0 2.0 1e-06 
0.0 0.5744 0 2.0 1e-06 
0.0 0.5745 0 2.0 1e-06 
0.0 0.5746 0 2.0 1e-06 
0.0 0.5747 0 2.0 1e-06 
0.0 0.5748 0 2.0 1e-06 
0.0 0.5749 0 2.0 1e-06 
0.0 0.575 0 2.0 1e-06 
0.0 0.5751 0 2.0 1e-06 
0.0 0.5752 0 2.0 1e-06 
0.0 0.5753 0 2.0 1e-06 
0.0 0.5754 0 2.0 1e-06 
0.0 0.5755 0 2.0 1e-06 
0.0 0.5756 0 2.0 1e-06 
0.0 0.5757 0 2.0 1e-06 
0.0 0.5758 0 2.0 1e-06 
0.0 0.5759 0 2.0 1e-06 
0.0 0.576 0 2.0 1e-06 
0.0 0.5761 0 2.0 1e-06 
0.0 0.5762 0 2.0 1e-06 
0.0 0.5763 0 2.0 1e-06 
0.0 0.5764 0 2.0 1e-06 
0.0 0.5765 0 2.0 1e-06 
0.0 0.5766 0 2.0 1e-06 
0.0 0.5767 0 2.0 1e-06 
0.0 0.5768 0 2.0 1e-06 
0.0 0.5769 0 2.0 1e-06 
0.0 0.577 0 2.0 1e-06 
0.0 0.5771 0 2.0 1e-06 
0.0 0.5772 0 2.0 1e-06 
0.0 0.5773 0 2.0 1e-06 
0.0 0.5774 0 2.0 1e-06 
0.0 0.5775 0 2.0 1e-06 
0.0 0.5776 0 2.0 1e-06 
0.0 0.5777 0 2.0 1e-06 
0.0 0.5778 0 2.0 1e-06 
0.0 0.5779 0 2.0 1e-06 
0.0 0.578 0 2.0 1e-06 
0.0 0.5781 0 2.0 1e-06 
0.0 0.5782 0 2.0 1e-06 
0.0 0.5783 0 2.0 1e-06 
0.0 0.5784 0 2.0 1e-06 
0.0 0.5785 0 2.0 1e-06 
0.0 0.5786 0 2.0 1e-06 
0.0 0.5787 0 2.0 1e-06 
0.0 0.5788 0 2.0 1e-06 
0.0 0.5789 0 2.0 1e-06 
0.0 0.579 0 2.0 1e-06 
0.0 0.5791 0 2.0 1e-06 
0.0 0.5792 0 2.0 1e-06 
0.0 0.5793 0 2.0 1e-06 
0.0 0.5794 0 2.0 1e-06 
0.0 0.5795 0 2.0 1e-06 
0.0 0.5796 0 2.0 1e-06 
0.0 0.5797 0 2.0 1e-06 
0.0 0.5798 0 2.0 1e-06 
0.0 0.5799 0 2.0 1e-06 
0.0 0.58 0 2.0 1e-06 
0.0 0.5801 0 2.0 1e-06 
0.0 0.5802 0 2.0 1e-06 
0.0 0.5803 0 2.0 1e-06 
0.0 0.5804 0 2.0 1e-06 
0.0 0.5805 0 2.0 1e-06 
0.0 0.5806 0 2.0 1e-06 
0.0 0.5807 0 2.0 1e-06 
0.0 0.5808 0 2.0 1e-06 
0.0 0.5809 0 2.0 1e-06 
0.0 0.581 0 2.0 1e-06 
0.0 0.5811 0 2.0 1e-06 
0.0 0.5812 0 2.0 1e-06 
0.0 0.5813 0 2.0 1e-06 
0.0 0.5814 0 2.0 1e-06 
0.0 0.5815 0 2.0 1e-06 
0.0 0.5816 0 2.0 1e-06 
0.0 0.5817 0 2.0 1e-06 
0.0 0.5818 0 2.0 1e-06 
0.0 0.5819 0 2.0 1e-06 
0.0 0.582 0 2.0 1e-06 
0.0 0.5821 0 2.0 1e-06 
0.0 0.5822 0 2.0 1e-06 
0.0 0.5823 0 2.0 1e-06 
0.0 0.5824 0 2.0 1e-06 
0.0 0.5825 0 2.0 1e-06 
0.0 0.5826 0 2.0 1e-06 
0.0 0.5827 0 2.0 1e-06 
0.0 0.5828 0 2.0 1e-06 
0.0 0.5829 0 2.0 1e-06 
0.0 0.583 0 2.0 1e-06 
0.0 0.5831 0 2.0 1e-06 
0.0 0.5832 0 2.0 1e-06 
0.0 0.5833 0 2.0 1e-06 
0.0 0.5834 0 2.0 1e-06 
0.0 0.5835 0 2.0 1e-06 
0.0 0.5836 0 2.0 1e-06 
0.0 0.5837 0 2.0 1e-06 
0.0 0.5838 0 2.0 1e-06 
0.0 0.5839 0 2.0 1e-06 
0.0 0.584 0 2.0 1e-06 
0.0 0.5841 0 2.0 1e-06 
0.0 0.5842 0 2.0 1e-06 
0.0 0.5843 0 2.0 1e-06 
0.0 0.5844 0 2.0 1e-06 
0.0 0.5845 0 2.0 1e-06 
0.0 0.5846 0 2.0 1e-06 
0.0 0.5847 0 2.0 1e-06 
0.0 0.5848 0 2.0 1e-06 
0.0 0.5849 0 2.0 1e-06 
0.0 0.585 0 2.0 1e-06 
0.0 0.5851 0 2.0 1e-06 
0.0 0.5852 0 2.0 1e-06 
0.0 0.5853 0 2.0 1e-06 
0.0 0.5854 0 2.0 1e-06 
0.0 0.5855 0 2.0 1e-06 
0.0 0.5856 0 2.0 1e-06 
0.0 0.5857 0 2.0 1e-06 
0.0 0.5858 0 2.0 1e-06 
0.0 0.5859 0 2.0 1e-06 
0.0 0.586 0 2.0 1e-06 
0.0 0.5861 0 2.0 1e-06 
0.0 0.5862 0 2.0 1e-06 
0.0 0.5863 0 2.0 1e-06 
0.0 0.5864 0 2.0 1e-06 
0.0 0.5865 0 2.0 1e-06 
0.0 0.5866 0 2.0 1e-06 
0.0 0.5867 0 2.0 1e-06 
0.0 0.5868 0 2.0 1e-06 
0.0 0.5869 0 2.0 1e-06 
0.0 0.587 0 2.0 1e-06 
0.0 0.5871 0 2.0 1e-06 
0.0 0.5872 0 2.0 1e-06 
0.0 0.5873 0 2.0 1e-06 
0.0 0.5874 0 2.0 1e-06 
0.0 0.5875 0 2.0 1e-06 
0.0 0.5876 0 2.0 1e-06 
0.0 0.5877 0 2.0 1e-06 
0.0 0.5878 0 2.0 1e-06 
0.0 0.5879 0 2.0 1e-06 
0.0 0.588 0 2.0 1e-06 
0.0 0.5881 0 2.0 1e-06 
0.0 0.5882 0 2.0 1e-06 
0.0 0.5883 0 2.0 1e-06 
0.0 0.5884 0 2.0 1e-06 
0.0 0.5885 0 2.0 1e-06 
0.0 0.5886 0 2.0 1e-06 
0.0 0.5887 0 2.0 1e-06 
0.0 0.5888 0 2.0 1e-06 
0.0 0.5889 0 2.0 1e-06 
0.0 0.589 0 2.0 1e-06 
0.0 0.5891 0 2.0 1e-06 
0.0 0.5892 0 2.0 1e-06 
0.0 0.5893 0 2.0 1e-06 
0.0 0.5894 0 2.0 1e-06 
0.0 0.5895 0 2.0 1e-06 
0.0 0.5896 0 2.0 1e-06 
0.0 0.5897 0 2.0 1e-06 
0.0 0.5898 0 2.0 1e-06 
0.0 0.5899 0 2.0 1e-06 
0.0 0.59 0 2.0 1e-06 
0.0 0.5901 0 2.0 1e-06 
0.0 0.5902 0 2.0 1e-06 
0.0 0.5903 0 2.0 1e-06 
0.0 0.5904 0 2.0 1e-06 
0.0 0.5905 0 2.0 1e-06 
0.0 0.5906 0 2.0 1e-06 
0.0 0.5907 0 2.0 1e-06 
0.0 0.5908 0 2.0 1e-06 
0.0 0.5909 0 2.0 1e-06 
0.0 0.591 0 2.0 1e-06 
0.0 0.5911 0 2.0 1e-06 
0.0 0.5912 0 2.0 1e-06 
0.0 0.5913 0 2.0 1e-06 
0.0 0.5914 0 2.0 1e-06 
0.0 0.5915 0 2.0 1e-06 
0.0 0.5916 0 2.0 1e-06 
0.0 0.5917 0 2.0 1e-06 
0.0 0.5918 0 2.0 1e-06 
0.0 0.5919 0 2.0 1e-06 
0.0 0.592 0 2.0 1e-06 
0.0 0.5921 0 2.0 1e-06 
0.0 0.5922 0 2.0 1e-06 
0.0 0.5923 0 2.0 1e-06 
0.0 0.5924 0 2.0 1e-06 
0.0 0.5925 0 2.0 1e-06 
0.0 0.5926 0 2.0 1e-06 
0.0 0.5927 0 2.0 1e-06 
0.0 0.5928 0 2.0 1e-06 
0.0 0.5929 0 2.0 1e-06 
0.0 0.593 0 2.0 1e-06 
0.0 0.5931 0 2.0 1e-06 
0.0 0.5932 0 2.0 1e-06 
0.0 0.5933 0 2.0 1e-06 
0.0 0.5934 0 2.0 1e-06 
0.0 0.5935 0 2.0 1e-06 
0.0 0.5936 0 2.0 1e-06 
0.0 0.5937 0 2.0 1e-06 
0.0 0.5938 0 2.0 1e-06 
0.0 0.5939 0 2.0 1e-06 
0.0 0.594 0 2.0 1e-06 
0.0 0.5941 0 2.0 1e-06 
0.0 0.5942 0 2.0 1e-06 
0.0 0.5943 0 2.0 1e-06 
0.0 0.5944 0 2.0 1e-06 
0.0 0.5945 0 2.0 1e-06 
0.0 0.5946 0 2.0 1e-06 
0.0 0.5947 0 2.0 1e-06 
0.0 0.5948 0 2.0 1e-06 
0.0 0.5949 0 2.0 1e-06 
0.0 0.595 0 2.0 1e-06 
0.0 0.5951 0 2.0 1e-06 
0.0 0.5952 0 2.0 1e-06 
0.0 0.5953 0 2.0 1e-06 
0.0 0.5954 0 2.0 1e-06 
0.0 0.5955 0 2.0 1e-06 
0.0 0.5956 0 2.0 1e-06 
0.0 0.5957 0 2.0 1e-06 
0.0 0.5958 0 2.0 1e-06 
0.0 0.5959 0 2.0 1e-06 
0.0 0.596 0 2.0 1e-06 
0.0 0.5961 0 2.0 1e-06 
0.0 0.5962 0 2.0 1e-06 
0.0 0.5963 0 2.0 1e-06 
0.0 0.5964 0 2.0 1e-06 
0.0 0.5965 0 2.0 1e-06 
0.0 0.5966 0 2.0 1e-06 
0.0 0.5967 0 2.0 1e-06 
0.0 0.5968 0 2.0 1e-06 
0.0 0.5969 0 2.0 1e-06 
0.0 0.597 0 2.0 1e-06 
0.0 0.5971 0 2.0 1e-06 
0.0 0.5972 0 2.0 1e-06 
0.0 0.5973 0 2.0 1e-06 
0.0 0.5974 0 2.0 1e-06 
0.0 0.5975 0 2.0 1e-06 
0.0 0.5976 0 2.0 1e-06 
0.0 0.5977 0 2.0 1e-06 
0.0 0.5978 0 2.0 1e-06 
0.0 0.5979 0 2.0 1e-06 
0.0 0.598 0 2.0 1e-06 
0.0 0.5981 0 2.0 1e-06 
0.0 0.5982 0 2.0 1e-06 
0.0 0.5983 0 2.0 1e-06 
0.0 0.5984 0 2.0 1e-06 
0.0 0.5985 0 2.0 1e-06 
0.0 0.5986 0 2.0 1e-06 
0.0 0.5987 0 2.0 1e-06 
0.0 0.5988 0 2.0 1e-06 
0.0 0.5989 0 2.0 1e-06 
0.0 0.599 0 2.0 1e-06 
0.0 0.5991 0 2.0 1e-06 
0.0 0.5992 0 2.0 1e-06 
0.0 0.5993 0 2.0 1e-06 
0.0 0.5994 0 2.0 1e-06 
0.0 0.5995 0 2.0 1e-06 
0.0 0.5996 0 2.0 1e-06 
0.0 0.5997 0 2.0 1e-06 
0.0 0.5998 0 2.0 1e-06 
0.0 0.5999 0 2.0 1e-06 
0.0 0.6 0 2.0 1e-06 
0.0 0.6001 0 2.0 1e-06 
0.0 0.6002 0 2.0 1e-06 
0.0 0.6003 0 2.0 1e-06 
0.0 0.6004 0 2.0 1e-06 
0.0 0.6005 0 2.0 1e-06 
0.0 0.6006 0 2.0 1e-06 
0.0 0.6007 0 2.0 1e-06 
0.0 0.6008 0 2.0 1e-06 
0.0 0.6009 0 2.0 1e-06 
0.0 0.601 0 2.0 1e-06 
0.0 0.6011 0 2.0 1e-06 
0.0 0.6012 0 2.0 1e-06 
0.0 0.6013 0 2.0 1e-06 
0.0 0.6014 0 2.0 1e-06 
0.0 0.6015 0 2.0 1e-06 
0.0 0.6016 0 2.0 1e-06 
0.0 0.6017 0 2.0 1e-06 
0.0 0.6018 0 2.0 1e-06 
0.0 0.6019 0 2.0 1e-06 
0.0 0.602 0 2.0 1e-06 
0.0 0.6021 0 2.0 1e-06 
0.0 0.6022 0 2.0 1e-06 
0.0 0.6023 0 2.0 1e-06 
0.0 0.6024 0 2.0 1e-06 
0.0 0.6025 0 2.0 1e-06 
0.0 0.6026 0 2.0 1e-06 
0.0 0.6027 0 2.0 1e-06 
0.0 0.6028 0 2.0 1e-06 
0.0 0.6029 0 2.0 1e-06 
0.0 0.603 0 2.0 1e-06 
0.0 0.6031 0 2.0 1e-06 
0.0 0.6032 0 2.0 1e-06 
0.0 0.6033 0 2.0 1e-06 
0.0 0.6034 0 2.0 1e-06 
0.0 0.6035 0 2.0 1e-06 
0.0 0.6036 0 2.0 1e-06 
0.0 0.6037 0 2.0 1e-06 
0.0 0.6038 0 2.0 1e-06 
0.0 0.6039 0 2.0 1e-06 
0.0 0.604 0 2.0 1e-06 
0.0 0.6041 0 2.0 1e-06 
0.0 0.6042 0 2.0 1e-06 
0.0 0.6043 0 2.0 1e-06 
0.0 0.6044 0 2.0 1e-06 
0.0 0.6045 0 2.0 1e-06 
0.0 0.6046 0 2.0 1e-06 
0.0 0.6047 0 2.0 1e-06 
0.0 0.6048 0 2.0 1e-06 
0.0 0.6049 0 2.0 1e-06 
0.0 0.605 0 2.0 1e-06 
0.0 0.6051 0 2.0 1e-06 
0.0 0.6052 0 2.0 1e-06 
0.0 0.6053 0 2.0 1e-06 
0.0 0.6054 0 2.0 1e-06 
0.0 0.6055 0 2.0 1e-06 
0.0 0.6056 0 2.0 1e-06 
0.0 0.6057 0 2.0 1e-06 
0.0 0.6058 0 2.0 1e-06 
0.0 0.6059 0 2.0 1e-06 
0.0 0.606 0 2.0 1e-06 
0.0 0.6061 0 2.0 1e-06 
0.0 0.6062 0 2.0 1e-06 
0.0 0.6063 0 2.0 1e-06 
0.0 0.6064 0 2.0 1e-06 
0.0 0.6065 0 2.0 1e-06 
0.0 0.6066 0 2.0 1e-06 
0.0 0.6067 0 2.0 1e-06 
0.0 0.6068 0 2.0 1e-06 
0.0 0.6069 0 2.0 1e-06 
0.0 0.607 0 2.0 1e-06 
0.0 0.6071 0 2.0 1e-06 
0.0 0.6072 0 2.0 1e-06 
0.0 0.6073 0 2.0 1e-06 
0.0 0.6074 0 2.0 1e-06 
0.0 0.6075 0 2.0 1e-06 
0.0 0.6076 0 2.0 1e-06 
0.0 0.6077 0 2.0 1e-06 
0.0 0.6078 0 2.0 1e-06 
0.0 0.6079 0 2.0 1e-06 
0.0 0.608 0 2.0 1e-06 
0.0 0.6081 0 2.0 1e-06 
0.0 0.6082 0 2.0 1e-06 
0.0 0.6083 0 2.0 1e-06 
0.0 0.6084 0 2.0 1e-06 
0.0 0.6085 0 2.0 1e-06 
0.0 0.6086 0 2.0 1e-06 
0.0 0.6087 0 2.0 1e-06 
0.0 0.6088 0 2.0 1e-06 
0.0 0.6089 0 2.0 1e-06 
0.0 0.609 0 2.0 1e-06 
0.0 0.6091 0 2.0 1e-06 
0.0 0.6092 0 2.0 1e-06 
0.0 0.6093 0 2.0 1e-06 
0.0 0.6094 0 2.0 1e-06 
0.0 0.6095 0 2.0 1e-06 
0.0 0.6096 0 2.0 1e-06 
0.0 0.6097 0 2.0 1e-06 
0.0 0.6098 0 2.0 1e-06 
0.0 0.6099 0 2.0 1e-06 
0.0 0.61 0 2.0 1e-06 
0.0 0.6101 0 2.0 1e-06 
0.0 0.6102 0 2.0 1e-06 
0.0 0.6103 0 2.0 1e-06 
0.0 0.6104 0 2.0 1e-06 
0.0 0.6105 0 2.0 1e-06 
0.0 0.6106 0 2.0 1e-06 
0.0 0.6107 0 2.0 1e-06 
0.0 0.6108 0 2.0 1e-06 
0.0 0.6109 0 2.0 1e-06 
0.0 0.611 0 2.0 1e-06 
0.0 0.6111 0 2.0 1e-06 
0.0 0.6112 0 2.0 1e-06 
0.0 0.6113 0 2.0 1e-06 
0.0 0.6114 0 2.0 1e-06 
0.0 0.6115 0 2.0 1e-06 
0.0 0.6116 0 2.0 1e-06 
0.0 0.6117 0 2.0 1e-06 
0.0 0.6118 0 2.0 1e-06 
0.0 0.6119 0 2.0 1e-06 
0.0 0.612 0 2.0 1e-06 
0.0 0.6121 0 2.0 1e-06 
0.0 0.6122 0 2.0 1e-06 
0.0 0.6123 0 2.0 1e-06 
0.0 0.6124 0 2.0 1e-06 
0.0 0.6125 0 2.0 1e-06 
0.0 0.6126 0 2.0 1e-06 
0.0 0.6127 0 2.0 1e-06 
0.0 0.6128 0 2.0 1e-06 
0.0 0.6129 0 2.0 1e-06 
0.0 0.613 0 2.0 1e-06 
0.0 0.6131 0 2.0 1e-06 
0.0 0.6132 0 2.0 1e-06 
0.0 0.6133 0 2.0 1e-06 
0.0 0.6134 0 2.0 1e-06 
0.0 0.6135 0 2.0 1e-06 
0.0 0.6136 0 2.0 1e-06 
0.0 0.6137 0 2.0 1e-06 
0.0 0.6138 0 2.0 1e-06 
0.0 0.6139 0 2.0 1e-06 
0.0 0.614 0 2.0 1e-06 
0.0 0.6141 0 2.0 1e-06 
0.0 0.6142 0 2.0 1e-06 
0.0 0.6143 0 2.0 1e-06 
0.0 0.6144 0 2.0 1e-06 
0.0 0.6145 0 2.0 1e-06 
0.0 0.6146 0 2.0 1e-06 
0.0 0.6147 0 2.0 1e-06 
0.0 0.6148 0 2.0 1e-06 
0.0 0.6149 0 2.0 1e-06 
0.0 0.615 0 2.0 1e-06 
0.0 0.6151 0 2.0 1e-06 
0.0 0.6152 0 2.0 1e-06 
0.0 0.6153 0 2.0 1e-06 
0.0 0.6154 0 2.0 1e-06 
0.0 0.6155 0 2.0 1e-06 
0.0 0.6156 0 2.0 1e-06 
0.0 0.6157 0 2.0 1e-06 
0.0 0.6158 0 2.0 1e-06 
0.0 0.6159 0 2.0 1e-06 
0.0 0.616 0 2.0 1e-06 
0.0 0.6161 0 2.0 1e-06 
0.0 0.6162 0 2.0 1e-06 
0.0 0.6163 0 2.0 1e-06 
0.0 0.6164 0 2.0 1e-06 
0.0 0.6165 0 2.0 1e-06 
0.0 0.6166 0 2.0 1e-06 
0.0 0.6167 0 2.0 1e-06 
0.0 0.6168 0 2.0 1e-06 
0.0 0.6169 0 2.0 1e-06 
0.0 0.617 0 2.0 1e-06 
0.0 0.6171 0 2.0 1e-06 
0.0 0.6172 0 2.0 1e-06 
0.0 0.6173 0 2.0 1e-06 
0.0 0.6174 0 2.0 1e-06 
0.0 0.6175 0 2.0 1e-06 
0.0 0.6176 0 2.0 1e-06 
0.0 0.6177 0 2.0 1e-06 
0.0 0.6178 0 2.0 1e-06 
0.0 0.6179 0 2.0 1e-06 
0.0 0.618 0 2.0 1e-06 
0.0 0.6181 0 2.0 1e-06 
0.0 0.6182 0 2.0 1e-06 
0.0 0.6183 0 2.0 1e-06 
0.0 0.6184 0 2.0 1e-06 
0.0 0.6185 0 2.0 1e-06 
0.0 0.6186 0 2.0 1e-06 
0.0 0.6187 0 2.0 1e-06 
0.0 0.6188 0 2.0 1e-06 
0.0 0.6189 0 2.0 1e-06 
0.0 0.619 0 2.0 1e-06 
0.0 0.6191 0 2.0 1e-06 
0.0 0.6192 0 2.0 1e-06 
0.0 0.6193 0 2.0 1e-06 
0.0 0.6194 0 2.0 1e-06 
0.0 0.6195 0 2.0 1e-06 
0.0 0.6196 0 2.0 1e-06 
0.0 0.6197 0 2.0 1e-06 
0.0 0.6198 0 2.0 1e-06 
0.0 0.6199 0 2.0 1e-06 
0.0 0.62 0 2.0 1e-06 
0.0 0.6201 0 2.0 1e-06 
0.0 0.6202 0 2.0 1e-06 
0.0 0.6203 0 2.0 1e-06 
0.0 0.6204 0 2.0 1e-06 
0.0 0.6205 0 2.0 1e-06 
0.0 0.6206 0 2.0 1e-06 
0.0 0.6207 0 2.0 1e-06 
0.0 0.6208 0 2.0 1e-06 
0.0 0.6209 0 2.0 1e-06 
0.0 0.621 0 2.0 1e-06 
0.0 0.6211 0 2.0 1e-06 
0.0 0.6212 0 2.0 1e-06 
0.0 0.6213 0 2.0 1e-06 
0.0 0.6214 0 2.0 1e-06 
0.0 0.6215 0 2.0 1e-06 
0.0 0.6216 0 2.0 1e-06 
0.0 0.6217 0 2.0 1e-06 
0.0 0.6218 0 2.0 1e-06 
0.0 0.6219 0 2.0 1e-06 
0.0 0.622 0 2.0 1e-06 
0.0 0.6221 0 2.0 1e-06 
0.0 0.6222 0 2.0 1e-06 
0.0 0.6223 0 2.0 1e-06 
0.0 0.6224 0 2.0 1e-06 
0.0 0.6225 0 2.0 1e-06 
0.0 0.6226 0 2.0 1e-06 
0.0 0.6227 0 2.0 1e-06 
0.0 0.6228 0 2.0 1e-06 
0.0 0.6229 0 2.0 1e-06 
0.0 0.623 0 2.0 1e-06 
0.0 0.6231 0 2.0 1e-06 
0.0 0.6232 0 2.0 1e-06 
0.0 0.6233 0 2.0 1e-06 
0.0 0.6234 0 2.0 1e-06 
0.0 0.6235 0 2.0 1e-06 
0.0 0.6236 0 2.0 1e-06 
0.0 0.6237 0 2.0 1e-06 
0.0 0.6238 0 2.0 1e-06 
0.0 0.6239 0 2.0 1e-06 
0.0 0.624 0 2.0 1e-06 
0.0 0.6241 0 2.0 1e-06 
0.0 0.6242 0 2.0 1e-06 
0.0 0.6243 0 2.0 1e-06 
0.0 0.6244 0 2.0 1e-06 
0.0 0.6245 0 2.0 1e-06 
0.0 0.6246 0 2.0 1e-06 
0.0 0.6247 0 2.0 1e-06 
0.0 0.6248 0 2.0 1e-06 
0.0 0.6249 0 2.0 1e-06 
0.0 0.625 0 2.0 1e-06 
0.0 0.6251 0 2.0 1e-06 
0.0 0.6252 0 2.0 1e-06 
0.0 0.6253 0 2.0 1e-06 
0.0 0.6254 0 2.0 1e-06 
0.0 0.6255 0 2.0 1e-06 
0.0 0.6256 0 2.0 1e-06 
0.0 0.6257 0 2.0 1e-06 
0.0 0.6258 0 2.0 1e-06 
0.0 0.6259 0 2.0 1e-06 
0.0 0.626 0 2.0 1e-06 
0.0 0.6261 0 2.0 1e-06 
0.0 0.6262 0 2.0 1e-06 
0.0 0.6263 0 2.0 1e-06 
0.0 0.6264 0 2.0 1e-06 
0.0 0.6265 0 2.0 1e-06 
0.0 0.6266 0 2.0 1e-06 
0.0 0.6267 0 2.0 1e-06 
0.0 0.6268 0 2.0 1e-06 
0.0 0.6269 0 2.0 1e-06 
0.0 0.627 0 2.0 1e-06 
0.0 0.6271 0 2.0 1e-06 
0.0 0.6272 0 2.0 1e-06 
0.0 0.6273 0 2.0 1e-06 
0.0 0.6274 0 2.0 1e-06 
0.0 0.6275 0 2.0 1e-06 
0.0 0.6276 0 2.0 1e-06 
0.0 0.6277 0 2.0 1e-06 
0.0 0.6278 0 2.0 1e-06 
0.0 0.6279 0 2.0 1e-06 
0.0 0.628 0 2.0 1e-06 
0.0 0.6281 0 2.0 1e-06 
0.0 0.6282 0 2.0 1e-06 
0.0 0.6283 0 2.0 1e-06 
0.0 0.6284 0 2.0 1e-06 
0.0 0.6285 0 2.0 1e-06 
0.0 0.6286 0 2.0 1e-06 
0.0 0.6287 0 2.0 1e-06 
0.0 0.6288 0 2.0 1e-06 
0.0 0.6289 0 2.0 1e-06 
0.0 0.629 0 2.0 1e-06 
0.0 0.6291 0 2.0 1e-06 
0.0 0.6292 0 2.0 1e-06 
0.0 0.6293 0 2.0 1e-06 
0.0 0.6294 0 2.0 1e-06 
0.0 0.6295 0 2.0 1e-06 
0.0 0.6296 0 2.0 1e-06 
0.0 0.6297 0 2.0 1e-06 
0.0 0.6298 0 2.0 1e-06 
0.0 0.6299 0 2.0 1e-06 
0.0 0.63 0 2.0 1e-06 
0.0 0.6301 0 2.0 1e-06 
0.0 0.6302 0 2.0 1e-06 
0.0 0.6303 0 2.0 1e-06 
0.0 0.6304 0 2.0 1e-06 
0.0 0.6305 0 2.0 1e-06 
0.0 0.6306 0 2.0 1e-06 
0.0 0.6307 0 2.0 1e-06 
0.0 0.6308 0 2.0 1e-06 
0.0 0.6309 0 2.0 1e-06 
0.0 0.631 0 2.0 1e-06 
0.0 0.6311 0 2.0 1e-06 
0.0 0.6312 0 2.0 1e-06 
0.0 0.6313 0 2.0 1e-06 
0.0 0.6314 0 2.0 1e-06 
0.0 0.6315 0 2.0 1e-06 
0.0 0.6316 0 2.0 1e-06 
0.0 0.6317 0 2.0 1e-06 
0.0 0.6318 0 2.0 1e-06 
0.0 0.6319 0 2.0 1e-06 
0.0 0.632 0 2.0 1e-06 
0.0 0.6321 0 2.0 1e-06 
0.0 0.6322 0 2.0 1e-06 
0.0 0.6323 0 2.0 1e-06 
0.0 0.6324 0 2.0 1e-06 
0.0 0.6325 0 2.0 1e-06 
0.0 0.6326 0 2.0 1e-06 
0.0 0.6327 0 2.0 1e-06 
0.0 0.6328 0 2.0 1e-06 
0.0 0.6329 0 2.0 1e-06 
0.0 0.633 0 2.0 1e-06 
0.0 0.6331 0 2.0 1e-06 
0.0 0.6332 0 2.0 1e-06 
0.0 0.6333 0 2.0 1e-06 
0.0 0.6334 0 2.0 1e-06 
0.0 0.6335 0 2.0 1e-06 
0.0 0.6336 0 2.0 1e-06 
0.0 0.6337 0 2.0 1e-06 
0.0 0.6338 0 2.0 1e-06 
0.0 0.6339 0 2.0 1e-06 
0.0 0.634 0 2.0 1e-06 
0.0 0.6341 0 2.0 1e-06 
0.0 0.6342 0 2.0 1e-06 
0.0 0.6343 0 2.0 1e-06 
0.0 0.6344 0 2.0 1e-06 
0.0 0.6345 0 2.0 1e-06 
0.0 0.6346 0 2.0 1e-06 
0.0 0.6347 0 2.0 1e-06 
0.0 0.6348 0 2.0 1e-06 
0.0 0.6349 0 2.0 1e-06 
0.0 0.635 0 2.0 1e-06 
0.0 0.6351 0 2.0 1e-06 
0.0 0.6352 0 2.0 1e-06 
0.0 0.6353 0 2.0 1e-06 
0.0 0.6354 0 2.0 1e-06 
0.0 0.6355 0 2.0 1e-06 
0.0 0.6356 0 2.0 1e-06 
0.0 0.6357 0 2.0 1e-06 
0.0 0.6358 0 2.0 1e-06 
0.0 0.6359 0 2.0 1e-06 
0.0 0.636 0 2.0 1e-06 
0.0 0.6361 0 2.0 1e-06 
0.0 0.6362 0 2.0 1e-06 
0.0 0.6363 0 2.0 1e-06 
0.0 0.6364 0 2.0 1e-06 
0.0 0.6365 0 2.0 1e-06 
0.0 0.6366 0 2.0 1e-06 
0.0 0.6367 0 2.0 1e-06 
0.0 0.6368 0 2.0 1e-06 
0.0 0.6369 0 2.0 1e-06 
0.0 0.637 0 2.0 1e-06 
0.0 0.6371 0 2.0 1e-06 
0.0 0.6372 0 2.0 1e-06 
0.0 0.6373 0 2.0 1e-06 
0.0 0.6374 0 2.0 1e-06 
0.0 0.6375 0 2.0 1e-06 
0.0 0.6376 0 2.0 1e-06 
0.0 0.6377 0 2.0 1e-06 
0.0 0.6378 0 2.0 1e-06 
0.0 0.6379 0 2.0 1e-06 
0.0 0.638 0 2.0 1e-06 
0.0 0.6381 0 2.0 1e-06 
0.0 0.6382 0 2.0 1e-06 
0.0 0.6383 0 2.0 1e-06 
0.0 0.6384 0 2.0 1e-06 
0.0 0.6385 0 2.0 1e-06 
0.0 0.6386 0 2.0 1e-06 
0.0 0.6387 0 2.0 1e-06 
0.0 0.6388 0 2.0 1e-06 
0.0 0.6389 0 2.0 1e-06 
0.0 0.639 0 2.0 1e-06 
0.0 0.6391 0 2.0 1e-06 
0.0 0.6392 0 2.0 1e-06 
0.0 0.6393 0 2.0 1e-06 
0.0 0.6394 0 2.0 1e-06 
0.0 0.6395 0 2.0 1e-06 
0.0 0.6396 0 2.0 1e-06 
0.0 0.6397 0 2.0 1e-06 
0.0 0.6398 0 2.0 1e-06 
0.0 0.6399 0 2.0 1e-06 
0.0 0.64 0 2.0 1e-06 
0.0 0.6401 0 2.0 1e-06 
0.0 0.6402 0 2.0 1e-06 
0.0 0.6403 0 2.0 1e-06 
0.0 0.6404 0 2.0 1e-06 
0.0 0.6405 0 2.0 1e-06 
0.0 0.6406 0 2.0 1e-06 
0.0 0.6407 0 2.0 1e-06 
0.0 0.6408 0 2.0 1e-06 
0.0 0.6409 0 2.0 1e-06 
0.0 0.641 0 2.0 1e-06 
0.0 0.6411 0 2.0 1e-06 
0.0 0.6412 0 2.0 1e-06 
0.0 0.6413 0 2.0 1e-06 
0.0 0.6414 0 2.0 1e-06 
0.0 0.6415 0 2.0 1e-06 
0.0 0.6416 0 2.0 1e-06 
0.0 0.6417 0 2.0 1e-06 
0.0 0.6418 0 2.0 1e-06 
0.0 0.6419 0 2.0 1e-06 
0.0 0.642 0 2.0 1e-06 
0.0 0.6421 0 2.0 1e-06 
0.0 0.6422 0 2.0 1e-06 
0.0 0.6423 0 2.0 1e-06 
0.0 0.6424 0 2.0 1e-06 
0.0 0.6425 0 2.0 1e-06 
0.0 0.6426 0 2.0 1e-06 
0.0 0.6427 0 2.0 1e-06 
0.0 0.6428 0 2.0 1e-06 
0.0 0.6429 0 2.0 1e-06 
0.0 0.643 0 2.0 1e-06 
0.0 0.6431 0 2.0 1e-06 
0.0 0.6432 0 2.0 1e-06 
0.0 0.6433 0 2.0 1e-06 
0.0 0.6434 0 2.0 1e-06 
0.0 0.6435 0 2.0 1e-06 
0.0 0.6436 0 2.0 1e-06 
0.0 0.6437 0 2.0 1e-06 
0.0 0.6438 0 2.0 1e-06 
0.0 0.6439 0 2.0 1e-06 
0.0 0.644 0 2.0 1e-06 
0.0 0.6441 0 2.0 1e-06 
0.0 0.6442 0 2.0 1e-06 
0.0 0.6443 0 2.0 1e-06 
0.0 0.6444 0 2.0 1e-06 
0.0 0.6445 0 2.0 1e-06 
0.0 0.6446 0 2.0 1e-06 
0.0 0.6447 0 2.0 1e-06 
0.0 0.6448 0 2.0 1e-06 
0.0 0.6449 0 2.0 1e-06 
0.0 0.645 0 2.0 1e-06 
0.0 0.6451 0 2.0 1e-06 
0.0 0.6452 0 2.0 1e-06 
0.0 0.6453 0 2.0 1e-06 
0.0 0.6454 0 2.0 1e-06 
0.0 0.6455 0 2.0 1e-06 
0.0 0.6456 0 2.0 1e-06 
0.0 0.6457 0 2.0 1e-06 
0.0 0.6458 0 2.0 1e-06 
0.0 0.6459 0 2.0 1e-06 
0.0 0.646 0 2.0 1e-06 
0.0 0.6461 0 2.0 1e-06 
0.0 0.6462 0 2.0 1e-06 
0.0 0.6463 0 2.0 1e-06 
0.0 0.6464 0 2.0 1e-06 
0.0 0.6465 0 2.0 1e-06 
0.0 0.6466 0 2.0 1e-06 
0.0 0.6467 0 2.0 1e-06 
0.0 0.6468 0 2.0 1e-06 
0.0 0.6469 0 2.0 1e-06 
0.0 0.647 0 2.0 1e-06 
0.0 0.6471 0 2.0 1e-06 
0.0 0.6472 0 2.0 1e-06 
0.0 0.6473 0 2.0 1e-06 
0.0 0.6474 0 2.0 1e-06 
0.0 0.6475 0 2.0 1e-06 
0.0 0.6476 0 2.0 1e-06 
0.0 0.6477 0 2.0 1e-06 
0.0 0.6478 0 2.0 1e-06 
0.0 0.6479 0 2.0 1e-06 
0.0 0.648 0 2.0 1e-06 
0.0 0.6481 0 2.0 1e-06 
0.0 0.6482 0 2.0 1e-06 
0.0 0.6483 0 2.0 1e-06 
0.0 0.6484 0 2.0 1e-06 
0.0 0.6485 0 2.0 1e-06 
0.0 0.6486 0 2.0 1e-06 
0.0 0.6487 0 2.0 1e-06 
0.0 0.6488 0 2.0 1e-06 
0.0 0.6489 0 2.0 1e-06 
0.0 0.649 0 2.0 1e-06 
0.0 0.6491 0 2.0 1e-06 
0.0 0.6492 0 2.0 1e-06 
0.0 0.6493 0 2.0 1e-06 
0.0 0.6494 0 2.0 1e-06 
0.0 0.6495 0 2.0 1e-06 
0.0 0.6496 0 2.0 1e-06 
0.0 0.6497 0 2.0 1e-06 
0.0 0.6498 0 2.0 1e-06 
0.0 0.6499 0 2.0 1e-06 
0.0 0.65 0 2.0 1e-06 
0.0 0.6501 0 2.0 1e-06 
0.0 0.6502 0 2.0 1e-06 
0.0 0.6503 0 2.0 1e-06 
0.0 0.6504 0 2.0 1e-06 
0.0 0.6505 0 2.0 1e-06 
0.0 0.6506 0 2.0 1e-06 
0.0 0.6507 0 2.0 1e-06 
0.0 0.6508 0 2.0 1e-06 
0.0 0.6509 0 2.0 1e-06 
0.0 0.651 0 2.0 1e-06 
0.0 0.6511 0 2.0 1e-06 
0.0 0.6512 0 2.0 1e-06 
0.0 0.6513 0 2.0 1e-06 
0.0 0.6514 0 2.0 1e-06 
0.0 0.6515 0 2.0 1e-06 
0.0 0.6516 0 2.0 1e-06 
0.0 0.6517 0 2.0 1e-06 
0.0 0.6518 0 2.0 1e-06 
0.0 0.6519 0 2.0 1e-06 
0.0 0.652 0 2.0 1e-06 
0.0 0.6521 0 2.0 1e-06 
0.0 0.6522 0 2.0 1e-06 
0.0 0.6523 0 2.0 1e-06 
0.0 0.6524 0 2.0 1e-06 
0.0 0.6525 0 2.0 1e-06 
0.0 0.6526 0 2.0 1e-06 
0.0 0.6527 0 2.0 1e-06 
0.0 0.6528 0 2.0 1e-06 
0.0 0.6529 0 2.0 1e-06 
0.0 0.653 0 2.0 1e-06 
0.0 0.6531 0 2.0 1e-06 
0.0 0.6532 0 2.0 1e-06 
0.0 0.6533 0 2.0 1e-06 
0.0 0.6534 0 2.0 1e-06 
0.0 0.6535 0 2.0 1e-06 
0.0 0.6536 0 2.0 1e-06 
0.0 0.6537 0 2.0 1e-06 
0.0 0.6538 0 2.0 1e-06 
0.0 0.6539 0 2.0 1e-06 
0.0 0.654 0 2.0 1e-06 
0.0 0.6541 0 2.0 1e-06 
0.0 0.6542 0 2.0 1e-06 
0.0 0.6543 0 2.0 1e-06 
0.0 0.6544 0 2.0 1e-06 
0.0 0.6545 0 2.0 1e-06 
0.0 0.6546 0 2.0 1e-06 
0.0 0.6547 0 2.0 1e-06 
0.0 0.6548 0 2.0 1e-06 
0.0 0.6549 0 2.0 1e-06 
0.0 0.655 0 2.0 1e-06 
0.0 0.6551 0 2.0 1e-06 
0.0 0.6552 0 2.0 1e-06 
0.0 0.6553 0 2.0 1e-06 
0.0 0.6554 0 2.0 1e-06 
0.0 0.6555 0 2.0 1e-06 
0.0 0.6556 0 2.0 1e-06 
0.0 0.6557 0 2.0 1e-06 
0.0 0.6558 0 2.0 1e-06 
0.0 0.6559 0 2.0 1e-06 
0.0 0.656 0 2.0 1e-06 
0.0 0.6561 0 2.0 1e-06 
0.0 0.6562 0 2.0 1e-06 
0.0 0.6563 0 2.0 1e-06 
0.0 0.6564 0 2.0 1e-06 
0.0 0.6565 0 2.0 1e-06 
0.0 0.6566 0 2.0 1e-06 
0.0 0.6567 0 2.0 1e-06 
0.0 0.6568 0 2.0 1e-06 
0.0 0.6569 0 2.0 1e-06 
0.0 0.657 0 2.0 1e-06 
0.0 0.6571 0 2.0 1e-06 
0.0 0.6572 0 2.0 1e-06 
0.0 0.6573 0 2.0 1e-06 
0.0 0.6574 0 2.0 1e-06 
0.0 0.6575 0 2.0 1e-06 
0.0 0.6576 0 2.0 1e-06 
0.0 0.6577 0 2.0 1e-06 
0.0 0.6578 0 2.0 1e-06 
0.0 0.6579 0 2.0 1e-06 
0.0 0.658 0 2.0 1e-06 
0.0 0.6581 0 2.0 1e-06 
0.0 0.6582 0 2.0 1e-06 
0.0 0.6583 0 2.0 1e-06 
0.0 0.6584 0 2.0 1e-06 
0.0 0.6585 0 2.0 1e-06 
0.0 0.6586 0 2.0 1e-06 
0.0 0.6587 0 2.0 1e-06 
0.0 0.6588 0 2.0 1e-06 
0.0 0.6589 0 2.0 1e-06 
0.0 0.659 0 2.0 1e-06 
0.0 0.6591 0 2.0 1e-06 
0.0 0.6592 0 2.0 1e-06 
0.0 0.6593 0 2.0 1e-06 
0.0 0.6594 0 2.0 1e-06 
0.0 0.6595 0 2.0 1e-06 
0.0 0.6596 0 2.0 1e-06 
0.0 0.6597 0 2.0 1e-06 
0.0 0.6598 0 2.0 1e-06 
0.0 0.6599 0 2.0 1e-06 
0.0 0.66 0 2.0 1e-06 
0.0 0.6601 0 2.0 1e-06 
0.0 0.6602 0 2.0 1e-06 
0.0 0.6603 0 2.0 1e-06 
0.0 0.6604 0 2.0 1e-06 
0.0 0.6605 0 2.0 1e-06 
0.0 0.6606 0 2.0 1e-06 
0.0 0.6607 0 2.0 1e-06 
0.0 0.6608 0 2.0 1e-06 
0.0 0.6609 0 2.0 1e-06 
0.0 0.661 0 2.0 1e-06 
0.0 0.6611 0 2.0 1e-06 
0.0 0.6612 0 2.0 1e-06 
0.0 0.6613 0 2.0 1e-06 
0.0 0.6614 0 2.0 1e-06 
0.0 0.6615 0 2.0 1e-06 
0.0 0.6616 0 2.0 1e-06 
0.0 0.6617 0 2.0 1e-06 
0.0 0.6618 0 2.0 1e-06 
0.0 0.6619 0 2.0 1e-06 
0.0 0.662 0 2.0 1e-06 
0.0 0.6621 0 2.0 1e-06 
0.0 0.6622 0 2.0 1e-06 
0.0 0.6623 0 2.0 1e-06 
0.0 0.6624 0 2.0 1e-06 
0.0 0.6625 0 2.0 1e-06 
0.0 0.6626 0 2.0 1e-06 
0.0 0.6627 0 2.0 1e-06 
0.0 0.6628 0 2.0 1e-06 
0.0 0.6629 0 2.0 1e-06 
0.0 0.663 0 2.0 1e-06 
0.0 0.6631 0 2.0 1e-06 
0.0 0.6632 0 2.0 1e-06 
0.0 0.6633 0 2.0 1e-06 
0.0 0.6634 0 2.0 1e-06 
0.0 0.6635 0 2.0 1e-06 
0.0 0.6636 0 2.0 1e-06 
0.0 0.6637 0 2.0 1e-06 
0.0 0.6638 0 2.0 1e-06 
0.0 0.6639 0 2.0 1e-06 
0.0 0.664 0 2.0 1e-06 
0.0 0.6641 0 2.0 1e-06 
0.0 0.6642 0 2.0 1e-06 
0.0 0.6643 0 2.0 1e-06 
0.0 0.6644 0 2.0 1e-06 
0.0 0.6645 0 2.0 1e-06 
0.0 0.6646 0 2.0 1e-06 
0.0 0.6647 0 2.0 1e-06 
0.0 0.6648 0 2.0 1e-06 
0.0 0.6649 0 2.0 1e-06 
0.0 0.665 0 2.0 1e-06 
0.0 0.6651 0 2.0 1e-06 
0.0 0.6652 0 2.0 1e-06 
0.0 0.6653 0 2.0 1e-06 
0.0 0.6654 0 2.0 1e-06 
0.0 0.6655 0 2.0 1e-06 
0.0 0.6656 0 2.0 1e-06 
0.0 0.6657 0 2.0 1e-06 
0.0 0.6658 0 2.0 1e-06 
0.0 0.6659 0 2.0 1e-06 
0.0 0.666 0 2.0 1e-06 
0.0 0.6661 0 2.0 1e-06 
0.0 0.6662 0 2.0 1e-06 
0.0 0.6663 0 2.0 1e-06 
0.0 0.6664 0 2.0 1e-06 
0.0 0.6665 0 2.0 1e-06 
0.0 0.6666 0 2.0 1e-06 
0.0 0.6667 0 2.0 1e-06 
0.0 0.6668 0 2.0 1e-06 
0.0 0.6669 0 2.0 1e-06 
0.0 0.667 0 2.0 1e-06 
0.0 0.6671 0 2.0 1e-06 
0.0 0.6672 0 2.0 1e-06 
0.0 0.6673 0 2.0 1e-06 
0.0 0.6674 0 2.0 1e-06 
0.0 0.6675 0 2.0 1e-06 
0.0 0.6676 0 2.0 1e-06 
0.0 0.6677 0 2.0 1e-06 
0.0 0.6678 0 2.0 1e-06 
0.0 0.6679 0 2.0 1e-06 
0.0 0.668 0 2.0 1e-06 
0.0 0.6681 0 2.0 1e-06 
0.0 0.6682 0 2.0 1e-06 
0.0 0.6683 0 2.0 1e-06 
0.0 0.6684 0 2.0 1e-06 
0.0 0.6685 0 2.0 1e-06 
0.0 0.6686 0 2.0 1e-06 
0.0 0.6687 0 2.0 1e-06 
0.0 0.6688 0 2.0 1e-06 
0.0 0.6689 0 2.0 1e-06 
0.0 0.669 0 2.0 1e-06 
0.0 0.6691 0 2.0 1e-06 
0.0 0.6692 0 2.0 1e-06 
0.0 0.6693 0 2.0 1e-06 
0.0 0.6694 0 2.0 1e-06 
0.0 0.6695 0 2.0 1e-06 
0.0 0.6696 0 2.0 1e-06 
0.0 0.6697 0 2.0 1e-06 
0.0 0.6698 0 2.0 1e-06 
0.0 0.6699 0 2.0 1e-06 
0.0 0.67 0 2.0 1e-06 
0.0 0.6701 0 2.0 1e-06 
0.0 0.6702 0 2.0 1e-06 
0.0 0.6703 0 2.0 1e-06 
0.0 0.6704 0 2.0 1e-06 
0.0 0.6705 0 2.0 1e-06 
0.0 0.6706 0 2.0 1e-06 
0.0 0.6707 0 2.0 1e-06 
0.0 0.6708 0 2.0 1e-06 
0.0 0.6709 0 2.0 1e-06 
0.0 0.671 0 2.0 1e-06 
0.0 0.6711 0 2.0 1e-06 
0.0 0.6712 0 2.0 1e-06 
0.0 0.6713 0 2.0 1e-06 
0.0 0.6714 0 2.0 1e-06 
0.0 0.6715 0 2.0 1e-06 
0.0 0.6716 0 2.0 1e-06 
0.0 0.6717 0 2.0 1e-06 
0.0 0.6718 0 2.0 1e-06 
0.0 0.6719 0 2.0 1e-06 
0.0 0.672 0 2.0 1e-06 
0.0 0.6721 0 2.0 1e-06 
0.0 0.6722 0 2.0 1e-06 
0.0 0.6723 0 2.0 1e-06 
0.0 0.6724 0 2.0 1e-06 
0.0 0.6725 0 2.0 1e-06 
0.0 0.6726 0 2.0 1e-06 
0.0 0.6727 0 2.0 1e-06 
0.0 0.6728 0 2.0 1e-06 
0.0 0.6729 0 2.0 1e-06 
0.0 0.673 0 2.0 1e-06 
0.0 0.6731 0 2.0 1e-06 
0.0 0.6732 0 2.0 1e-06 
0.0 0.6733 0 2.0 1e-06 
0.0 0.6734 0 2.0 1e-06 
0.0 0.6735 0 2.0 1e-06 
0.0 0.6736 0 2.0 1e-06 
0.0 0.6737 0 2.0 1e-06 
0.0 0.6738 0 2.0 1e-06 
0.0 0.6739 0 2.0 1e-06 
0.0 0.674 0 2.0 1e-06 
0.0 0.6741 0 2.0 1e-06 
0.0 0.6742 0 2.0 1e-06 
0.0 0.6743 0 2.0 1e-06 
0.0 0.6744 0 2.0 1e-06 
0.0 0.6745 0 2.0 1e-06 
0.0 0.6746 0 2.0 1e-06 
0.0 0.6747 0 2.0 1e-06 
0.0 0.6748 0 2.0 1e-06 
0.0 0.6749 0 2.0 1e-06 
0.0 0.675 0 2.0 1e-06 
0.0 0.6751 0 2.0 1e-06 
0.0 0.6752 0 2.0 1e-06 
0.0 0.6753 0 2.0 1e-06 
0.0 0.6754 0 2.0 1e-06 
0.0 0.6755 0 2.0 1e-06 
0.0 0.6756 0 2.0 1e-06 
0.0 0.6757 0 2.0 1e-06 
0.0 0.6758 0 2.0 1e-06 
0.0 0.6759 0 2.0 1e-06 
0.0 0.676 0 2.0 1e-06 
0.0 0.6761 0 2.0 1e-06 
0.0 0.6762 0 2.0 1e-06 
0.0 0.6763 0 2.0 1e-06 
0.0 0.6764 0 2.0 1e-06 
0.0 0.6765 0 2.0 1e-06 
0.0 0.6766 0 2.0 1e-06 
0.0 0.6767 0 2.0 1e-06 
0.0 0.6768 0 2.0 1e-06 
0.0 0.6769 0 2.0 1e-06 
0.0 0.677 0 2.0 1e-06 
0.0 0.6771 0 2.0 1e-06 
0.0 0.6772 0 2.0 1e-06 
0.0 0.6773 0 2.0 1e-06 
0.0 0.6774 0 2.0 1e-06 
0.0 0.6775 0 2.0 1e-06 
0.0 0.6776 0 2.0 1e-06 
0.0 0.6777 0 2.0 1e-06 
0.0 0.6778 0 2.0 1e-06 
0.0 0.6779 0 2.0 1e-06 
0.0 0.678 0 2.0 1e-06 
0.0 0.6781 0 2.0 1e-06 
0.0 0.6782 0 2.0 1e-06 
0.0 0.6783 0 2.0 1e-06 
0.0 0.6784 0 2.0 1e-06 
0.0 0.6785 0 2.0 1e-06 
0.0 0.6786 0 2.0 1e-06 
0.0 0.6787 0 2.0 1e-06 
0.0 0.6788 0 2.0 1e-06 
0.0 0.6789 0 2.0 1e-06 
0.0 0.679 0 2.0 1e-06 
0.0 0.6791 0 2.0 1e-06 
0.0 0.6792 0 2.0 1e-06 
0.0 0.6793 0 2.0 1e-06 
0.0 0.6794 0 2.0 1e-06 
0.0 0.6795 0 2.0 1e-06 
0.0 0.6796 0 2.0 1e-06 
0.0 0.6797 0 2.0 1e-06 
0.0 0.6798 0 2.0 1e-06 
0.0 0.6799 0 2.0 1e-06 
0.0 0.68 0 2.0 1e-06 
0.0 0.6801 0 2.0 1e-06 
0.0 0.6802 0 2.0 1e-06 
0.0 0.6803 0 2.0 1e-06 
0.0 0.6804 0 2.0 1e-06 
0.0 0.6805 0 2.0 1e-06 
0.0 0.6806 0 2.0 1e-06 
0.0 0.6807 0 2.0 1e-06 
0.0 0.6808 0 2.0 1e-06 
0.0 0.6809 0 2.0 1e-06 
0.0 0.681 0 2.0 1e-06 
0.0 0.6811 0 2.0 1e-06 
0.0 0.6812 0 2.0 1e-06 
0.0 0.6813 0 2.0 1e-06 
0.0 0.6814 0 2.0 1e-06 
0.0 0.6815 0 2.0 1e-06 
0.0 0.6816 0 2.0 1e-06 
0.0 0.6817 0 2.0 1e-06 
0.0 0.6818 0 2.0 1e-06 
0.0 0.6819 0 2.0 1e-06 
0.0 0.682 0 2.0 1e-06 
0.0 0.6821 0 2.0 1e-06 
0.0 0.6822 0 2.0 1e-06 
0.0 0.6823 0 2.0 1e-06 
0.0 0.6824 0 2.0 1e-06 
0.0 0.6825 0 2.0 1e-06 
0.0 0.6826 0 2.0 1e-06 
0.0 0.6827 0 2.0 1e-06 
0.0 0.6828 0 2.0 1e-06 
0.0 0.6829 0 2.0 1e-06 
0.0 0.683 0 2.0 1e-06 
0.0 0.6831 0 2.0 1e-06 
0.0 0.6832 0 2.0 1e-06 
0.0 0.6833 0 2.0 1e-06 
0.0 0.6834 0 2.0 1e-06 
0.0 0.6835 0 2.0 1e-06 
0.0 0.6836 0 2.0 1e-06 
0.0 0.6837 0 2.0 1e-06 
0.0 0.6838 0 2.0 1e-06 
0.0 0.6839 0 2.0 1e-06 
0.0 0.684 0 2.0 1e-06 
0.0 0.6841 0 2.0 1e-06 
0.0 0.6842 0 2.0 1e-06 
0.0 0.6843 0 2.0 1e-06 
0.0 0.6844 0 2.0 1e-06 
0.0 0.6845 0 2.0 1e-06 
0.0 0.6846 0 2.0 1e-06 
0.0 0.6847 0 2.0 1e-06 
0.0 0.6848 0 2.0 1e-06 
0.0 0.6849 0 2.0 1e-06 
0.0 0.685 0 2.0 1e-06 
0.0 0.6851 0 2.0 1e-06 
0.0 0.6852 0 2.0 1e-06 
0.0 0.6853 0 2.0 1e-06 
0.0 0.6854 0 2.0 1e-06 
0.0 0.6855 0 2.0 1e-06 
0.0 0.6856 0 2.0 1e-06 
0.0 0.6857 0 2.0 1e-06 
0.0 0.6858 0 2.0 1e-06 
0.0 0.6859 0 2.0 1e-06 
0.0 0.686 0 2.0 1e-06 
0.0 0.6861 0 2.0 1e-06 
0.0 0.6862 0 2.0 1e-06 
0.0 0.6863 0 2.0 1e-06 
0.0 0.6864 0 2.0 1e-06 
0.0 0.6865 0 2.0 1e-06 
0.0 0.6866 0 2.0 1e-06 
0.0 0.6867 0 2.0 1e-06 
0.0 0.6868 0 2.0 1e-06 
0.0 0.6869 0 2.0 1e-06 
0.0 0.687 0 2.0 1e-06 
0.0 0.6871 0 2.0 1e-06 
0.0 0.6872 0 2.0 1e-06 
0.0 0.6873 0 2.0 1e-06 
0.0 0.6874 0 2.0 1e-06 
0.0 0.6875 0 2.0 1e-06 
0.0 0.6876 0 2.0 1e-06 
0.0 0.6877 0 2.0 1e-06 
0.0 0.6878 0 2.0 1e-06 
0.0 0.6879 0 2.0 1e-06 
0.0 0.688 0 2.0 1e-06 
0.0 0.6881 0 2.0 1e-06 
0.0 0.6882 0 2.0 1e-06 
0.0 0.6883 0 2.0 1e-06 
0.0 0.6884 0 2.0 1e-06 
0.0 0.6885 0 2.0 1e-06 
0.0 0.6886 0 2.0 1e-06 
0.0 0.6887 0 2.0 1e-06 
0.0 0.6888 0 2.0 1e-06 
0.0 0.6889 0 2.0 1e-06 
0.0 0.689 0 2.0 1e-06 
0.0 0.6891 0 2.0 1e-06 
0.0 0.6892 0 2.0 1e-06 
0.0 0.6893 0 2.0 1e-06 
0.0 0.6894 0 2.0 1e-06 
0.0 0.6895 0 2.0 1e-06 
0.0 0.6896 0 2.0 1e-06 
0.0 0.6897 0 2.0 1e-06 
0.0 0.6898 0 2.0 1e-06 
0.0 0.6899 0 2.0 1e-06 
0.0 0.69 0 2.0 1e-06 
0.0 0.6901 0 2.0 1e-06 
0.0 0.6902 0 2.0 1e-06 
0.0 0.6903 0 2.0 1e-06 
0.0 0.6904 0 2.0 1e-06 
0.0 0.6905 0 2.0 1e-06 
0.0 0.6906 0 2.0 1e-06 
0.0 0.6907 0 2.0 1e-06 
0.0 0.6908 0 2.0 1e-06 
0.0 0.6909 0 2.0 1e-06 
0.0 0.691 0 2.0 1e-06 
0.0 0.6911 0 2.0 1e-06 
0.0 0.6912 0 2.0 1e-06 
0.0 0.6913 0 2.0 1e-06 
0.0 0.6914 0 2.0 1e-06 
0.0 0.6915 0 2.0 1e-06 
0.0 0.6916 0 2.0 1e-06 
0.0 0.6917 0 2.0 1e-06 
0.0 0.6918 0 2.0 1e-06 
0.0 0.6919 0 2.0 1e-06 
0.0 0.692 0 2.0 1e-06 
0.0 0.6921 0 2.0 1e-06 
0.0 0.6922 0 2.0 1e-06 
0.0 0.6923 0 2.0 1e-06 
0.0 0.6924 0 2.0 1e-06 
0.0 0.6925 0 2.0 1e-06 
0.0 0.6926 0 2.0 1e-06 
0.0 0.6927 0 2.0 1e-06 
0.0 0.6928 0 2.0 1e-06 
0.0 0.6929 0 2.0 1e-06 
0.0 0.693 0 2.0 1e-06 
0.0 0.6931 0 2.0 1e-06 
0.0 0.6932 0 2.0 1e-06 
0.0 0.6933 0 2.0 1e-06 
0.0 0.6934 0 2.0 1e-06 
0.0 0.6935 0 2.0 1e-06 
0.0 0.6936 0 2.0 1e-06 
0.0 0.6937 0 2.0 1e-06 
0.0 0.6938 0 2.0 1e-06 
0.0 0.6939 0 2.0 1e-06 
0.0 0.694 0 2.0 1e-06 
0.0 0.6941 0 2.0 1e-06 
0.0 0.6942 0 2.0 1e-06 
0.0 0.6943 0 2.0 1e-06 
0.0 0.6944 0 2.0 1e-06 
0.0 0.6945 0 2.0 1e-06 
0.0 0.6946 0 2.0 1e-06 
0.0 0.6947 0 2.0 1e-06 
0.0 0.6948 0 2.0 1e-06 
0.0 0.6949 0 2.0 1e-06 
0.0 0.695 0 2.0 1e-06 
0.0 0.6951 0 2.0 1e-06 
0.0 0.6952 0 2.0 1e-06 
0.0 0.6953 0 2.0 1e-06 
0.0 0.6954 0 2.0 1e-06 
0.0 0.6955 0 2.0 1e-06 
0.0 0.6956 0 2.0 1e-06 
0.0 0.6957 0 2.0 1e-06 
0.0 0.6958 0 2.0 1e-06 
0.0 0.6959 0 2.0 1e-06 
0.0 0.696 0 2.0 1e-06 
0.0 0.6961 0 2.0 1e-06 
0.0 0.6962 0 2.0 1e-06 
0.0 0.6963 0 2.0 1e-06 
0.0 0.6964 0 2.0 1e-06 
0.0 0.6965 0 2.0 1e-06 
0.0 0.6966 0 2.0 1e-06 
0.0 0.6967 0 2.0 1e-06 
0.0 0.6968 0 2.0 1e-06 
0.0 0.6969 0 2.0 1e-06 
0.0 0.697 0 2.0 1e-06 
0.0 0.6971 0 2.0 1e-06 
0.0 0.6972 0 2.0 1e-06 
0.0 0.6973 0 2.0 1e-06 
0.0 0.6974 0 2.0 1e-06 
0.0 0.6975 0 2.0 1e-06 
0.0 0.6976 0 2.0 1e-06 
0.0 0.6977 0 2.0 1e-06 
0.0 0.6978 0 2.0 1e-06 
0.0 0.6979 0 2.0 1e-06 
0.0 0.698 0 2.0 1e-06 
0.0 0.6981 0 2.0 1e-06 
0.0 0.6982 0 2.0 1e-06 
0.0 0.6983 0 2.0 1e-06 
0.0 0.6984 0 2.0 1e-06 
0.0 0.6985 0 2.0 1e-06 
0.0 0.6986 0 2.0 1e-06 
0.0 0.6987 0 2.0 1e-06 
0.0 0.6988 0 2.0 1e-06 
0.0 0.6989 0 2.0 1e-06 
0.0 0.699 0 2.0 1e-06 
0.0 0.6991 0 2.0 1e-06 
0.0 0.6992 0 2.0 1e-06 
0.0 0.6993 0 2.0 1e-06 
0.0 0.6994 0 2.0 1e-06 
0.0 0.6995 0 2.0 1e-06 
0.0 0.6996 0 2.0 1e-06 
0.0 0.6997 0 2.0 1e-06 
0.0 0.6998 0 2.0 1e-06 
0.0 0.6999 0 2.0 1e-06 
0.0 0.7 0 2.0 1e-06 
0.0 0.7001 0 2.0 1e-06 
0.0 0.7002 0 2.0 1e-06 
0.0 0.7003 0 2.0 1e-06 
0.0 0.7004 0 2.0 1e-06 
0.0 0.7005 0 2.0 1e-06 
0.0 0.7006 0 2.0 1e-06 
0.0 0.7007 0 2.0 1e-06 
0.0 0.7008 0 2.0 1e-06 
0.0 0.7009 0 2.0 1e-06 
0.0 0.701 0 2.0 1e-06 
0.0 0.7011 0 2.0 1e-06 
0.0 0.7012 0 2.0 1e-06 
0.0 0.7013 0 2.0 1e-06 
0.0 0.7014 0 2.0 1e-06 
0.0 0.7015 0 2.0 1e-06 
0.0 0.7016 0 2.0 1e-06 
0.0 0.7017 0 2.0 1e-06 
0.0 0.7018 0 2.0 1e-06 
0.0 0.7019 0 2.0 1e-06 
0.0 0.702 0 2.0 1e-06 
0.0 0.7021 0 2.0 1e-06 
0.0 0.7022 0 2.0 1e-06 
0.0 0.7023 0 2.0 1e-06 
0.0 0.7024 0 2.0 1e-06 
0.0 0.7025 0 2.0 1e-06 
0.0 0.7026 0 2.0 1e-06 
0.0 0.7027 0 2.0 1e-06 
0.0 0.7028 0 2.0 1e-06 
0.0 0.7029 0 2.0 1e-06 
0.0 0.703 0 2.0 1e-06 
0.0 0.7031 0 2.0 1e-06 
0.0 0.7032 0 2.0 1e-06 
0.0 0.7033 0 2.0 1e-06 
0.0 0.7034 0 2.0 1e-06 
0.0 0.7035 0 2.0 1e-06 
0.0 0.7036 0 2.0 1e-06 
0.0 0.7037 0 2.0 1e-06 
0.0 0.7038 0 2.0 1e-06 
0.0 0.7039 0 2.0 1e-06 
0.0 0.704 0 2.0 1e-06 
0.0 0.7041 0 2.0 1e-06 
0.0 0.7042 0 2.0 1e-06 
0.0 0.7043 0 2.0 1e-06 
0.0 0.7044 0 2.0 1e-06 
0.0 0.7045 0 2.0 1e-06 
0.0 0.7046 0 2.0 1e-06 
0.0 0.7047 0 2.0 1e-06 
0.0 0.7048 0 2.0 1e-06 
0.0 0.7049 0 2.0 1e-06 
0.0 0.705 0 2.0 1e-06 
0.0 0.7051 0 2.0 1e-06 
0.0 0.7052 0 2.0 1e-06 
0.0 0.7053 0 2.0 1e-06 
0.0 0.7054 0 2.0 1e-06 
0.0 0.7055 0 2.0 1e-06 
0.0 0.7056 0 2.0 1e-06 
0.0 0.7057 0 2.0 1e-06 
0.0 0.7058 0 2.0 1e-06 
0.0 0.7059 0 2.0 1e-06 
0.0 0.706 0 2.0 1e-06 
0.0 0.7061 0 2.0 1e-06 
0.0 0.7062 0 2.0 1e-06 
0.0 0.7063 0 2.0 1e-06 
0.0 0.7064 0 2.0 1e-06 
0.0 0.7065 0 2.0 1e-06 
0.0 0.7066 0 2.0 1e-06 
0.0 0.7067 0 2.0 1e-06 
0.0 0.7068 0 2.0 1e-06 
0.0 0.7069 0 2.0 1e-06 
0.0 0.707 0 2.0 1e-06 
0.0 0.7071 0 2.0 1e-06 
0.0 0.7072 0 2.0 1e-06 
0.0 0.7073 0 2.0 1e-06 
0.0 0.7074 0 2.0 1e-06 
0.0 0.7075 0 2.0 1e-06 
0.0 0.7076 0 2.0 1e-06 
0.0 0.7077 0 2.0 1e-06 
0.0 0.7078 0 2.0 1e-06 
0.0 0.7079 0 2.0 1e-06 
0.0 0.708 0 2.0 1e-06 
0.0 0.7081 0 2.0 1e-06 
0.0 0.7082 0 2.0 1e-06 
0.0 0.7083 0 2.0 1e-06 
0.0 0.7084 0 2.0 1e-06 
0.0 0.7085 0 2.0 1e-06 
0.0 0.7086 0 2.0 1e-06 
0.0 0.7087 0 2.0 1e-06 
0.0 0.7088 0 2.0 1e-06 
0.0 0.7089 0 2.0 1e-06 
0.0 0.709 0 2.0 1e-06 
0.0 0.7091 0 2.0 1e-06 
0.0 0.7092 0 2.0 1e-06 
0.0 0.7093 0 2.0 1e-06 
0.0 0.7094 0 2.0 1e-06 
0.0 0.7095 0 2.0 1e-06 
0.0 0.7096 0 2.0 1e-06 
0.0 0.7097 0 2.0 1e-06 
0.0 0.7098 0 2.0 1e-06 
0.0 0.7099 0 2.0 1e-06 
0.0 0.71 0 2.0 1e-06 
0.0 0.7101 0 2.0 1e-06 
0.0 0.7102 0 2.0 1e-06 
0.0 0.7103 0 2.0 1e-06 
0.0 0.7104 0 2.0 1e-06 
0.0 0.7105 0 2.0 1e-06 
0.0 0.7106 0 2.0 1e-06 
0.0 0.7107 0 2.0 1e-06 
0.0 0.7108 0 2.0 1e-06 
0.0 0.7109 0 2.0 1e-06 
0.0 0.711 0 2.0 1e-06 
0.0 0.7111 0 2.0 1e-06 
0.0 0.7112 0 2.0 1e-06 
0.0 0.7113 0 2.0 1e-06 
0.0 0.7114 0 2.0 1e-06 
0.0 0.7115 0 2.0 1e-06 
0.0 0.7116 0 2.0 1e-06 
0.0 0.7117 0 2.0 1e-06 
0.0 0.7118 0 2.0 1e-06 
0.0 0.7119 0 2.0 1e-06 
0.0 0.712 0 2.0 1e-06 
0.0 0.7121 0 2.0 1e-06 
0.0 0.7122 0 2.0 1e-06 
0.0 0.7123 0 2.0 1e-06 
0.0 0.7124 0 2.0 1e-06 
0.0 0.7125 0 2.0 1e-06 
0.0 0.7126 0 2.0 1e-06 
0.0 0.7127 0 2.0 1e-06 
0.0 0.7128 0 2.0 1e-06 
0.0 0.7129 0 2.0 1e-06 
0.0 0.713 0 2.0 1e-06 
0.0 0.7131 0 2.0 1e-06 
0.0 0.7132 0 2.0 1e-06 
0.0 0.7133 0 2.0 1e-06 
0.0 0.7134 0 2.0 1e-06 
0.0 0.7135 0 2.0 1e-06 
0.0 0.7136 0 2.0 1e-06 
0.0 0.7137 0 2.0 1e-06 
0.0 0.7138 0 2.0 1e-06 
0.0 0.7139 0 2.0 1e-06 
0.0 0.714 0 2.0 1e-06 
0.0 0.7141 0 2.0 1e-06 
0.0 0.7142 0 2.0 1e-06 
0.0 0.7143 0 2.0 1e-06 
0.0 0.7144 0 2.0 1e-06 
0.0 0.7145 0 2.0 1e-06 
0.0 0.7146 0 2.0 1e-06 
0.0 0.7147 0 2.0 1e-06 
0.0 0.7148 0 2.0 1e-06 
0.0 0.7149 0 2.0 1e-06 
0.0 0.715 0 2.0 1e-06 
0.0 0.7151 0 2.0 1e-06 
0.0 0.7152 0 2.0 1e-06 
0.0 0.7153 0 2.0 1e-06 
0.0 0.7154 0 2.0 1e-06 
0.0 0.7155 0 2.0 1e-06 
0.0 0.7156 0 2.0 1e-06 
0.0 0.7157 0 2.0 1e-06 
0.0 0.7158 0 2.0 1e-06 
0.0 0.7159 0 2.0 1e-06 
0.0 0.716 0 2.0 1e-06 
0.0 0.7161 0 2.0 1e-06 
0.0 0.7162 0 2.0 1e-06 
0.0 0.7163 0 2.0 1e-06 
0.0 0.7164 0 2.0 1e-06 
0.0 0.7165 0 2.0 1e-06 
0.0 0.7166 0 2.0 1e-06 
0.0 0.7167 0 2.0 1e-06 
0.0 0.7168 0 2.0 1e-06 
0.0 0.7169 0 2.0 1e-06 
0.0 0.717 0 2.0 1e-06 
0.0 0.7171 0 2.0 1e-06 
0.0 0.7172 0 2.0 1e-06 
0.0 0.7173 0 2.0 1e-06 
0.0 0.7174 0 2.0 1e-06 
0.0 0.7175 0 2.0 1e-06 
0.0 0.7176 0 2.0 1e-06 
0.0 0.7177 0 2.0 1e-06 
0.0 0.7178 0 2.0 1e-06 
0.0 0.7179 0 2.0 1e-06 
0.0 0.718 0 2.0 1e-06 
0.0 0.7181 0 2.0 1e-06 
0.0 0.7182 0 2.0 1e-06 
0.0 0.7183 0 2.0 1e-06 
0.0 0.7184 0 2.0 1e-06 
0.0 0.7185 0 2.0 1e-06 
0.0 0.7186 0 2.0 1e-06 
0.0 0.7187 0 2.0 1e-06 
0.0 0.7188 0 2.0 1e-06 
0.0 0.7189 0 2.0 1e-06 
0.0 0.719 0 2.0 1e-06 
0.0 0.7191 0 2.0 1e-06 
0.0 0.7192 0 2.0 1e-06 
0.0 0.7193 0 2.0 1e-06 
0.0 0.7194 0 2.0 1e-06 
0.0 0.7195 0 2.0 1e-06 
0.0 0.7196 0 2.0 1e-06 
0.0 0.7197 0 2.0 1e-06 
0.0 0.7198 0 2.0 1e-06 
0.0 0.7199 0 2.0 1e-06 
0.0 0.72 0 2.0 1e-06 
0.0 0.7201 0 2.0 1e-06 
0.0 0.7202 0 2.0 1e-06 
0.0 0.7203 0 2.0 1e-06 
0.0 0.7204 0 2.0 1e-06 
0.0 0.7205 0 2.0 1e-06 
0.0 0.7206 0 2.0 1e-06 
0.0 0.7207 0 2.0 1e-06 
0.0 0.7208 0 2.0 1e-06 
0.0 0.7209 0 2.0 1e-06 
0.0 0.721 0 2.0 1e-06 
0.0 0.7211 0 2.0 1e-06 
0.0 0.7212 0 2.0 1e-06 
0.0 0.7213 0 2.0 1e-06 
0.0 0.7214 0 2.0 1e-06 
0.0 0.7215 0 2.0 1e-06 
0.0 0.7216 0 2.0 1e-06 
0.0 0.7217 0 2.0 1e-06 
0.0 0.7218 0 2.0 1e-06 
0.0 0.7219 0 2.0 1e-06 
0.0 0.722 0 2.0 1e-06 
0.0 0.7221 0 2.0 1e-06 
0.0 0.7222 0 2.0 1e-06 
0.0 0.7223 0 2.0 1e-06 
0.0 0.7224 0 2.0 1e-06 
0.0 0.7225 0 2.0 1e-06 
0.0 0.7226 0 2.0 1e-06 
0.0 0.7227 0 2.0 1e-06 
0.0 0.7228 0 2.0 1e-06 
0.0 0.7229 0 2.0 1e-06 
0.0 0.723 0 2.0 1e-06 
0.0 0.7231 0 2.0 1e-06 
0.0 0.7232 0 2.0 1e-06 
0.0 0.7233 0 2.0 1e-06 
0.0 0.7234 0 2.0 1e-06 
0.0 0.7235 0 2.0 1e-06 
0.0 0.7236 0 2.0 1e-06 
0.0 0.7237 0 2.0 1e-06 
0.0 0.7238 0 2.0 1e-06 
0.0 0.7239 0 2.0 1e-06 
0.0 0.724 0 2.0 1e-06 
0.0 0.7241 0 2.0 1e-06 
0.0 0.7242 0 2.0 1e-06 
0.0 0.7243 0 2.0 1e-06 
0.0 0.7244 0 2.0 1e-06 
0.0 0.7245 0 2.0 1e-06 
0.0 0.7246 0 2.0 1e-06 
0.0 0.7247 0 2.0 1e-06 
0.0 0.7248 0 2.0 1e-06 
0.0 0.7249 0 2.0 1e-06 
0.0 0.725 0 2.0 1e-06 
0.0 0.7251 0 2.0 1e-06 
0.0 0.7252 0 2.0 1e-06 
0.0 0.7253 0 2.0 1e-06 
0.0 0.7254 0 2.0 1e-06 
0.0 0.7255 0 2.0 1e-06 
0.0 0.7256 0 2.0 1e-06 
0.0 0.7257 0 2.0 1e-06 
0.0 0.7258 0 2.0 1e-06 
0.0 0.7259 0 2.0 1e-06 
0.0 0.726 0 2.0 1e-06 
0.0 0.7261 0 2.0 1e-06 
0.0 0.7262 0 2.0 1e-06 
0.0 0.7263 0 2.0 1e-06 
0.0 0.7264 0 2.0 1e-06 
0.0 0.7265 0 2.0 1e-06 
0.0 0.7266 0 2.0 1e-06 
0.0 0.7267 0 2.0 1e-06 
0.0 0.7268 0 2.0 1e-06 
0.0 0.7269 0 2.0 1e-06 
0.0 0.727 0 2.0 1e-06 
0.0 0.7271 0 2.0 1e-06 
0.0 0.7272 0 2.0 1e-06 
0.0 0.7273 0 2.0 1e-06 
0.0 0.7274 0 2.0 1e-06 
0.0 0.7275 0 2.0 1e-06 
0.0 0.7276 0 2.0 1e-06 
0.0 0.7277 0 2.0 1e-06 
0.0 0.7278 0 2.0 1e-06 
0.0 0.7279 0 2.0 1e-06 
0.0 0.728 0 2.0 1e-06 
0.0 0.7281 0 2.0 1e-06 
0.0 0.7282 0 2.0 1e-06 
0.0 0.7283 0 2.0 1e-06 
0.0 0.7284 0 2.0 1e-06 
0.0 0.7285 0 2.0 1e-06 
0.0 0.7286 0 2.0 1e-06 
0.0 0.7287 0 2.0 1e-06 
0.0 0.7288 0 2.0 1e-06 
0.0 0.7289 0 2.0 1e-06 
0.0 0.729 0 2.0 1e-06 
0.0 0.7291 0 2.0 1e-06 
0.0 0.7292 0 2.0 1e-06 
0.0 0.7293 0 2.0 1e-06 
0.0 0.7294 0 2.0 1e-06 
0.0 0.7295 0 2.0 1e-06 
0.0 0.7296 0 2.0 1e-06 
0.0 0.7297 0 2.0 1e-06 
0.0 0.7298 0 2.0 1e-06 
0.0 0.7299 0 2.0 1e-06 
0.0 0.73 0 2.0 1e-06 
0.0 0.7301 0 2.0 1e-06 
0.0 0.7302 0 2.0 1e-06 
0.0 0.7303 0 2.0 1e-06 
0.0 0.7304 0 2.0 1e-06 
0.0 0.7305 0 2.0 1e-06 
0.0 0.7306 0 2.0 1e-06 
0.0 0.7307 0 2.0 1e-06 
0.0 0.7308 0 2.0 1e-06 
0.0 0.7309 0 2.0 1e-06 
0.0 0.731 0 2.0 1e-06 
0.0 0.7311 0 2.0 1e-06 
0.0 0.7312 0 2.0 1e-06 
0.0 0.7313 0 2.0 1e-06 
0.0 0.7314 0 2.0 1e-06 
0.0 0.7315 0 2.0 1e-06 
0.0 0.7316 0 2.0 1e-06 
0.0 0.7317 0 2.0 1e-06 
0.0 0.7318 0 2.0 1e-06 
0.0 0.7319 0 2.0 1e-06 
0.0 0.732 0 2.0 1e-06 
0.0 0.7321 0 2.0 1e-06 
0.0 0.7322 0 2.0 1e-06 
0.0 0.7323 0 2.0 1e-06 
0.0 0.7324 0 2.0 1e-06 
0.0 0.7325 0 2.0 1e-06 
0.0 0.7326 0 2.0 1e-06 
0.0 0.7327 0 2.0 1e-06 
0.0 0.7328 0 2.0 1e-06 
0.0 0.7329 0 2.0 1e-06 
0.0 0.733 0 2.0 1e-06 
0.0 0.7331 0 2.0 1e-06 
0.0 0.7332 0 2.0 1e-06 
0.0 0.7333 0 2.0 1e-06 
0.0 0.7334 0 2.0 1e-06 
0.0 0.7335 0 2.0 1e-06 
0.0 0.7336 0 2.0 1e-06 
0.0 0.7337 0 2.0 1e-06 
0.0 0.7338 0 2.0 1e-06 
0.0 0.7339 0 2.0 1e-06 
0.0 0.734 0 2.0 1e-06 
0.0 0.7341 0 2.0 1e-06 
0.0 0.7342 0 2.0 1e-06 
0.0 0.7343 0 2.0 1e-06 
0.0 0.7344 0 2.0 1e-06 
0.0 0.7345 0 2.0 1e-06 
0.0 0.7346 0 2.0 1e-06 
0.0 0.7347 0 2.0 1e-06 
0.0 0.7348 0 2.0 1e-06 
0.0 0.7349 0 2.0 1e-06 
0.0 0.735 0 2.0 1e-06 
0.0 0.7351 0 2.0 1e-06 
0.0 0.7352 0 2.0 1e-06 
0.0 0.7353 0 2.0 1e-06 
0.0 0.7354 0 2.0 1e-06 
0.0 0.7355 0 2.0 1e-06 
0.0 0.7356 0 2.0 1e-06 
0.0 0.7357 0 2.0 1e-06 
0.0 0.7358 0 2.0 1e-06 
0.0 0.7359 0 2.0 1e-06 
0.0 0.736 0 2.0 1e-06 
0.0 0.7361 0 2.0 1e-06 
0.0 0.7362 0 2.0 1e-06 
0.0 0.7363 0 2.0 1e-06 
0.0 0.7364 0 2.0 1e-06 
0.0 0.7365 0 2.0 1e-06 
0.0 0.7366 0 2.0 1e-06 
0.0 0.7367 0 2.0 1e-06 
0.0 0.7368 0 2.0 1e-06 
0.0 0.7369 0 2.0 1e-06 
0.0 0.737 0 2.0 1e-06 
0.0 0.7371 0 2.0 1e-06 
0.0 0.7372 0 2.0 1e-06 
0.0 0.7373 0 2.0 1e-06 
0.0 0.7374 0 2.0 1e-06 
0.0 0.7375 0 2.0 1e-06 
0.0 0.7376 0 2.0 1e-06 
0.0 0.7377 0 2.0 1e-06 
0.0 0.7378 0 2.0 1e-06 
0.0 0.7379 0 2.0 1e-06 
0.0 0.738 0 2.0 1e-06 
0.0 0.7381 0 2.0 1e-06 
0.0 0.7382 0 2.0 1e-06 
0.0 0.7383 0 2.0 1e-06 
0.0 0.7384 0 2.0 1e-06 
0.0 0.7385 0 2.0 1e-06 
0.0 0.7386 0 2.0 1e-06 
0.0 0.7387 0 2.0 1e-06 
0.0 0.7388 0 2.0 1e-06 
0.0 0.7389 0 2.0 1e-06 
0.0 0.739 0 2.0 1e-06 
0.0 0.7391 0 2.0 1e-06 
0.0 0.7392 0 2.0 1e-06 
0.0 0.7393 0 2.0 1e-06 
0.0 0.7394 0 2.0 1e-06 
0.0 0.7395 0 2.0 1e-06 
0.0 0.7396 0 2.0 1e-06 
0.0 0.7397 0 2.0 1e-06 
0.0 0.7398 0 2.0 1e-06 
0.0 0.7399 0 2.0 1e-06 
0.0 0.74 0 2.0 1e-06 
0.0 0.7401 0 2.0 1e-06 
0.0 0.7402 0 2.0 1e-06 
0.0 0.7403 0 2.0 1e-06 
0.0 0.7404 0 2.0 1e-06 
0.0 0.7405 0 2.0 1e-06 
0.0 0.7406 0 2.0 1e-06 
0.0 0.7407 0 2.0 1e-06 
0.0 0.7408 0 2.0 1e-06 
0.0 0.7409 0 2.0 1e-06 
0.0 0.741 0 2.0 1e-06 
0.0 0.7411 0 2.0 1e-06 
0.0 0.7412 0 2.0 1e-06 
0.0 0.7413 0 2.0 1e-06 
0.0 0.7414 0 2.0 1e-06 
0.0 0.7415 0 2.0 1e-06 
0.0 0.7416 0 2.0 1e-06 
0.0 0.7417 0 2.0 1e-06 
0.0 0.7418 0 2.0 1e-06 
0.0 0.7419 0 2.0 1e-06 
0.0 0.742 0 2.0 1e-06 
0.0 0.7421 0 2.0 1e-06 
0.0 0.7422 0 2.0 1e-06 
0.0 0.7423 0 2.0 1e-06 
0.0 0.7424 0 2.0 1e-06 
0.0 0.7425 0 2.0 1e-06 
0.0 0.7426 0 2.0 1e-06 
0.0 0.7427 0 2.0 1e-06 
0.0 0.7428 0 2.0 1e-06 
0.0 0.7429 0 2.0 1e-06 
0.0 0.743 0 2.0 1e-06 
0.0 0.7431 0 2.0 1e-06 
0.0 0.7432 0 2.0 1e-06 
0.0 0.7433 0 2.0 1e-06 
0.0 0.7434 0 2.0 1e-06 
0.0 0.7435 0 2.0 1e-06 
0.0 0.7436 0 2.0 1e-06 
0.0 0.7437 0 2.0 1e-06 
0.0 0.7438 0 2.0 1e-06 
0.0 0.7439 0 2.0 1e-06 
0.0 0.744 0 2.0 1e-06 
0.0 0.7441 0 2.0 1e-06 
0.0 0.7442 0 2.0 1e-06 
0.0 0.7443 0 2.0 1e-06 
0.0 0.7444 0 2.0 1e-06 
0.0 0.7445 0 2.0 1e-06 
0.0 0.7446 0 2.0 1e-06 
0.0 0.7447 0 2.0 1e-06 
0.0 0.7448 0 2.0 1e-06 
0.0 0.7449 0 2.0 1e-06 
0.0 0.745 0 2.0 1e-06 
0.0 0.7451 0 2.0 1e-06 
0.0 0.7452 0 2.0 1e-06 
0.0 0.7453 0 2.0 1e-06 
0.0 0.7454 0 2.0 1e-06 
0.0 0.7455 0 2.0 1e-06 
0.0 0.7456 0 2.0 1e-06 
0.0 0.7457 0 2.0 1e-06 
0.0 0.7458 0 2.0 1e-06 
0.0 0.7459 0 2.0 1e-06 
0.0 0.746 0 2.0 1e-06 
0.0 0.7461 0 2.0 1e-06 
0.0 0.7462 0 2.0 1e-06 
0.0 0.7463 0 2.0 1e-06 
0.0 0.7464 0 2.0 1e-06 
0.0 0.7465 0 2.0 1e-06 
0.0 0.7466 0 2.0 1e-06 
0.0 0.7467 0 2.0 1e-06 
0.0 0.7468 0 2.0 1e-06 
0.0 0.7469 0 2.0 1e-06 
0.0 0.747 0 2.0 1e-06 
0.0 0.7471 0 2.0 1e-06 
0.0 0.7472 0 2.0 1e-06 
0.0 0.7473 0 2.0 1e-06 
0.0 0.7474 0 2.0 1e-06 
0.0 0.7475 0 2.0 1e-06 
0.0 0.7476 0 2.0 1e-06 
0.0 0.7477 0 2.0 1e-06 
0.0 0.7478 0 2.0 1e-06 
0.0 0.7479 0 2.0 1e-06 
0.0 0.748 0 2.0 1e-06 
0.0 0.7481 0 2.0 1e-06 
0.0 0.7482 0 2.0 1e-06 
0.0 0.7483 0 2.0 1e-06 
0.0 0.7484 0 2.0 1e-06 
0.0 0.7485 0 2.0 1e-06 
0.0 0.7486 0 2.0 1e-06 
0.0 0.7487 0 2.0 1e-06 
0.0 0.7488 0 2.0 1e-06 
0.0 0.7489 0 2.0 1e-06 
0.0 0.749 0 2.0 1e-06 
0.0 0.7491 0 2.0 1e-06 
0.0 0.7492 0 2.0 1e-06 
0.0 0.7493 0 2.0 1e-06 
0.0 0.7494 0 2.0 1e-06 
0.0 0.7495 0 2.0 1e-06 
0.0 0.7496 0 2.0 1e-06 
0.0 0.7497 0 2.0 1e-06 
0.0 0.7498 0 2.0 1e-06 
0.0 0.7499 0 2.0 1e-06 
0.0 0.75 0 2.0 1e-06 
0.0 0.7501 0 2.0 1e-06 
0.0 0.7502 0 2.0 1e-06 
0.0 0.7503 0 2.0 1e-06 
0.0 0.7504 0 2.0 1e-06 
0.0 0.7505 0 2.0 1e-06 
0.0 0.7506 0 2.0 1e-06 
0.0 0.7507 0 2.0 1e-06 
0.0 0.7508 0 2.0 1e-06 
0.0 0.7509 0 2.0 1e-06 
0.0 0.751 0 2.0 1e-06 
0.0 0.7511 0 2.0 1e-06 
0.0 0.7512 0 2.0 1e-06 
0.0 0.7513 0 2.0 1e-06 
0.0 0.7514 0 2.0 1e-06 
0.0 0.7515 0 2.0 1e-06 
0.0 0.7516 0 2.0 1e-06 
0.0 0.7517 0 2.0 1e-06 
0.0 0.7518 0 2.0 1e-06 
0.0 0.7519 0 2.0 1e-06 
0.0 0.752 0 2.0 1e-06 
0.0 0.7521 0 2.0 1e-06 
0.0 0.7522 0 2.0 1e-06 
0.0 0.7523 0 2.0 1e-06 
0.0 0.7524 0 2.0 1e-06 
0.0 0.7525 0 2.0 1e-06 
0.0 0.7526 0 2.0 1e-06 
0.0 0.7527 0 2.0 1e-06 
0.0 0.7528 0 2.0 1e-06 
0.0 0.7529 0 2.0 1e-06 
0.0 0.753 0 2.0 1e-06 
0.0 0.7531 0 2.0 1e-06 
0.0 0.7532 0 2.0 1e-06 
0.0 0.7533 0 2.0 1e-06 
0.0 0.7534 0 2.0 1e-06 
0.0 0.7535 0 2.0 1e-06 
0.0 0.7536 0 2.0 1e-06 
0.0 0.7537 0 2.0 1e-06 
0.0 0.7538 0 2.0 1e-06 
0.0 0.7539 0 2.0 1e-06 
0.0 0.754 0 2.0 1e-06 
0.0 0.7541 0 2.0 1e-06 
0.0 0.7542 0 2.0 1e-06 
0.0 0.7543 0 2.0 1e-06 
0.0 0.7544 0 2.0 1e-06 
0.0 0.7545 0 2.0 1e-06 
0.0 0.7546 0 2.0 1e-06 
0.0 0.7547 0 2.0 1e-06 
0.0 0.7548 0 2.0 1e-06 
0.0 0.7549 0 2.0 1e-06 
0.0 0.755 0 2.0 1e-06 
0.0 0.7551 0 2.0 1e-06 
0.0 0.7552 0 2.0 1e-06 
0.0 0.7553 0 2.0 1e-06 
0.0 0.7554 0 2.0 1e-06 
0.0 0.7555 0 2.0 1e-06 
0.0 0.7556 0 2.0 1e-06 
0.0 0.7557 0 2.0 1e-06 
0.0 0.7558 0 2.0 1e-06 
0.0 0.7559 0 2.0 1e-06 
0.0 0.756 0 2.0 1e-06 
0.0 0.7561 0 2.0 1e-06 
0.0 0.7562 0 2.0 1e-06 
0.0 0.7563 0 2.0 1e-06 
0.0 0.7564 0 2.0 1e-06 
0.0 0.7565 0 2.0 1e-06 
0.0 0.7566 0 2.0 1e-06 
0.0 0.7567 0 2.0 1e-06 
0.0 0.7568 0 2.0 1e-06 
0.0 0.7569 0 2.0 1e-06 
0.0 0.757 0 2.0 1e-06 
0.0 0.7571 0 2.0 1e-06 
0.0 0.7572 0 2.0 1e-06 
0.0 0.7573 0 2.0 1e-06 
0.0 0.7574 0 2.0 1e-06 
0.0 0.7575 0 2.0 1e-06 
0.0 0.7576 0 2.0 1e-06 
0.0 0.7577 0 2.0 1e-06 
0.0 0.7578 0 2.0 1e-06 
0.0 0.7579 0 2.0 1e-06 
0.0 0.758 0 2.0 1e-06 
0.0 0.7581 0 2.0 1e-06 
0.0 0.7582 0 2.0 1e-06 
0.0 0.7583 0 2.0 1e-06 
0.0 0.7584 0 2.0 1e-06 
0.0 0.7585 0 2.0 1e-06 
0.0 0.7586 0 2.0 1e-06 
0.0 0.7587 0 2.0 1e-06 
0.0 0.7588 0 2.0 1e-06 
0.0 0.7589 0 2.0 1e-06 
0.0 0.759 0 2.0 1e-06 
0.0 0.7591 0 2.0 1e-06 
0.0 0.7592 0 2.0 1e-06 
0.0 0.7593 0 2.0 1e-06 
0.0 0.7594 0 2.0 1e-06 
0.0 0.7595 0 2.0 1e-06 
0.0 0.7596 0 2.0 1e-06 
0.0 0.7597 0 2.0 1e-06 
0.0 0.7598 0 2.0 1e-06 
0.0 0.7599 0 2.0 1e-06 
0.0 0.76 0 2.0 1e-06 
0.0 0.7601 0 2.0 1e-06 
0.0 0.7602 0 2.0 1e-06 
0.0 0.7603 0 2.0 1e-06 
0.0 0.7604 0 2.0 1e-06 
0.0 0.7605 0 2.0 1e-06 
0.0 0.7606 0 2.0 1e-06 
0.0 0.7607 0 2.0 1e-06 
0.0 0.7608 0 2.0 1e-06 
0.0 0.7609 0 2.0 1e-06 
0.0 0.761 0 2.0 1e-06 
0.0 0.7611 0 2.0 1e-06 
0.0 0.7612 0 2.0 1e-06 
0.0 0.7613 0 2.0 1e-06 
0.0 0.7614 0 2.0 1e-06 
0.0 0.7615 0 2.0 1e-06 
0.0 0.7616 0 2.0 1e-06 
0.0 0.7617 0 2.0 1e-06 
0.0 0.7618 0 2.0 1e-06 
0.0 0.7619 0 2.0 1e-06 
0.0 0.762 0 2.0 1e-06 
0.0 0.7621 0 2.0 1e-06 
0.0 0.7622 0 2.0 1e-06 
0.0 0.7623 0 2.0 1e-06 
0.0 0.7624 0 2.0 1e-06 
0.0 0.7625 0 2.0 1e-06 
0.0 0.7626 0 2.0 1e-06 
0.0 0.7627 0 2.0 1e-06 
0.0 0.7628 0 2.0 1e-06 
0.0 0.7629 0 2.0 1e-06 
0.0 0.763 0 2.0 1e-06 
0.0 0.7631 0 2.0 1e-06 
0.0 0.7632 0 2.0 1e-06 
0.0 0.7633 0 2.0 1e-06 
0.0 0.7634 0 2.0 1e-06 
0.0 0.7635 0 2.0 1e-06 
0.0 0.7636 0 2.0 1e-06 
0.0 0.7637 0 2.0 1e-06 
0.0 0.7638 0 2.0 1e-06 
0.0 0.7639 0 2.0 1e-06 
0.0 0.764 0 2.0 1e-06 
0.0 0.7641 0 2.0 1e-06 
0.0 0.7642 0 2.0 1e-06 
0.0 0.7643 0 2.0 1e-06 
0.0 0.7644 0 2.0 1e-06 
0.0 0.7645 0 2.0 1e-06 
0.0 0.7646 0 2.0 1e-06 
0.0 0.7647 0 2.0 1e-06 
0.0 0.7648 0 2.0 1e-06 
0.0 0.7649 0 2.0 1e-06 
0.0 0.765 0 2.0 1e-06 
0.0 0.7651 0 2.0 1e-06 
0.0 0.7652 0 2.0 1e-06 
0.0 0.7653 0 2.0 1e-06 
0.0 0.7654 0 2.0 1e-06 
0.0 0.7655 0 2.0 1e-06 
0.0 0.7656 0 2.0 1e-06 
0.0 0.7657 0 2.0 1e-06 
0.0 0.7658 0 2.0 1e-06 
0.0 0.7659 0 2.0 1e-06 
0.0 0.766 0 2.0 1e-06 
0.0 0.7661 0 2.0 1e-06 
0.0 0.7662 0 2.0 1e-06 
0.0 0.7663 0 2.0 1e-06 
0.0 0.7664 0 2.0 1e-06 
0.0 0.7665 0 2.0 1e-06 
0.0 0.7666 0 2.0 1e-06 
0.0 0.7667 0 2.0 1e-06 
0.0 0.7668 0 2.0 1e-06 
0.0 0.7669 0 2.0 1e-06 
0.0 0.767 0 2.0 1e-06 
0.0 0.7671 0 2.0 1e-06 
0.0 0.7672 0 2.0 1e-06 
0.0 0.7673 0 2.0 1e-06 
0.0 0.7674 0 2.0 1e-06 
0.0 0.7675 0 2.0 1e-06 
0.0 0.7676 0 2.0 1e-06 
0.0 0.7677 0 2.0 1e-06 
0.0 0.7678 0 2.0 1e-06 
0.0 0.7679 0 2.0 1e-06 
0.0 0.768 0 2.0 1e-06 
0.0 0.7681 0 2.0 1e-06 
0.0 0.7682 0 2.0 1e-06 
0.0 0.7683 0 2.0 1e-06 
0.0 0.7684 0 2.0 1e-06 
0.0 0.7685 0 2.0 1e-06 
0.0 0.7686 0 2.0 1e-06 
0.0 0.7687 0 2.0 1e-06 
0.0 0.7688 0 2.0 1e-06 
0.0 0.7689 0 2.0 1e-06 
0.0 0.769 0 2.0 1e-06 
0.0 0.7691 0 2.0 1e-06 
0.0 0.7692 0 2.0 1e-06 
0.0 0.7693 0 2.0 1e-06 
0.0 0.7694 0 2.0 1e-06 
0.0 0.7695 0 2.0 1e-06 
0.0 0.7696 0 2.0 1e-06 
0.0 0.7697 0 2.0 1e-06 
0.0 0.7698 0 2.0 1e-06 
0.0 0.7699 0 2.0 1e-06 
0.0 0.77 0 2.0 1e-06 
0.0 0.7701 0 2.0 1e-06 
0.0 0.7702 0 2.0 1e-06 
0.0 0.7703 0 2.0 1e-06 
0.0 0.7704 0 2.0 1e-06 
0.0 0.7705 0 2.0 1e-06 
0.0 0.7706 0 2.0 1e-06 
0.0 0.7707 0 2.0 1e-06 
0.0 0.7708 0 2.0 1e-06 
0.0 0.7709 0 2.0 1e-06 
0.0 0.771 0 2.0 1e-06 
0.0 0.7711 0 2.0 1e-06 
0.0 0.7712 0 2.0 1e-06 
0.0 0.7713 0 2.0 1e-06 
0.0 0.7714 0 2.0 1e-06 
0.0 0.7715 0 2.0 1e-06 
0.0 0.7716 0 2.0 1e-06 
0.0 0.7717 0 2.0 1e-06 
0.0 0.7718 0 2.0 1e-06 
0.0 0.7719 0 2.0 1e-06 
0.0 0.772 0 2.0 1e-06 
0.0 0.7721 0 2.0 1e-06 
0.0 0.7722 0 2.0 1e-06 
0.0 0.7723 0 2.0 1e-06 
0.0 0.7724 0 2.0 1e-06 
0.0 0.7725 0 2.0 1e-06 
0.0 0.7726 0 2.0 1e-06 
0.0 0.7727 0 2.0 1e-06 
0.0 0.7728 0 2.0 1e-06 
0.0 0.7729 0 2.0 1e-06 
0.0 0.773 0 2.0 1e-06 
0.0 0.7731 0 2.0 1e-06 
0.0 0.7732 0 2.0 1e-06 
0.0 0.7733 0 2.0 1e-06 
0.0 0.7734 0 2.0 1e-06 
0.0 0.7735 0 2.0 1e-06 
0.0 0.7736 0 2.0 1e-06 
0.0 0.7737 0 2.0 1e-06 
0.0 0.7738 0 2.0 1e-06 
0.0 0.7739 0 2.0 1e-06 
0.0 0.774 0 2.0 1e-06 
0.0 0.7741 0 2.0 1e-06 
0.0 0.7742 0 2.0 1e-06 
0.0 0.7743 0 2.0 1e-06 
0.0 0.7744 0 2.0 1e-06 
0.0 0.7745 0 2.0 1e-06 
0.0 0.7746 0 2.0 1e-06 
0.0 0.7747 0 2.0 1e-06 
0.0 0.7748 0 2.0 1e-06 
0.0 0.7749 0 2.0 1e-06 
0.0 0.775 0 2.0 1e-06 
0.0 0.7751 0 2.0 1e-06 
0.0 0.7752 0 2.0 1e-06 
0.0 0.7753 0 2.0 1e-06 
0.0 0.7754 0 2.0 1e-06 
0.0 0.7755 0 2.0 1e-06 
0.0 0.7756 0 2.0 1e-06 
0.0 0.7757 0 2.0 1e-06 
0.0 0.7758 0 2.0 1e-06 
0.0 0.7759 0 2.0 1e-06 
0.0 0.776 0 2.0 1e-06 
0.0 0.7761 0 2.0 1e-06 
0.0 0.7762 0 2.0 1e-06 
0.0 0.7763 0 2.0 1e-06 
0.0 0.7764 0 2.0 1e-06 
0.0 0.7765 0 2.0 1e-06 
0.0 0.7766 0 2.0 1e-06 
0.0 0.7767 0 2.0 1e-06 
0.0 0.7768 0 2.0 1e-06 
0.0 0.7769 0 2.0 1e-06 
0.0 0.777 0 2.0 1e-06 
0.0 0.7771 0 2.0 1e-06 
0.0 0.7772 0 2.0 1e-06 
0.0 0.7773 0 2.0 1e-06 
0.0 0.7774 0 2.0 1e-06 
0.0 0.7775 0 2.0 1e-06 
0.0 0.7776 0 2.0 1e-06 
0.0 0.7777 0 2.0 1e-06 
0.0 0.7778 0 2.0 1e-06 
0.0 0.7779 0 2.0 1e-06 
0.0 0.778 0 2.0 1e-06 
0.0 0.7781 0 2.0 1e-06 
0.0 0.7782 0 2.0 1e-06 
0.0 0.7783 0 2.0 1e-06 
0.0 0.7784 0 2.0 1e-06 
0.0 0.7785 0 2.0 1e-06 
0.0 0.7786 0 2.0 1e-06 
0.0 0.7787 0 2.0 1e-06 
0.0 0.7788 0 2.0 1e-06 
0.0 0.7789 0 2.0 1e-06 
0.0 0.779 0 2.0 1e-06 
0.0 0.7791 0 2.0 1e-06 
0.0 0.7792 0 2.0 1e-06 
0.0 0.7793 0 2.0 1e-06 
0.0 0.7794 0 2.0 1e-06 
0.0 0.7795 0 2.0 1e-06 
0.0 0.7796 0 2.0 1e-06 
0.0 0.7797 0 2.0 1e-06 
0.0 0.7798 0 2.0 1e-06 
0.0 0.7799 0 2.0 1e-06 
0.0 0.78 0 2.0 1e-06 
0.0 0.7801 0 2.0 1e-06 
0.0 0.7802 0 2.0 1e-06 
0.0 0.7803 0 2.0 1e-06 
0.0 0.7804 0 2.0 1e-06 
0.0 0.7805 0 2.0 1e-06 
0.0 0.7806 0 2.0 1e-06 
0.0 0.7807 0 2.0 1e-06 
0.0 0.7808 0 2.0 1e-06 
0.0 0.7809 0 2.0 1e-06 
0.0 0.781 0 2.0 1e-06 
0.0 0.7811 0 2.0 1e-06 
0.0 0.7812 0 2.0 1e-06 
0.0 0.7813 0 2.0 1e-06 
0.0 0.7814 0 2.0 1e-06 
0.0 0.7815 0 2.0 1e-06 
0.0 0.7816 0 2.0 1e-06 
0.0 0.7817 0 2.0 1e-06 
0.0 0.7818 0 2.0 1e-06 
0.0 0.7819 0 2.0 1e-06 
0.0 0.782 0 2.0 1e-06 
0.0 0.7821 0 2.0 1e-06 
0.0 0.7822 0 2.0 1e-06 
0.0 0.7823 0 2.0 1e-06 
0.0 0.7824 0 2.0 1e-06 
0.0 0.7825 0 2.0 1e-06 
0.0 0.7826 0 2.0 1e-06 
0.0 0.7827 0 2.0 1e-06 
0.0 0.7828 0 2.0 1e-06 
0.0 0.7829 0 2.0 1e-06 
0.0 0.783 0 2.0 1e-06 
0.0 0.7831 0 2.0 1e-06 
0.0 0.7832 0 2.0 1e-06 
0.0 0.7833 0 2.0 1e-06 
0.0 0.7834 0 2.0 1e-06 
0.0 0.7835 0 2.0 1e-06 
0.0 0.7836 0 2.0 1e-06 
0.0 0.7837 0 2.0 1e-06 
0.0 0.7838 0 2.0 1e-06 
0.0 0.7839 0 2.0 1e-06 
0.0 0.784 0 2.0 1e-06 
0.0 0.7841 0 2.0 1e-06 
0.0 0.7842 0 2.0 1e-06 
0.0 0.7843 0 2.0 1e-06 
0.0 0.7844 0 2.0 1e-06 
0.0 0.7845 0 2.0 1e-06 
0.0 0.7846 0 2.0 1e-06 
0.0 0.7847 0 2.0 1e-06 
0.0 0.7848 0 2.0 1e-06 
0.0 0.7849 0 2.0 1e-06 
0.0 0.785 0 2.0 1e-06 
0.0 0.7851 0 2.0 1e-06 
0.0 0.7852 0 2.0 1e-06 
0.0 0.7853 0 2.0 1e-06 
0.0 0.7854 0 2.0 1e-06 
0.0 0.7855 0 2.0 1e-06 
0.0 0.7856 0 2.0 1e-06 
0.0 0.7857 0 2.0 1e-06 
0.0 0.7858 0 2.0 1e-06 
0.0 0.7859 0 2.0 1e-06 
0.0 0.786 0 2.0 1e-06 
0.0 0.7861 0 2.0 1e-06 
0.0 0.7862 0 2.0 1e-06 
0.0 0.7863 0 2.0 1e-06 
0.0 0.7864 0 2.0 1e-06 
0.0 0.7865 0 2.0 1e-06 
0.0 0.7866 0 2.0 1e-06 
0.0 0.7867 0 2.0 1e-06 
0.0 0.7868 0 2.0 1e-06 
0.0 0.7869 0 2.0 1e-06 
0.0 0.787 0 2.0 1e-06 
0.0 0.7871 0 2.0 1e-06 
0.0 0.7872 0 2.0 1e-06 
0.0 0.7873 0 2.0 1e-06 
0.0 0.7874 0 2.0 1e-06 
0.0 0.7875 0 2.0 1e-06 
0.0 0.7876 0 2.0 1e-06 
0.0 0.7877 0 2.0 1e-06 
0.0 0.7878 0 2.0 1e-06 
0.0 0.7879 0 2.0 1e-06 
0.0 0.788 0 2.0 1e-06 
0.0 0.7881 0 2.0 1e-06 
0.0 0.7882 0 2.0 1e-06 
0.0 0.7883 0 2.0 1e-06 
0.0 0.7884 0 2.0 1e-06 
0.0 0.7885 0 2.0 1e-06 
0.0 0.7886 0 2.0 1e-06 
0.0 0.7887 0 2.0 1e-06 
0.0 0.7888 0 2.0 1e-06 
0.0 0.7889 0 2.0 1e-06 
0.0 0.789 0 2.0 1e-06 
0.0 0.7891 0 2.0 1e-06 
0.0 0.7892 0 2.0 1e-06 
0.0 0.7893 0 2.0 1e-06 
0.0 0.7894 0 2.0 1e-06 
0.0 0.7895 0 2.0 1e-06 
0.0 0.7896 0 2.0 1e-06 
0.0 0.7897 0 2.0 1e-06 
0.0 0.7898 0 2.0 1e-06 
0.0 0.7899 0 2.0 1e-06 
0.0 0.79 0 2.0 1e-06 
0.0 0.7901 0 2.0 1e-06 
0.0 0.7902 0 2.0 1e-06 
0.0 0.7903 0 2.0 1e-06 
0.0 0.7904 0 2.0 1e-06 
0.0 0.7905 0 2.0 1e-06 
0.0 0.7906 0 2.0 1e-06 
0.0 0.7907 0 2.0 1e-06 
0.0 0.7908 0 2.0 1e-06 
0.0 0.7909 0 2.0 1e-06 
0.0 0.791 0 2.0 1e-06 
0.0 0.7911 0 2.0 1e-06 
0.0 0.7912 0 2.0 1e-06 
0.0 0.7913 0 2.0 1e-06 
0.0 0.7914 0 2.0 1e-06 
0.0 0.7915 0 2.0 1e-06 
0.0 0.7916 0 2.0 1e-06 
0.0 0.7917 0 2.0 1e-06 
0.0 0.7918 0 2.0 1e-06 
0.0 0.7919 0 2.0 1e-06 
0.0 0.792 0 2.0 1e-06 
0.0 0.7921 0 2.0 1e-06 
0.0 0.7922 0 2.0 1e-06 
0.0 0.7923 0 2.0 1e-06 
0.0 0.7924 0 2.0 1e-06 
0.0 0.7925 0 2.0 1e-06 
0.0 0.7926 0 2.0 1e-06 
0.0 0.7927 0 2.0 1e-06 
0.0 0.7928 0 2.0 1e-06 
0.0 0.7929 0 2.0 1e-06 
0.0 0.793 0 2.0 1e-06 
0.0 0.7931 0 2.0 1e-06 
0.0 0.7932 0 2.0 1e-06 
0.0 0.7933 0 2.0 1e-06 
0.0 0.7934 0 2.0 1e-06 
0.0 0.7935 0 2.0 1e-06 
0.0 0.7936 0 2.0 1e-06 
0.0 0.7937 0 2.0 1e-06 
0.0 0.7938 0 2.0 1e-06 
0.0 0.7939 0 2.0 1e-06 
0.0 0.794 0 2.0 1e-06 
0.0 0.7941 0 2.0 1e-06 
0.0 0.7942 0 2.0 1e-06 
0.0 0.7943 0 2.0 1e-06 
0.0 0.7944 0 2.0 1e-06 
0.0 0.7945 0 2.0 1e-06 
0.0 0.7946 0 2.0 1e-06 
0.0 0.7947 0 2.0 1e-06 
0.0 0.7948 0 2.0 1e-06 
0.0 0.7949 0 2.0 1e-06 
0.0 0.795 0 2.0 1e-06 
0.0 0.7951 0 2.0 1e-06 
0.0 0.7952 0 2.0 1e-06 
0.0 0.7953 0 2.0 1e-06 
0.0 0.7954 0 2.0 1e-06 
0.0 0.7955 0 2.0 1e-06 
0.0 0.7956 0 2.0 1e-06 
0.0 0.7957 0 2.0 1e-06 
0.0 0.7958 0 2.0 1e-06 
0.0 0.7959 0 2.0 1e-06 
0.0 0.796 0 2.0 1e-06 
0.0 0.7961 0 2.0 1e-06 
0.0 0.7962 0 2.0 1e-06 
0.0 0.7963 0 2.0 1e-06 
0.0 0.7964 0 2.0 1e-06 
0.0 0.7965 0 2.0 1e-06 
0.0 0.7966 0 2.0 1e-06 
0.0 0.7967 0 2.0 1e-06 
0.0 0.7968 0 2.0 1e-06 
0.0 0.7969 0 2.0 1e-06 
0.0 0.797 0 2.0 1e-06 
0.0 0.7971 0 2.0 1e-06 
0.0 0.7972 0 2.0 1e-06 
0.0 0.7973 0 2.0 1e-06 
0.0 0.7974 0 2.0 1e-06 
0.0 0.7975 0 2.0 1e-06 
0.0 0.7976 0 2.0 1e-06 
0.0 0.7977 0 2.0 1e-06 
0.0 0.7978 0 2.0 1e-06 
0.0 0.7979 0 2.0 1e-06 
0.0 0.798 0 2.0 1e-06 
0.0 0.7981 0 2.0 1e-06 
0.0 0.7982 0 2.0 1e-06 
0.0 0.7983 0 2.0 1e-06 
0.0 0.7984 0 2.0 1e-06 
0.0 0.7985 0 2.0 1e-06 
0.0 0.7986 0 2.0 1e-06 
0.0 0.7987 0 2.0 1e-06 
0.0 0.7988 0 2.0 1e-06 
0.0 0.7989 0 2.0 1e-06 
0.0 0.799 0 2.0 1e-06 
0.0 0.7991 0 2.0 1e-06 
0.0 0.7992 0 2.0 1e-06 
0.0 0.7993 0 2.0 1e-06 
0.0 0.7994 0 2.0 1e-06 
0.0 0.7995 0 2.0 1e-06 
0.0 0.7996 0 2.0 1e-06 
0.0 0.7997 0 2.0 1e-06 
0.0 0.7998 0 2.0 1e-06 
0.0 0.7999 0 2.0 1e-06 
0.0 0.8 0 2.0 1e-06 
0.0 0.8001 0 2.0 1e-06 
0.0 0.8002 0 2.0 1e-06 
0.0 0.8003 0 2.0 1e-06 
0.0 0.8004 0 2.0 1e-06 
0.0 0.8005 0 2.0 1e-06 
0.0 0.8006 0 2.0 1e-06 
0.0 0.8007 0 2.0 1e-06 
0.0 0.8008 0 2.0 1e-06 
0.0 0.8009 0 2.0 1e-06 
0.0 0.801 0 2.0 1e-06 
0.0 0.8011 0 2.0 1e-06 
0.0 0.8012 0 2.0 1e-06 
0.0 0.8013 0 2.0 1e-06 
0.0 0.8014 0 2.0 1e-06 
0.0 0.8015 0 2.0 1e-06 
0.0 0.8016 0 2.0 1e-06 
0.0 0.8017 0 2.0 1e-06 
0.0 0.8018 0 2.0 1e-06 
0.0 0.8019 0 2.0 1e-06 
0.0 0.802 0 2.0 1e-06 
0.0 0.8021 0 2.0 1e-06 
0.0 0.8022 0 2.0 1e-06 
0.0 0.8023 0 2.0 1e-06 
0.0 0.8024 0 2.0 1e-06 
0.0 0.8025 0 2.0 1e-06 
0.0 0.8026 0 2.0 1e-06 
0.0 0.8027 0 2.0 1e-06 
0.0 0.8028 0 2.0 1e-06 
0.0 0.8029 0 2.0 1e-06 
0.0 0.803 0 2.0 1e-06 
0.0 0.8031 0 2.0 1e-06 
0.0 0.8032 0 2.0 1e-06 
0.0 0.8033 0 2.0 1e-06 
0.0 0.8034 0 2.0 1e-06 
0.0 0.8035 0 2.0 1e-06 
0.0 0.8036 0 2.0 1e-06 
0.0 0.8037 0 2.0 1e-06 
0.0 0.8038 0 2.0 1e-06 
0.0 0.8039 0 2.0 1e-06 
0.0 0.804 0 2.0 1e-06 
0.0 0.8041 0 2.0 1e-06 
0.0 0.8042 0 2.0 1e-06 
0.0 0.8043 0 2.0 1e-06 
0.0 0.8044 0 2.0 1e-06 
0.0 0.8045 0 2.0 1e-06 
0.0 0.8046 0 2.0 1e-06 
0.0 0.8047 0 2.0 1e-06 
0.0 0.8048 0 2.0 1e-06 
0.0 0.8049 0 2.0 1e-06 
0.0 0.805 0 2.0 1e-06 
0.0 0.8051 0 2.0 1e-06 
0.0 0.8052 0 2.0 1e-06 
0.0 0.8053 0 2.0 1e-06 
0.0 0.8054 0 2.0 1e-06 
0.0 0.8055 0 2.0 1e-06 
0.0 0.8056 0 2.0 1e-06 
0.0 0.8057 0 2.0 1e-06 
0.0 0.8058 0 2.0 1e-06 
0.0 0.8059 0 2.0 1e-06 
0.0 0.806 0 2.0 1e-06 
0.0 0.8061 0 2.0 1e-06 
0.0 0.8062 0 2.0 1e-06 
0.0 0.8063 0 2.0 1e-06 
0.0 0.8064 0 2.0 1e-06 
0.0 0.8065 0 2.0 1e-06 
0.0 0.8066 0 2.0 1e-06 
0.0 0.8067 0 2.0 1e-06 
0.0 0.8068 0 2.0 1e-06 
0.0 0.8069 0 2.0 1e-06 
0.0 0.807 0 2.0 1e-06 
0.0 0.8071 0 2.0 1e-06 
0.0 0.8072 0 2.0 1e-06 
0.0 0.8073 0 2.0 1e-06 
0.0 0.8074 0 2.0 1e-06 
0.0 0.8075 0 2.0 1e-06 
0.0 0.8076 0 2.0 1e-06 
0.0 0.8077 0 2.0 1e-06 
0.0 0.8078 0 2.0 1e-06 
0.0 0.8079 0 2.0 1e-06 
0.0 0.808 0 2.0 1e-06 
0.0 0.8081 0 2.0 1e-06 
0.0 0.8082 0 2.0 1e-06 
0.0 0.8083 0 2.0 1e-06 
0.0 0.8084 0 2.0 1e-06 
0.0 0.8085 0 2.0 1e-06 
0.0 0.8086 0 2.0 1e-06 
0.0 0.8087 0 2.0 1e-06 
0.0 0.8088 0 2.0 1e-06 
0.0 0.8089 0 2.0 1e-06 
0.0 0.809 0 2.0 1e-06 
0.0 0.8091 0 2.0 1e-06 
0.0 0.8092 0 2.0 1e-06 
0.0 0.8093 0 2.0 1e-06 
0.0 0.8094 0 2.0 1e-06 
0.0 0.8095 0 2.0 1e-06 
0.0 0.8096 0 2.0 1e-06 
0.0 0.8097 0 2.0 1e-06 
0.0 0.8098 0 2.0 1e-06 
0.0 0.8099 0 2.0 1e-06 
0.0 0.81 0 2.0 1e-06 
0.0 0.8101 0 2.0 1e-06 
0.0 0.8102 0 2.0 1e-06 
0.0 0.8103 0 2.0 1e-06 
0.0 0.8104 0 2.0 1e-06 
0.0 0.8105 0 2.0 1e-06 
0.0 0.8106 0 2.0 1e-06 
0.0 0.8107 0 2.0 1e-06 
0.0 0.8108 0 2.0 1e-06 
0.0 0.8109 0 2.0 1e-06 
0.0 0.811 0 2.0 1e-06 
0.0 0.8111 0 2.0 1e-06 
0.0 0.8112 0 2.0 1e-06 
0.0 0.8113 0 2.0 1e-06 
0.0 0.8114 0 2.0 1e-06 
0.0 0.8115 0 2.0 1e-06 
0.0 0.8116 0 2.0 1e-06 
0.0 0.8117 0 2.0 1e-06 
0.0 0.8118 0 2.0 1e-06 
0.0 0.8119 0 2.0 1e-06 
0.0 0.812 0 2.0 1e-06 
0.0 0.8121 0 2.0 1e-06 
0.0 0.8122 0 2.0 1e-06 
0.0 0.8123 0 2.0 1e-06 
0.0 0.8124 0 2.0 1e-06 
0.0 0.8125 0 2.0 1e-06 
0.0 0.8126 0 2.0 1e-06 
0.0 0.8127 0 2.0 1e-06 
0.0 0.8128 0 2.0 1e-06 
0.0 0.8129 0 2.0 1e-06 
0.0 0.813 0 2.0 1e-06 
0.0 0.8131 0 2.0 1e-06 
0.0 0.8132 0 2.0 1e-06 
0.0 0.8133 0 2.0 1e-06 
0.0 0.8134 0 2.0 1e-06 
0.0 0.8135 0 2.0 1e-06 
0.0 0.8136 0 2.0 1e-06 
0.0 0.8137 0 2.0 1e-06 
0.0 0.8138 0 2.0 1e-06 
0.0 0.8139 0 2.0 1e-06 
0.0 0.814 0 2.0 1e-06 
0.0 0.8141 0 2.0 1e-06 
0.0 0.8142 0 2.0 1e-06 
0.0 0.8143 0 2.0 1e-06 
0.0 0.8144 0 2.0 1e-06 
0.0 0.8145 0 2.0 1e-06 
0.0 0.8146 0 2.0 1e-06 
0.0 0.8147 0 2.0 1e-06 
0.0 0.8148 0 2.0 1e-06 
0.0 0.8149 0 2.0 1e-06 
0.0 0.815 0 2.0 1e-06 
0.0 0.8151 0 2.0 1e-06 
0.0 0.8152 0 2.0 1e-06 
0.0 0.8153 0 2.0 1e-06 
0.0 0.8154 0 2.0 1e-06 
0.0 0.8155 0 2.0 1e-06 
0.0 0.8156 0 2.0 1e-06 
0.0 0.8157 0 2.0 1e-06 
0.0 0.8158 0 2.0 1e-06 
0.0 0.8159 0 2.0 1e-06 
0.0 0.816 0 2.0 1e-06 
0.0 0.8161 0 2.0 1e-06 
0.0 0.8162 0 2.0 1e-06 
0.0 0.8163 0 2.0 1e-06 
0.0 0.8164 0 2.0 1e-06 
0.0 0.8165 0 2.0 1e-06 
0.0 0.8166 0 2.0 1e-06 
0.0 0.8167 0 2.0 1e-06 
0.0 0.8168 0 2.0 1e-06 
0.0 0.8169 0 2.0 1e-06 
0.0 0.817 0 2.0 1e-06 
0.0 0.8171 0 2.0 1e-06 
0.0 0.8172 0 2.0 1e-06 
0.0 0.8173 0 2.0 1e-06 
0.0 0.8174 0 2.0 1e-06 
0.0 0.8175 0 2.0 1e-06 
0.0 0.8176 0 2.0 1e-06 
0.0 0.8177 0 2.0 1e-06 
0.0 0.8178 0 2.0 1e-06 
0.0 0.8179 0 2.0 1e-06 
0.0 0.818 0 2.0 1e-06 
0.0 0.8181 0 2.0 1e-06 
0.0 0.8182 0 2.0 1e-06 
0.0 0.8183 0 2.0 1e-06 
0.0 0.8184 0 2.0 1e-06 
0.0 0.8185 0 2.0 1e-06 
0.0 0.8186 0 2.0 1e-06 
0.0 0.8187 0 2.0 1e-06 
0.0 0.8188 0 2.0 1e-06 
0.0 0.8189 0 2.0 1e-06 
0.0 0.819 0 2.0 1e-06 
0.0 0.8191 0 2.0 1e-06 
0.0 0.8192 0 2.0 1e-06 
0.0 0.8193 0 2.0 1e-06 
0.0 0.8194 0 2.0 1e-06 
0.0 0.8195 0 2.0 1e-06 
0.0 0.8196 0 2.0 1e-06 
0.0 0.8197 0 2.0 1e-06 
0.0 0.8198 0 2.0 1e-06 
0.0 0.8199 0 2.0 1e-06 
0.0 0.82 0 2.0 1e-06 
0.0 0.8201 0 2.0 1e-06 
0.0 0.8202 0 2.0 1e-06 
0.0 0.8203 0 2.0 1e-06 
0.0 0.8204 0 2.0 1e-06 
0.0 0.8205 0 2.0 1e-06 
0.0 0.8206 0 2.0 1e-06 
0.0 0.8207 0 2.0 1e-06 
0.0 0.8208 0 2.0 1e-06 
0.0 0.8209 0 2.0 1e-06 
0.0 0.821 0 2.0 1e-06 
0.0 0.8211 0 2.0 1e-06 
0.0 0.8212 0 2.0 1e-06 
0.0 0.8213 0 2.0 1e-06 
0.0 0.8214 0 2.0 1e-06 
0.0 0.8215 0 2.0 1e-06 
0.0 0.8216 0 2.0 1e-06 
0.0 0.8217 0 2.0 1e-06 
0.0 0.8218 0 2.0 1e-06 
0.0 0.8219 0 2.0 1e-06 
0.0 0.822 0 2.0 1e-06 
0.0 0.8221 0 2.0 1e-06 
0.0 0.8222 0 2.0 1e-06 
0.0 0.8223 0 2.0 1e-06 
0.0 0.8224 0 2.0 1e-06 
0.0 0.8225 0 2.0 1e-06 
0.0 0.8226 0 2.0 1e-06 
0.0 0.8227 0 2.0 1e-06 
0.0 0.8228 0 2.0 1e-06 
0.0 0.8229 0 2.0 1e-06 
0.0 0.823 0 2.0 1e-06 
0.0 0.8231 0 2.0 1e-06 
0.0 0.8232 0 2.0 1e-06 
0.0 0.8233 0 2.0 1e-06 
0.0 0.8234 0 2.0 1e-06 
0.0 0.8235 0 2.0 1e-06 
0.0 0.8236 0 2.0 1e-06 
0.0 0.8237 0 2.0 1e-06 
0.0 0.8238 0 2.0 1e-06 
0.0 0.8239 0 2.0 1e-06 
0.0 0.824 0 2.0 1e-06 
0.0 0.8241 0 2.0 1e-06 
0.0 0.8242 0 2.0 1e-06 
0.0 0.8243 0 2.0 1e-06 
0.0 0.8244 0 2.0 1e-06 
0.0 0.8245 0 2.0 1e-06 
0.0 0.8246 0 2.0 1e-06 
0.0 0.8247 0 2.0 1e-06 
0.0 0.8248 0 2.0 1e-06 
0.0 0.8249 0 2.0 1e-06 
0.0 0.825 0 2.0 1e-06 
0.0 0.8251 0 2.0 1e-06 
0.0 0.8252 0 2.0 1e-06 
0.0 0.8253 0 2.0 1e-06 
0.0 0.8254 0 2.0 1e-06 
0.0 0.8255 0 2.0 1e-06 
0.0 0.8256 0 2.0 1e-06 
0.0 0.8257 0 2.0 1e-06 
0.0 0.8258 0 2.0 1e-06 
0.0 0.8259 0 2.0 1e-06 
0.0 0.826 0 2.0 1e-06 
0.0 0.8261 0 2.0 1e-06 
0.0 0.8262 0 2.0 1e-06 
0.0 0.8263 0 2.0 1e-06 
0.0 0.8264 0 2.0 1e-06 
0.0 0.8265 0 2.0 1e-06 
0.0 0.8266 0 2.0 1e-06 
0.0 0.8267 0 2.0 1e-06 
0.0 0.8268 0 2.0 1e-06 
0.0 0.8269 0 2.0 1e-06 
0.0 0.827 0 2.0 1e-06 
0.0 0.8271 0 2.0 1e-06 
0.0 0.8272 0 2.0 1e-06 
0.0 0.8273 0 2.0 1e-06 
0.0 0.8274 0 2.0 1e-06 
0.0 0.8275 0 2.0 1e-06 
0.0 0.8276 0 2.0 1e-06 
0.0 0.8277 0 2.0 1e-06 
0.0 0.8278 0 2.0 1e-06 
0.0 0.8279 0 2.0 1e-06 
0.0 0.828 0 2.0 1e-06 
0.0 0.8281 0 2.0 1e-06 
0.0 0.8282 0 2.0 1e-06 
0.0 0.8283 0 2.0 1e-06 
0.0 0.8284 0 2.0 1e-06 
0.0 0.8285 0 2.0 1e-06 
0.0 0.8286 0 2.0 1e-06 
0.0 0.8287 0 2.0 1e-06 
0.0 0.8288 0 2.0 1e-06 
0.0 0.8289 0 2.0 1e-06 
0.0 0.829 0 2.0 1e-06 
0.0 0.8291 0 2.0 1e-06 
0.0 0.8292 0 2.0 1e-06 
0.0 0.8293 0 2.0 1e-06 
0.0 0.8294 0 2.0 1e-06 
0.0 0.8295 0 2.0 1e-06 
0.0 0.8296 0 2.0 1e-06 
0.0 0.8297 0 2.0 1e-06 
0.0 0.8298 0 2.0 1e-06 
0.0 0.8299 0 2.0 1e-06 
0.0 0.83 0 2.0 1e-06 
0.0 0.8301 0 2.0 1e-06 
0.0 0.8302 0 2.0 1e-06 
0.0 0.8303 0 2.0 1e-06 
0.0 0.8304 0 2.0 1e-06 
0.0 0.8305 0 2.0 1e-06 
0.0 0.8306 0 2.0 1e-06 
0.0 0.8307 0 2.0 1e-06 
0.0 0.8308 0 2.0 1e-06 
0.0 0.8309 0 2.0 1e-06 
0.0 0.831 0 2.0 1e-06 
0.0 0.8311 0 2.0 1e-06 
0.0 0.8312 0 2.0 1e-06 
0.0 0.8313 0 2.0 1e-06 
0.0 0.8314 0 2.0 1e-06 
0.0 0.8315 0 2.0 1e-06 
0.0 0.8316 0 2.0 1e-06 
0.0 0.8317 0 2.0 1e-06 
0.0 0.8318 0 2.0 1e-06 
0.0 0.8319 0 2.0 1e-06 
0.0 0.832 0 2.0 1e-06 
0.0 0.8321 0 2.0 1e-06 
0.0 0.8322 0 2.0 1e-06 
0.0 0.8323 0 2.0 1e-06 
0.0 0.8324 0 2.0 1e-06 
0.0 0.8325 0 2.0 1e-06 
0.0 0.8326 0 2.0 1e-06 
0.0 0.8327 0 2.0 1e-06 
0.0 0.8328 0 2.0 1e-06 
0.0 0.8329 0 2.0 1e-06 
0.0 0.833 0 2.0 1e-06 
0.0 0.8331 0 2.0 1e-06 
0.0 0.8332 0 2.0 1e-06 
0.0 0.8333 0 2.0 1e-06 
0.0 0.8334 0 2.0 1e-06 
0.0 0.8335 0 2.0 1e-06 
0.0 0.8336 0 2.0 1e-06 
0.0 0.8337 0 2.0 1e-06 
0.0 0.8338 0 2.0 1e-06 
0.0 0.8339 0 2.0 1e-06 
0.0 0.834 0 2.0 1e-06 
0.0 0.8341 0 2.0 1e-06 
0.0 0.8342 0 2.0 1e-06 
0.0 0.8343 0 2.0 1e-06 
0.0 0.8344 0 2.0 1e-06 
0.0 0.8345 0 2.0 1e-06 
0.0 0.8346 0 2.0 1e-06 
0.0 0.8347 0 2.0 1e-06 
0.0 0.8348 0 2.0 1e-06 
0.0 0.8349 0 2.0 1e-06 
0.0 0.835 0 2.0 1e-06 
0.0 0.8351 0 2.0 1e-06 
0.0 0.8352 0 2.0 1e-06 
0.0 0.8353 0 2.0 1e-06 
0.0 0.8354 0 2.0 1e-06 
0.0 0.8355 0 2.0 1e-06 
0.0 0.8356 0 2.0 1e-06 
0.0 0.8357 0 2.0 1e-06 
0.0 0.8358 0 2.0 1e-06 
0.0 0.8359 0 2.0 1e-06 
0.0 0.836 0 2.0 1e-06 
0.0 0.8361 0 2.0 1e-06 
0.0 0.8362 0 2.0 1e-06 
0.0 0.8363 0 2.0 1e-06 
0.0 0.8364 0 2.0 1e-06 
0.0 0.8365 0 2.0 1e-06 
0.0 0.8366 0 2.0 1e-06 
0.0 0.8367 0 2.0 1e-06 
0.0 0.8368 0 2.0 1e-06 
0.0 0.8369 0 2.0 1e-06 
0.0 0.837 0 2.0 1e-06 
0.0 0.8371 0 2.0 1e-06 
0.0 0.8372 0 2.0 1e-06 
0.0 0.8373 0 2.0 1e-06 
0.0 0.8374 0 2.0 1e-06 
0.0 0.8375 0 2.0 1e-06 
0.0 0.8376 0 2.0 1e-06 
0.0 0.8377 0 2.0 1e-06 
0.0 0.8378 0 2.0 1e-06 
0.0 0.8379 0 2.0 1e-06 
0.0 0.838 0 2.0 1e-06 
0.0 0.8381 0 2.0 1e-06 
0.0 0.8382 0 2.0 1e-06 
0.0 0.8383 0 2.0 1e-06 
0.0 0.8384 0 2.0 1e-06 
0.0 0.8385 0 2.0 1e-06 
0.0 0.8386 0 2.0 1e-06 
0.0 0.8387 0 2.0 1e-06 
0.0 0.8388 0 2.0 1e-06 
0.0 0.8389 0 2.0 1e-06 
0.0 0.839 0 2.0 1e-06 
0.0 0.8391 0 2.0 1e-06 
0.0 0.8392 0 2.0 1e-06 
0.0 0.8393 0 2.0 1e-06 
0.0 0.8394 0 2.0 1e-06 
0.0 0.8395 0 2.0 1e-06 
0.0 0.8396 0 2.0 1e-06 
0.0 0.8397 0 2.0 1e-06 
0.0 0.8398 0 2.0 1e-06 
0.0 0.8399 0 2.0 1e-06 
0.0 0.84 0 2.0 1e-06 
0.0 0.8401 0 2.0 1e-06 
0.0 0.8402 0 2.0 1e-06 
0.0 0.8403 0 2.0 1e-06 
0.0 0.8404 0 2.0 1e-06 
0.0 0.8405 0 2.0 1e-06 
0.0 0.8406 0 2.0 1e-06 
0.0 0.8407 0 2.0 1e-06 
0.0 0.8408 0 2.0 1e-06 
0.0 0.8409 0 2.0 1e-06 
0.0 0.841 0 2.0 1e-06 
0.0 0.8411 0 2.0 1e-06 
0.0 0.8412 0 2.0 1e-06 
0.0 0.8413 0 2.0 1e-06 
0.0 0.8414 0 2.0 1e-06 
0.0 0.8415 0 2.0 1e-06 
0.0 0.8416 0 2.0 1e-06 
0.0 0.8417 0 2.0 1e-06 
0.0 0.8418 0 2.0 1e-06 
0.0 0.8419 0 2.0 1e-06 
0.0 0.842 0 2.0 1e-06 
0.0 0.8421 0 2.0 1e-06 
0.0 0.8422 0 2.0 1e-06 
0.0 0.8423 0 2.0 1e-06 
0.0 0.8424 0 2.0 1e-06 
0.0 0.8425 0 2.0 1e-06 
0.0 0.8426 0 2.0 1e-06 
0.0 0.8427 0 2.0 1e-06 
0.0 0.8428 0 2.0 1e-06 
0.0 0.8429 0 2.0 1e-06 
0.0 0.843 0 2.0 1e-06 
0.0 0.8431 0 2.0 1e-06 
0.0 0.8432 0 2.0 1e-06 
0.0 0.8433 0 2.0 1e-06 
0.0 0.8434 0 2.0 1e-06 
0.0 0.8435 0 2.0 1e-06 
0.0 0.8436 0 2.0 1e-06 
0.0 0.8437 0 2.0 1e-06 
0.0 0.8438 0 2.0 1e-06 
0.0 0.8439 0 2.0 1e-06 
0.0 0.844 0 2.0 1e-06 
0.0 0.8441 0 2.0 1e-06 
0.0 0.8442 0 2.0 1e-06 
0.0 0.8443 0 2.0 1e-06 
0.0 0.8444 0 2.0 1e-06 
0.0 0.8445 0 2.0 1e-06 
0.0 0.8446 0 2.0 1e-06 
0.0 0.8447 0 2.0 1e-06 
0.0 0.8448 0 2.0 1e-06 
0.0 0.8449 0 2.0 1e-06 
0.0 0.845 0 2.0 1e-06 
0.0 0.8451 0 2.0 1e-06 
0.0 0.8452 0 2.0 1e-06 
0.0 0.8453 0 2.0 1e-06 
0.0 0.8454 0 2.0 1e-06 
0.0 0.8455 0 2.0 1e-06 
0.0 0.8456 0 2.0 1e-06 
0.0 0.8457 0 2.0 1e-06 
0.0 0.8458 0 2.0 1e-06 
0.0 0.8459 0 2.0 1e-06 
0.0 0.846 0 2.0 1e-06 
0.0 0.8461 0 2.0 1e-06 
0.0 0.8462 0 2.0 1e-06 
0.0 0.8463 0 2.0 1e-06 
0.0 0.8464 0 2.0 1e-06 
0.0 0.8465 0 2.0 1e-06 
0.0 0.8466 0 2.0 1e-06 
0.0 0.8467 0 2.0 1e-06 
0.0 0.8468 0 2.0 1e-06 
0.0 0.8469 0 2.0 1e-06 
0.0 0.847 0 2.0 1e-06 
0.0 0.8471 0 2.0 1e-06 
0.0 0.8472 0 2.0 1e-06 
0.0 0.8473 0 2.0 1e-06 
0.0 0.8474 0 2.0 1e-06 
0.0 0.8475 0 2.0 1e-06 
0.0 0.8476 0 2.0 1e-06 
0.0 0.8477 0 2.0 1e-06 
0.0 0.8478 0 2.0 1e-06 
0.0 0.8479 0 2.0 1e-06 
0.0 0.848 0 2.0 1e-06 
0.0 0.8481 0 2.0 1e-06 
0.0 0.8482 0 2.0 1e-06 
0.0 0.8483 0 2.0 1e-06 
0.0 0.8484 0 2.0 1e-06 
0.0 0.8485 0 2.0 1e-06 
0.0 0.8486 0 2.0 1e-06 
0.0 0.8487 0 2.0 1e-06 
0.0 0.8488 0 2.0 1e-06 
0.0 0.8489 0 2.0 1e-06 
0.0 0.849 0 2.0 1e-06 
0.0 0.8491 0 2.0 1e-06 
0.0 0.8492 0 2.0 1e-06 
0.0 0.8493 0 2.0 1e-06 
0.0 0.8494 0 2.0 1e-06 
0.0 0.8495 0 2.0 1e-06 
0.0 0.8496 0 2.0 1e-06 
0.0 0.8497 0 2.0 1e-06 
0.0 0.8498 0 2.0 1e-06 
0.0 0.8499 0 2.0 1e-06 
0.0 0.85 0 2.0 1e-06 
0.0 0.8501 0 2.0 1e-06 
0.0 0.8502 0 2.0 1e-06 
0.0 0.8503 0 2.0 1e-06 
0.0 0.8504 0 2.0 1e-06 
0.0 0.8505 0 2.0 1e-06 
0.0 0.8506 0 2.0 1e-06 
0.0 0.8507 0 2.0 1e-06 
0.0 0.8508 0 2.0 1e-06 
0.0 0.8509 0 2.0 1e-06 
0.0 0.851 0 2.0 1e-06 
0.0 0.8511 0 2.0 1e-06 
0.0 0.8512 0 2.0 1e-06 
0.0 0.8513 0 2.0 1e-06 
0.0 0.8514 0 2.0 1e-06 
0.0 0.8515 0 2.0 1e-06 
0.0 0.8516 0 2.0 1e-06 
0.0 0.8517 0 2.0 1e-06 
0.0 0.8518 0 2.0 1e-06 
0.0 0.8519 0 2.0 1e-06 
0.0 0.852 0 2.0 1e-06 
0.0 0.8521 0 2.0 1e-06 
0.0 0.8522 0 2.0 1e-06 
0.0 0.8523 0 2.0 1e-06 
0.0 0.8524 0 2.0 1e-06 
0.0 0.8525 0 2.0 1e-06 
0.0 0.8526 0 2.0 1e-06 
0.0 0.8527 0 2.0 1e-06 
0.0 0.8528 0 2.0 1e-06 
0.0 0.8529 0 2.0 1e-06 
0.0 0.853 0 2.0 1e-06 
0.0 0.8531 0 2.0 1e-06 
0.0 0.8532 0 2.0 1e-06 
0.0 0.8533 0 2.0 1e-06 
0.0 0.8534 0 2.0 1e-06 
0.0 0.8535 0 2.0 1e-06 
0.0 0.8536 0 2.0 1e-06 
0.0 0.8537 0 2.0 1e-06 
0.0 0.8538 0 2.0 1e-06 
0.0 0.8539 0 2.0 1e-06 
0.0 0.854 0 2.0 1e-06 
0.0 0.8541 0 2.0 1e-06 
0.0 0.8542 0 2.0 1e-06 
0.0 0.8543 0 2.0 1e-06 
0.0 0.8544 0 2.0 1e-06 
0.0 0.8545 0 2.0 1e-06 
0.0 0.8546 0 2.0 1e-06 
0.0 0.8547 0 2.0 1e-06 
0.0 0.8548 0 2.0 1e-06 
0.0 0.8549 0 2.0 1e-06 
0.0 0.855 0 2.0 1e-06 
0.0 0.8551 0 2.0 1e-06 
0.0 0.8552 0 2.0 1e-06 
0.0 0.8553 0 2.0 1e-06 
0.0 0.8554 0 2.0 1e-06 
0.0 0.8555 0 2.0 1e-06 
0.0 0.8556 0 2.0 1e-06 
0.0 0.8557 0 2.0 1e-06 
0.0 0.8558 0 2.0 1e-06 
0.0 0.8559 0 2.0 1e-06 
0.0 0.856 0 2.0 1e-06 
0.0 0.8561 0 2.0 1e-06 
0.0 0.8562 0 2.0 1e-06 
0.0 0.8563 0 2.0 1e-06 
0.0 0.8564 0 2.0 1e-06 
0.0 0.8565 0 2.0 1e-06 
0.0 0.8566 0 2.0 1e-06 
0.0 0.8567 0 2.0 1e-06 
0.0 0.8568 0 2.0 1e-06 
0.0 0.8569 0 2.0 1e-06 
0.0 0.857 0 2.0 1e-06 
0.0 0.8571 0 2.0 1e-06 
0.0 0.8572 0 2.0 1e-06 
0.0 0.8573 0 2.0 1e-06 
0.0 0.8574 0 2.0 1e-06 
0.0 0.8575 0 2.0 1e-06 
0.0 0.8576 0 2.0 1e-06 
0.0 0.8577 0 2.0 1e-06 
0.0 0.8578 0 2.0 1e-06 
0.0 0.8579 0 2.0 1e-06 
0.0 0.858 0 2.0 1e-06 
0.0 0.8581 0 2.0 1e-06 
0.0 0.8582 0 2.0 1e-06 
0.0 0.8583 0 2.0 1e-06 
0.0 0.8584 0 2.0 1e-06 
0.0 0.8585 0 2.0 1e-06 
0.0 0.8586 0 2.0 1e-06 
0.0 0.8587 0 2.0 1e-06 
0.0 0.8588 0 2.0 1e-06 
0.0 0.8589 0 2.0 1e-06 
0.0 0.859 0 2.0 1e-06 
0.0 0.8591 0 2.0 1e-06 
0.0 0.8592 0 2.0 1e-06 
0.0 0.8593 0 2.0 1e-06 
0.0 0.8594 0 2.0 1e-06 
0.0 0.8595 0 2.0 1e-06 
0.0 0.8596 0 2.0 1e-06 
0.0 0.8597 0 2.0 1e-06 
0.0 0.8598 0 2.0 1e-06 
0.0 0.8599 0 2.0 1e-06 
0.0 0.86 0 2.0 1e-06 
0.0 0.8601 0 2.0 1e-06 
0.0 0.8602 0 2.0 1e-06 
0.0 0.8603 0 2.0 1e-06 
0.0 0.8604 0 2.0 1e-06 
0.0 0.8605 0 2.0 1e-06 
0.0 0.8606 0 2.0 1e-06 
0.0 0.8607 0 2.0 1e-06 
0.0 0.8608 0 2.0 1e-06 
0.0 0.8609 0 2.0 1e-06 
0.0 0.861 0 2.0 1e-06 
0.0 0.8611 0 2.0 1e-06 
0.0 0.8612 0 2.0 1e-06 
0.0 0.8613 0 2.0 1e-06 
0.0 0.8614 0 2.0 1e-06 
0.0 0.8615 0 2.0 1e-06 
0.0 0.8616 0 2.0 1e-06 
0.0 0.8617 0 2.0 1e-06 
0.0 0.8618 0 2.0 1e-06 
0.0 0.8619 0 2.0 1e-06 
0.0 0.862 0 2.0 1e-06 
0.0 0.8621 0 2.0 1e-06 
0.0 0.8622 0 2.0 1e-06 
0.0 0.8623 0 2.0 1e-06 
0.0 0.8624 0 2.0 1e-06 
0.0 0.8625 0 2.0 1e-06 
0.0 0.8626 0 2.0 1e-06 
0.0 0.8627 0 2.0 1e-06 
0.0 0.8628 0 2.0 1e-06 
0.0 0.8629 0 2.0 1e-06 
0.0 0.863 0 2.0 1e-06 
0.0 0.8631 0 2.0 1e-06 
0.0 0.8632 0 2.0 1e-06 
0.0 0.8633 0 2.0 1e-06 
0.0 0.8634 0 2.0 1e-06 
0.0 0.8635 0 2.0 1e-06 
0.0 0.8636 0 2.0 1e-06 
0.0 0.8637 0 2.0 1e-06 
0.0 0.8638 0 2.0 1e-06 
0.0 0.8639 0 2.0 1e-06 
0.0 0.864 0 2.0 1e-06 
0.0 0.8641 0 2.0 1e-06 
0.0 0.8642 0 2.0 1e-06 
0.0 0.8643 0 2.0 1e-06 
0.0 0.8644 0 2.0 1e-06 
0.0 0.8645 0 2.0 1e-06 
0.0 0.8646 0 2.0 1e-06 
0.0 0.8647 0 2.0 1e-06 
0.0 0.8648 0 2.0 1e-06 
0.0 0.8649 0 2.0 1e-06 
0.0 0.865 0 2.0 1e-06 
0.0 0.8651 0 2.0 1e-06 
0.0 0.8652 0 2.0 1e-06 
0.0 0.8653 0 2.0 1e-06 
0.0 0.8654 0 2.0 1e-06 
0.0 0.8655 0 2.0 1e-06 
0.0 0.8656 0 2.0 1e-06 
0.0 0.8657 0 2.0 1e-06 
0.0 0.8658 0 2.0 1e-06 
0.0 0.8659 0 2.0 1e-06 
0.0 0.866 0 2.0 1e-06 
0.0 0.8661 0 2.0 1e-06 
0.0 0.8662 0 2.0 1e-06 
0.0 0.8663 0 2.0 1e-06 
0.0 0.8664 0 2.0 1e-06 
0.0 0.8665 0 2.0 1e-06 
0.0 0.8666 0 2.0 1e-06 
0.0 0.8667 0 2.0 1e-06 
0.0 0.8668 0 2.0 1e-06 
0.0 0.8669 0 2.0 1e-06 
0.0 0.867 0 2.0 1e-06 
0.0 0.8671 0 2.0 1e-06 
0.0 0.8672 0 2.0 1e-06 
0.0 0.8673 0 2.0 1e-06 
0.0 0.8674 0 2.0 1e-06 
0.0 0.8675 0 2.0 1e-06 
0.0 0.8676 0 2.0 1e-06 
0.0 0.8677 0 2.0 1e-06 
0.0 0.8678 0 2.0 1e-06 
0.0 0.8679 0 2.0 1e-06 
0.0 0.868 0 2.0 1e-06 
0.0 0.8681 0 2.0 1e-06 
0.0 0.8682 0 2.0 1e-06 
0.0 0.8683 0 2.0 1e-06 
0.0 0.8684 0 2.0 1e-06 
0.0 0.8685 0 2.0 1e-06 
0.0 0.8686 0 2.0 1e-06 
0.0 0.8687 0 2.0 1e-06 
0.0 0.8688 0 2.0 1e-06 
0.0 0.8689 0 2.0 1e-06 
0.0 0.869 0 2.0 1e-06 
0.0 0.8691 0 2.0 1e-06 
0.0 0.8692 0 2.0 1e-06 
0.0 0.8693 0 2.0 1e-06 
0.0 0.8694 0 2.0 1e-06 
0.0 0.8695 0 2.0 1e-06 
0.0 0.8696 0 2.0 1e-06 
0.0 0.8697 0 2.0 1e-06 
0.0 0.8698 0 2.0 1e-06 
0.0 0.8699 0 2.0 1e-06 
0.0 0.87 0 2.0 1e-06 
0.0 0.8701 0 2.0 1e-06 
0.0 0.8702 0 2.0 1e-06 
0.0 0.8703 0 2.0 1e-06 
0.0 0.8704 0 2.0 1e-06 
0.0 0.8705 0 2.0 1e-06 
0.0 0.8706 0 2.0 1e-06 
0.0 0.8707 0 2.0 1e-06 
0.0 0.8708 0 2.0 1e-06 
0.0 0.8709 0 2.0 1e-06 
0.0 0.871 0 2.0 1e-06 
0.0 0.8711 0 2.0 1e-06 
0.0 0.8712 0 2.0 1e-06 
0.0 0.8713 0 2.0 1e-06 
0.0 0.8714 0 2.0 1e-06 
0.0 0.8715 0 2.0 1e-06 
0.0 0.8716 0 2.0 1e-06 
0.0 0.8717 0 2.0 1e-06 
0.0 0.8718 0 2.0 1e-06 
0.0 0.8719 0 2.0 1e-06 
0.0 0.872 0 2.0 1e-06 
0.0 0.8721 0 2.0 1e-06 
0.0 0.8722 0 2.0 1e-06 
0.0 0.8723 0 2.0 1e-06 
0.0 0.8724 0 2.0 1e-06 
0.0 0.8725 0 2.0 1e-06 
0.0 0.8726 0 2.0 1e-06 
0.0 0.8727 0 2.0 1e-06 
0.0 0.8728 0 2.0 1e-06 
0.0 0.8729 0 2.0 1e-06 
0.0 0.873 0 2.0 1e-06 
0.0 0.8731 0 2.0 1e-06 
0.0 0.8732 0 2.0 1e-06 
0.0 0.8733 0 2.0 1e-06 
0.0 0.8734 0 2.0 1e-06 
0.0 0.8735 0 2.0 1e-06 
0.0 0.8736 0 2.0 1e-06 
0.0 0.8737 0 2.0 1e-06 
0.0 0.8738 0 2.0 1e-06 
0.0 0.8739 0 2.0 1e-06 
0.0 0.874 0 2.0 1e-06 
0.0 0.8741 0 2.0 1e-06 
0.0 0.8742 0 2.0 1e-06 
0.0 0.8743 0 2.0 1e-06 
0.0 0.8744 0 2.0 1e-06 
0.0 0.8745 0 2.0 1e-06 
0.0 0.8746 0 2.0 1e-06 
0.0 0.8747 0 2.0 1e-06 
0.0 0.8748 0 2.0 1e-06 
0.0 0.8749 0 2.0 1e-06 
0.0 0.875 0 2.0 1e-06 
0.0 0.8751 0 2.0 1e-06 
0.0 0.8752 0 2.0 1e-06 
0.0 0.8753 0 2.0 1e-06 
0.0 0.8754 0 2.0 1e-06 
0.0 0.8755 0 2.0 1e-06 
0.0 0.8756 0 2.0 1e-06 
0.0 0.8757 0 2.0 1e-06 
0.0 0.8758 0 2.0 1e-06 
0.0 0.8759 0 2.0 1e-06 
0.0 0.876 0 2.0 1e-06 
0.0 0.8761 0 2.0 1e-06 
0.0 0.8762 0 2.0 1e-06 
0.0 0.8763 0 2.0 1e-06 
0.0 0.8764 0 2.0 1e-06 
0.0 0.8765 0 2.0 1e-06 
0.0 0.8766 0 2.0 1e-06 
0.0 0.8767 0 2.0 1e-06 
0.0 0.8768 0 2.0 1e-06 
0.0 0.8769 0 2.0 1e-06 
0.0 0.877 0 2.0 1e-06 
0.0 0.8771 0 2.0 1e-06 
0.0 0.8772 0 2.0 1e-06 
0.0 0.8773 0 2.0 1e-06 
0.0 0.8774 0 2.0 1e-06 
0.0 0.8775 0 2.0 1e-06 
0.0 0.8776 0 2.0 1e-06 
0.0 0.8777 0 2.0 1e-06 
0.0 0.8778 0 2.0 1e-06 
0.0 0.8779 0 2.0 1e-06 
0.0 0.878 0 2.0 1e-06 
0.0 0.8781 0 2.0 1e-06 
0.0 0.8782 0 2.0 1e-06 
0.0 0.8783 0 2.0 1e-06 
0.0 0.8784 0 2.0 1e-06 
0.0 0.8785 0 2.0 1e-06 
0.0 0.8786 0 2.0 1e-06 
0.0 0.8787 0 2.0 1e-06 
0.0 0.8788 0 2.0 1e-06 
0.0 0.8789 0 2.0 1e-06 
0.0 0.879 0 2.0 1e-06 
0.0 0.8791 0 2.0 1e-06 
0.0 0.8792 0 2.0 1e-06 
0.0 0.8793 0 2.0 1e-06 
0.0 0.8794 0 2.0 1e-06 
0.0 0.8795 0 2.0 1e-06 
0.0 0.8796 0 2.0 1e-06 
0.0 0.8797 0 2.0 1e-06 
0.0 0.8798 0 2.0 1e-06 
0.0 0.8799 0 2.0 1e-06 
0.0 0.88 0 2.0 1e-06 
0.0 0.8801 0 2.0 1e-06 
0.0 0.8802 0 2.0 1e-06 
0.0 0.8803 0 2.0 1e-06 
0.0 0.8804 0 2.0 1e-06 
0.0 0.8805 0 2.0 1e-06 
0.0 0.8806 0 2.0 1e-06 
0.0 0.8807 0 2.0 1e-06 
0.0 0.8808 0 2.0 1e-06 
0.0 0.8809 0 2.0 1e-06 
0.0 0.881 0 2.0 1e-06 
0.0 0.8811 0 2.0 1e-06 
0.0 0.8812 0 2.0 1e-06 
0.0 0.8813 0 2.0 1e-06 
0.0 0.8814 0 2.0 1e-06 
0.0 0.8815 0 2.0 1e-06 
0.0 0.8816 0 2.0 1e-06 
0.0 0.8817 0 2.0 1e-06 
0.0 0.8818 0 2.0 1e-06 
0.0 0.8819 0 2.0 1e-06 
0.0 0.882 0 2.0 1e-06 
0.0 0.8821 0 2.0 1e-06 
0.0 0.8822 0 2.0 1e-06 
0.0 0.8823 0 2.0 1e-06 
0.0 0.8824 0 2.0 1e-06 
0.0 0.8825 0 2.0 1e-06 
0.0 0.8826 0 2.0 1e-06 
0.0 0.8827 0 2.0 1e-06 
0.0 0.8828 0 2.0 1e-06 
0.0 0.8829 0 2.0 1e-06 
0.0 0.883 0 2.0 1e-06 
0.0 0.8831 0 2.0 1e-06 
0.0 0.8832 0 2.0 1e-06 
0.0 0.8833 0 2.0 1e-06 
0.0 0.8834 0 2.0 1e-06 
0.0 0.8835 0 2.0 1e-06 
0.0 0.8836 0 2.0 1e-06 
0.0 0.8837 0 2.0 1e-06 
0.0 0.8838 0 2.0 1e-06 
0.0 0.8839 0 2.0 1e-06 
0.0 0.884 0 2.0 1e-06 
0.0 0.8841 0 2.0 1e-06 
0.0 0.8842 0 2.0 1e-06 
0.0 0.8843 0 2.0 1e-06 
0.0 0.8844 0 2.0 1e-06 
0.0 0.8845 0 2.0 1e-06 
0.0 0.8846 0 2.0 1e-06 
0.0 0.8847 0 2.0 1e-06 
0.0 0.8848 0 2.0 1e-06 
0.0 0.8849 0 2.0 1e-06 
0.0 0.885 0 2.0 1e-06 
0.0 0.8851 0 2.0 1e-06 
0.0 0.8852 0 2.0 1e-06 
0.0 0.8853 0 2.0 1e-06 
0.0 0.8854 0 2.0 1e-06 
0.0 0.8855 0 2.0 1e-06 
0.0 0.8856 0 2.0 1e-06 
0.0 0.8857 0 2.0 1e-06 
0.0 0.8858 0 2.0 1e-06 
0.0 0.8859 0 2.0 1e-06 
0.0 0.886 0 2.0 1e-06 
0.0 0.8861 0 2.0 1e-06 
0.0 0.8862 0 2.0 1e-06 
0.0 0.8863 0 2.0 1e-06 
0.0 0.8864 0 2.0 1e-06 
0.0 0.8865 0 2.0 1e-06 
0.0 0.8866 0 2.0 1e-06 
0.0 0.8867 0 2.0 1e-06 
0.0 0.8868 0 2.0 1e-06 
0.0 0.8869 0 2.0 1e-06 
0.0 0.887 0 2.0 1e-06 
0.0 0.8871 0 2.0 1e-06 
0.0 0.8872 0 2.0 1e-06 
0.0 0.8873 0 2.0 1e-06 
0.0 0.8874 0 2.0 1e-06 
0.0 0.8875 0 2.0 1e-06 
0.0 0.8876 0 2.0 1e-06 
0.0 0.8877 0 2.0 1e-06 
0.0 0.8878 0 2.0 1e-06 
0.0 0.8879 0 2.0 1e-06 
0.0 0.888 0 2.0 1e-06 
0.0 0.8881 0 2.0 1e-06 
0.0 0.8882 0 2.0 1e-06 
0.0 0.8883 0 2.0 1e-06 
0.0 0.8884 0 2.0 1e-06 
0.0 0.8885 0 2.0 1e-06 
0.0 0.8886 0 2.0 1e-06 
0.0 0.8887 0 2.0 1e-06 
0.0 0.8888 0 2.0 1e-06 
0.0 0.8889 0 2.0 1e-06 
0.0 0.889 0 2.0 1e-06 
0.0 0.8891 0 2.0 1e-06 
0.0 0.8892 0 2.0 1e-06 
0.0 0.8893 0 2.0 1e-06 
0.0 0.8894 0 2.0 1e-06 
0.0 0.8895 0 2.0 1e-06 
0.0 0.8896 0 2.0 1e-06 
0.0 0.8897 0 2.0 1e-06 
0.0 0.8898 0 2.0 1e-06 
0.0 0.8899 0 2.0 1e-06 
0.0 0.89 0 2.0 1e-06 
0.0 0.8901 0 2.0 1e-06 
0.0 0.8902 0 2.0 1e-06 
0.0 0.8903 0 2.0 1e-06 
0.0 0.8904 0 2.0 1e-06 
0.0 0.8905 0 2.0 1e-06 
0.0 0.8906 0 2.0 1e-06 
0.0 0.8907 0 2.0 1e-06 
0.0 0.8908 0 2.0 1e-06 
0.0 0.8909 0 2.0 1e-06 
0.0 0.891 0 2.0 1e-06 
0.0 0.8911 0 2.0 1e-06 
0.0 0.8912 0 2.0 1e-06 
0.0 0.8913 0 2.0 1e-06 
0.0 0.8914 0 2.0 1e-06 
0.0 0.8915 0 2.0 1e-06 
0.0 0.8916 0 2.0 1e-06 
0.0 0.8917 0 2.0 1e-06 
0.0 0.8918 0 2.0 1e-06 
0.0 0.8919 0 2.0 1e-06 
0.0 0.892 0 2.0 1e-06 
0.0 0.8921 0 2.0 1e-06 
0.0 0.8922 0 2.0 1e-06 
0.0 0.8923 0 2.0 1e-06 
0.0 0.8924 0 2.0 1e-06 
0.0 0.8925 0 2.0 1e-06 
0.0 0.8926 0 2.0 1e-06 
0.0 0.8927 0 2.0 1e-06 
0.0 0.8928 0 2.0 1e-06 
0.0 0.8929 0 2.0 1e-06 
0.0 0.893 0 2.0 1e-06 
0.0 0.8931 0 2.0 1e-06 
0.0 0.8932 0 2.0 1e-06 
0.0 0.8933 0 2.0 1e-06 
0.0 0.8934 0 2.0 1e-06 
0.0 0.8935 0 2.0 1e-06 
0.0 0.8936 0 2.0 1e-06 
0.0 0.8937 0 2.0 1e-06 
0.0 0.8938 0 2.0 1e-06 
0.0 0.8939 0 2.0 1e-06 
0.0 0.894 0 2.0 1e-06 
0.0 0.8941 0 2.0 1e-06 
0.0 0.8942 0 2.0 1e-06 
0.0 0.8943 0 2.0 1e-06 
0.0 0.8944 0 2.0 1e-06 
0.0 0.8945 0 2.0 1e-06 
0.0 0.8946 0 2.0 1e-06 
0.0 0.8947 0 2.0 1e-06 
0.0 0.8948 0 2.0 1e-06 
0.0 0.8949 0 2.0 1e-06 
0.0 0.895 0 2.0 1e-06 
0.0 0.8951 0 2.0 1e-06 
0.0 0.8952 0 2.0 1e-06 
0.0 0.8953 0 2.0 1e-06 
0.0 0.8954 0 2.0 1e-06 
0.0 0.8955 0 2.0 1e-06 
0.0 0.8956 0 2.0 1e-06 
0.0 0.8957 0 2.0 1e-06 
0.0 0.8958 0 2.0 1e-06 
0.0 0.8959 0 2.0 1e-06 
0.0 0.896 0 2.0 1e-06 
0.0 0.8961 0 2.0 1e-06 
0.0 0.8962 0 2.0 1e-06 
0.0 0.8963 0 2.0 1e-06 
0.0 0.8964 0 2.0 1e-06 
0.0 0.8965 0 2.0 1e-06 
0.0 0.8966 0 2.0 1e-06 
0.0 0.8967 0 2.0 1e-06 
0.0 0.8968 0 2.0 1e-06 
0.0 0.8969 0 2.0 1e-06 
0.0 0.897 0 2.0 1e-06 
0.0 0.8971 0 2.0 1e-06 
0.0 0.8972 0 2.0 1e-06 
0.0 0.8973 0 2.0 1e-06 
0.0 0.8974 0 2.0 1e-06 
0.0 0.8975 0 2.0 1e-06 
0.0 0.8976 0 2.0 1e-06 
0.0 0.8977 0 2.0 1e-06 
0.0 0.8978 0 2.0 1e-06 
0.0 0.8979 0 2.0 1e-06 
0.0 0.898 0 2.0 1e-06 
0.0 0.8981 0 2.0 1e-06 
0.0 0.8982 0 2.0 1e-06 
0.0 0.8983 0 2.0 1e-06 
0.0 0.8984 0 2.0 1e-06 
0.0 0.8985 0 2.0 1e-06 
0.0 0.8986 0 2.0 1e-06 
0.0 0.8987 0 2.0 1e-06 
0.0 0.8988 0 2.0 1e-06 
0.0 0.8989 0 2.0 1e-06 
0.0 0.899 0 2.0 1e-06 
0.0 0.8991 0 2.0 1e-06 
0.0 0.8992 0 2.0 1e-06 
0.0 0.8993 0 2.0 1e-06 
0.0 0.8994 0 2.0 1e-06 
0.0 0.8995 0 2.0 1e-06 
0.0 0.8996 0 2.0 1e-06 
0.0 0.8997 0 2.0 1e-06 
0.0 0.8998 0 2.0 1e-06 
0.0 0.8999 0 2.0 1e-06 
0.0 0.9 0 2.0 1e-06 
0.0 0.9001 0 2.0 1e-06 
0.0 0.9002 0 2.0 1e-06 
0.0 0.9003 0 2.0 1e-06 
0.0 0.9004 0 2.0 1e-06 
0.0 0.9005 0 2.0 1e-06 
0.0 0.9006 0 2.0 1e-06 
0.0 0.9007 0 2.0 1e-06 
0.0 0.9008 0 2.0 1e-06 
0.0 0.9009 0 2.0 1e-06 
0.0 0.901 0 2.0 1e-06 
0.0 0.9011 0 2.0 1e-06 
0.0 0.9012 0 2.0 1e-06 
0.0 0.9013 0 2.0 1e-06 
0.0 0.9014 0 2.0 1e-06 
0.0 0.9015 0 2.0 1e-06 
0.0 0.9016 0 2.0 1e-06 
0.0 0.9017 0 2.0 1e-06 
0.0 0.9018 0 2.0 1e-06 
0.0 0.9019 0 2.0 1e-06 
0.0 0.902 0 2.0 1e-06 
0.0 0.9021 0 2.0 1e-06 
0.0 0.9022 0 2.0 1e-06 
0.0 0.9023 0 2.0 1e-06 
0.0 0.9024 0 2.0 1e-06 
0.0 0.9025 0 2.0 1e-06 
0.0 0.9026 0 2.0 1e-06 
0.0 0.9027 0 2.0 1e-06 
0.0 0.9028 0 2.0 1e-06 
0.0 0.9029 0 2.0 1e-06 
0.0 0.903 0 2.0 1e-06 
0.0 0.9031 0 2.0 1e-06 
0.0 0.9032 0 2.0 1e-06 
0.0 0.9033 0 2.0 1e-06 
0.0 0.9034 0 2.0 1e-06 
0.0 0.9035 0 2.0 1e-06 
0.0 0.9036 0 2.0 1e-06 
0.0 0.9037 0 2.0 1e-06 
0.0 0.9038 0 2.0 1e-06 
0.0 0.9039 0 2.0 1e-06 
0.0 0.904 0 2.0 1e-06 
0.0 0.9041 0 2.0 1e-06 
0.0 0.9042 0 2.0 1e-06 
0.0 0.9043 0 2.0 1e-06 
0.0 0.9044 0 2.0 1e-06 
0.0 0.9045 0 2.0 1e-06 
0.0 0.9046 0 2.0 1e-06 
0.0 0.9047 0 2.0 1e-06 
0.0 0.9048 0 2.0 1e-06 
0.0 0.9049 0 2.0 1e-06 
0.0 0.905 0 2.0 1e-06 
0.0 0.9051 0 2.0 1e-06 
0.0 0.9052 0 2.0 1e-06 
0.0 0.9053 0 2.0 1e-06 
0.0 0.9054 0 2.0 1e-06 
0.0 0.9055 0 2.0 1e-06 
0.0 0.9056 0 2.0 1e-06 
0.0 0.9057 0 2.0 1e-06 
0.0 0.9058 0 2.0 1e-06 
0.0 0.9059 0 2.0 1e-06 
0.0 0.906 0 2.0 1e-06 
0.0 0.9061 0 2.0 1e-06 
0.0 0.9062 0 2.0 1e-06 
0.0 0.9063 0 2.0 1e-06 
0.0 0.9064 0 2.0 1e-06 
0.0 0.9065 0 2.0 1e-06 
0.0 0.9066 0 2.0 1e-06 
0.0 0.9067 0 2.0 1e-06 
0.0 0.9068 0 2.0 1e-06 
0.0 0.9069 0 2.0 1e-06 
0.0 0.907 0 2.0 1e-06 
0.0 0.9071 0 2.0 1e-06 
0.0 0.9072 0 2.0 1e-06 
0.0 0.9073 0 2.0 1e-06 
0.0 0.9074 0 2.0 1e-06 
0.0 0.9075 0 2.0 1e-06 
0.0 0.9076 0 2.0 1e-06 
0.0 0.9077 0 2.0 1e-06 
0.0 0.9078 0 2.0 1e-06 
0.0 0.9079 0 2.0 1e-06 
0.0 0.908 0 2.0 1e-06 
0.0 0.9081 0 2.0 1e-06 
0.0 0.9082 0 2.0 1e-06 
0.0 0.9083 0 2.0 1e-06 
0.0 0.9084 0 2.0 1e-06 
0.0 0.9085 0 2.0 1e-06 
0.0 0.9086 0 2.0 1e-06 
0.0 0.9087 0 2.0 1e-06 
0.0 0.9088 0 2.0 1e-06 
0.0 0.9089 0 2.0 1e-06 
0.0 0.909 0 2.0 1e-06 
0.0 0.9091 0 2.0 1e-06 
0.0 0.9092 0 2.0 1e-06 
0.0 0.9093 0 2.0 1e-06 
0.0 0.9094 0 2.0 1e-06 
0.0 0.9095 0 2.0 1e-06 
0.0 0.9096 0 2.0 1e-06 
0.0 0.9097 0 2.0 1e-06 
0.0 0.9098 0 2.0 1e-06 
0.0 0.9099 0 2.0 1e-06 
0.0 0.91 0 2.0 1e-06 
0.0 0.9101 0 2.0 1e-06 
0.0 0.9102 0 2.0 1e-06 
0.0 0.9103 0 2.0 1e-06 
0.0 0.9104 0 2.0 1e-06 
0.0 0.9105 0 2.0 1e-06 
0.0 0.9106 0 2.0 1e-06 
0.0 0.9107 0 2.0 1e-06 
0.0 0.9108 0 2.0 1e-06 
0.0 0.9109 0 2.0 1e-06 
0.0 0.911 0 2.0 1e-06 
0.0 0.9111 0 2.0 1e-06 
0.0 0.9112 0 2.0 1e-06 
0.0 0.9113 0 2.0 1e-06 
0.0 0.9114 0 2.0 1e-06 
0.0 0.9115 0 2.0 1e-06 
0.0 0.9116 0 2.0 1e-06 
0.0 0.9117 0 2.0 1e-06 
0.0 0.9118 0 2.0 1e-06 
0.0 0.9119 0 2.0 1e-06 
0.0 0.912 0 2.0 1e-06 
0.0 0.9121 0 2.0 1e-06 
0.0 0.9122 0 2.0 1e-06 
0.0 0.9123 0 2.0 1e-06 
0.0 0.9124 0 2.0 1e-06 
0.0 0.9125 0 2.0 1e-06 
0.0 0.9126 0 2.0 1e-06 
0.0 0.9127 0 2.0 1e-06 
0.0 0.9128 0 2.0 1e-06 
0.0 0.9129 0 2.0 1e-06 
0.0 0.913 0 2.0 1e-06 
0.0 0.9131 0 2.0 1e-06 
0.0 0.9132 0 2.0 1e-06 
0.0 0.9133 0 2.0 1e-06 
0.0 0.9134 0 2.0 1e-06 
0.0 0.9135 0 2.0 1e-06 
0.0 0.9136 0 2.0 1e-06 
0.0 0.9137 0 2.0 1e-06 
0.0 0.9138 0 2.0 1e-06 
0.0 0.9139 0 2.0 1e-06 
0.0 0.914 0 2.0 1e-06 
0.0 0.9141 0 2.0 1e-06 
0.0 0.9142 0 2.0 1e-06 
0.0 0.9143 0 2.0 1e-06 
0.0 0.9144 0 2.0 1e-06 
0.0 0.9145 0 2.0 1e-06 
0.0 0.9146 0 2.0 1e-06 
0.0 0.9147 0 2.0 1e-06 
0.0 0.9148 0 2.0 1e-06 
0.0 0.9149 0 2.0 1e-06 
0.0 0.915 0 2.0 1e-06 
0.0 0.9151 0 2.0 1e-06 
0.0 0.9152 0 2.0 1e-06 
0.0 0.9153 0 2.0 1e-06 
0.0 0.9154 0 2.0 1e-06 
0.0 0.9155 0 2.0 1e-06 
0.0 0.9156 0 2.0 1e-06 
0.0 0.9157 0 2.0 1e-06 
0.0 0.9158 0 2.0 1e-06 
0.0 0.9159 0 2.0 1e-06 
0.0 0.916 0 2.0 1e-06 
0.0 0.9161 0 2.0 1e-06 
0.0 0.9162 0 2.0 1e-06 
0.0 0.9163 0 2.0 1e-06 
0.0 0.9164 0 2.0 1e-06 
0.0 0.9165 0 2.0 1e-06 
0.0 0.9166 0 2.0 1e-06 
0.0 0.9167 0 2.0 1e-06 
0.0 0.9168 0 2.0 1e-06 
0.0 0.9169 0 2.0 1e-06 
0.0 0.917 0 2.0 1e-06 
0.0 0.9171 0 2.0 1e-06 
0.0 0.9172 0 2.0 1e-06 
0.0 0.9173 0 2.0 1e-06 
0.0 0.9174 0 2.0 1e-06 
0.0 0.9175 0 2.0 1e-06 
0.0 0.9176 0 2.0 1e-06 
0.0 0.9177 0 2.0 1e-06 
0.0 0.9178 0 2.0 1e-06 
0.0 0.9179 0 2.0 1e-06 
0.0 0.918 0 2.0 1e-06 
0.0 0.9181 0 2.0 1e-06 
0.0 0.9182 0 2.0 1e-06 
0.0 0.9183 0 2.0 1e-06 
0.0 0.9184 0 2.0 1e-06 
0.0 0.9185 0 2.0 1e-06 
0.0 0.9186 0 2.0 1e-06 
0.0 0.9187 0 2.0 1e-06 
0.0 0.9188 0 2.0 1e-06 
0.0 0.9189 0 2.0 1e-06 
0.0 0.919 0 2.0 1e-06 
0.0 0.9191 0 2.0 1e-06 
0.0 0.9192 0 2.0 1e-06 
0.0 0.9193 0 2.0 1e-06 
0.0 0.9194 0 2.0 1e-06 
0.0 0.9195 0 2.0 1e-06 
0.0 0.9196 0 2.0 1e-06 
0.0 0.9197 0 2.0 1e-06 
0.0 0.9198 0 2.0 1e-06 
0.0 0.9199 0 2.0 1e-06 
0.0 0.92 0 2.0 1e-06 
0.0 0.9201 0 2.0 1e-06 
0.0 0.9202 0 2.0 1e-06 
0.0 0.9203 0 2.0 1e-06 
0.0 0.9204 0 2.0 1e-06 
0.0 0.9205 0 2.0 1e-06 
0.0 0.9206 0 2.0 1e-06 
0.0 0.9207 0 2.0 1e-06 
0.0 0.9208 0 2.0 1e-06 
0.0 0.9209 0 2.0 1e-06 
0.0 0.921 0 2.0 1e-06 
0.0 0.9211 0 2.0 1e-06 
0.0 0.9212 0 2.0 1e-06 
0.0 0.9213 0 2.0 1e-06 
0.0 0.9214 0 2.0 1e-06 
0.0 0.9215 0 2.0 1e-06 
0.0 0.9216 0 2.0 1e-06 
0.0 0.9217 0 2.0 1e-06 
0.0 0.9218 0 2.0 1e-06 
0.0 0.9219 0 2.0 1e-06 
0.0 0.922 0 2.0 1e-06 
0.0 0.9221 0 2.0 1e-06 
0.0 0.9222 0 2.0 1e-06 
0.0 0.9223 0 2.0 1e-06 
0.0 0.9224 0 2.0 1e-06 
0.0 0.9225 0 2.0 1e-06 
0.0 0.9226 0 2.0 1e-06 
0.0 0.9227 0 2.0 1e-06 
0.0 0.9228 0 2.0 1e-06 
0.0 0.9229 0 2.0 1e-06 
0.0 0.923 0 2.0 1e-06 
0.0 0.9231 0 2.0 1e-06 
0.0 0.9232 0 2.0 1e-06 
0.0 0.9233 0 2.0 1e-06 
0.0 0.9234 0 2.0 1e-06 
0.0 0.9235 0 2.0 1e-06 
0.0 0.9236 0 2.0 1e-06 
0.0 0.9237 0 2.0 1e-06 
0.0 0.9238 0 2.0 1e-06 
0.0 0.9239 0 2.0 1e-06 
0.0 0.924 0 2.0 1e-06 
0.0 0.9241 0 2.0 1e-06 
0.0 0.9242 0 2.0 1e-06 
0.0 0.9243 0 2.0 1e-06 
0.0 0.9244 0 2.0 1e-06 
0.0 0.9245 0 2.0 1e-06 
0.0 0.9246 0 2.0 1e-06 
0.0 0.9247 0 2.0 1e-06 
0.0 0.9248 0 2.0 1e-06 
0.0 0.9249 0 2.0 1e-06 
0.0 0.925 0 2.0 1e-06 
0.0 0.9251 0 2.0 1e-06 
0.0 0.9252 0 2.0 1e-06 
0.0 0.9253 0 2.0 1e-06 
0.0 0.9254 0 2.0 1e-06 
0.0 0.9255 0 2.0 1e-06 
0.0 0.9256 0 2.0 1e-06 
0.0 0.9257 0 2.0 1e-06 
0.0 0.9258 0 2.0 1e-06 
0.0 0.9259 0 2.0 1e-06 
0.0 0.926 0 2.0 1e-06 
0.0 0.9261 0 2.0 1e-06 
0.0 0.9262 0 2.0 1e-06 
0.0 0.9263 0 2.0 1e-06 
0.0 0.9264 0 2.0 1e-06 
0.0 0.9265 0 2.0 1e-06 
0.0 0.9266 0 2.0 1e-06 
0.0 0.9267 0 2.0 1e-06 
0.0 0.9268 0 2.0 1e-06 
0.0 0.9269 0 2.0 1e-06 
0.0 0.927 0 2.0 1e-06 
0.0 0.9271 0 2.0 1e-06 
0.0 0.9272 0 2.0 1e-06 
0.0 0.9273 0 2.0 1e-06 
0.0 0.9274 0 2.0 1e-06 
0.0 0.9275 0 2.0 1e-06 
0.0 0.9276 0 2.0 1e-06 
0.0 0.9277 0 2.0 1e-06 
0.0 0.9278 0 2.0 1e-06 
0.0 0.9279 0 2.0 1e-06 
0.0 0.928 0 2.0 1e-06 
0.0 0.9281 0 2.0 1e-06 
0.0 0.9282 0 2.0 1e-06 
0.0 0.9283 0 2.0 1e-06 
0.0 0.9284 0 2.0 1e-06 
0.0 0.9285 0 2.0 1e-06 
0.0 0.9286 0 2.0 1e-06 
0.0 0.9287 0 2.0 1e-06 
0.0 0.9288 0 2.0 1e-06 
0.0 0.9289 0 2.0 1e-06 
0.0 0.929 0 2.0 1e-06 
0.0 0.9291 0 2.0 1e-06 
0.0 0.9292 0 2.0 1e-06 
0.0 0.9293 0 2.0 1e-06 
0.0 0.9294 0 2.0 1e-06 
0.0 0.9295 0 2.0 1e-06 
0.0 0.9296 0 2.0 1e-06 
0.0 0.9297 0 2.0 1e-06 
0.0 0.9298 0 2.0 1e-06 
0.0 0.9299 0 2.0 1e-06 
0.0 0.93 0 2.0 1e-06 
0.0 0.9301 0 2.0 1e-06 
0.0 0.9302 0 2.0 1e-06 
0.0 0.9303 0 2.0 1e-06 
0.0 0.9304 0 2.0 1e-06 
0.0 0.9305 0 2.0 1e-06 
0.0 0.9306 0 2.0 1e-06 
0.0 0.9307 0 2.0 1e-06 
0.0 0.9308 0 2.0 1e-06 
0.0 0.9309 0 2.0 1e-06 
0.0 0.931 0 2.0 1e-06 
0.0 0.9311 0 2.0 1e-06 
0.0 0.9312 0 2.0 1e-06 
0.0 0.9313 0 2.0 1e-06 
0.0 0.9314 0 2.0 1e-06 
0.0 0.9315 0 2.0 1e-06 
0.0 0.9316 0 2.0 1e-06 
0.0 0.9317 0 2.0 1e-06 
0.0 0.9318 0 2.0 1e-06 
0.0 0.9319 0 2.0 1e-06 
0.0 0.932 0 2.0 1e-06 
0.0 0.9321 0 2.0 1e-06 
0.0 0.9322 0 2.0 1e-06 
0.0 0.9323 0 2.0 1e-06 
0.0 0.9324 0 2.0 1e-06 
0.0 0.9325 0 2.0 1e-06 
0.0 0.9326 0 2.0 1e-06 
0.0 0.9327 0 2.0 1e-06 
0.0 0.9328 0 2.0 1e-06 
0.0 0.9329 0 2.0 1e-06 
0.0 0.933 0 2.0 1e-06 
0.0 0.9331 0 2.0 1e-06 
0.0 0.9332 0 2.0 1e-06 
0.0 0.9333 0 2.0 1e-06 
0.0 0.9334 0 2.0 1e-06 
0.0 0.9335 0 2.0 1e-06 
0.0 0.9336 0 2.0 1e-06 
0.0 0.9337 0 2.0 1e-06 
0.0 0.9338 0 2.0 1e-06 
0.0 0.9339 0 2.0 1e-06 
0.0 0.934 0 2.0 1e-06 
0.0 0.9341 0 2.0 1e-06 
0.0 0.9342 0 2.0 1e-06 
0.0 0.9343 0 2.0 1e-06 
0.0 0.9344 0 2.0 1e-06 
0.0 0.9345 0 2.0 1e-06 
0.0 0.9346 0 2.0 1e-06 
0.0 0.9347 0 2.0 1e-06 
0.0 0.9348 0 2.0 1e-06 
0.0 0.9349 0 2.0 1e-06 
0.0 0.935 0 2.0 1e-06 
0.0 0.9351 0 2.0 1e-06 
0.0 0.9352 0 2.0 1e-06 
0.0 0.9353 0 2.0 1e-06 
0.0 0.9354 0 2.0 1e-06 
0.0 0.9355 0 2.0 1e-06 
0.0 0.9356 0 2.0 1e-06 
0.0 0.9357 0 2.0 1e-06 
0.0 0.9358 0 2.0 1e-06 
0.0 0.9359 0 2.0 1e-06 
0.0 0.936 0 2.0 1e-06 
0.0 0.9361 0 2.0 1e-06 
0.0 0.9362 0 2.0 1e-06 
0.0 0.9363 0 2.0 1e-06 
0.0 0.9364 0 2.0 1e-06 
0.0 0.9365 0 2.0 1e-06 
0.0 0.9366 0 2.0 1e-06 
0.0 0.9367 0 2.0 1e-06 
0.0 0.9368 0 2.0 1e-06 
0.0 0.9369 0 2.0 1e-06 
0.0 0.937 0 2.0 1e-06 
0.0 0.9371 0 2.0 1e-06 
0.0 0.9372 0 2.0 1e-06 
0.0 0.9373 0 2.0 1e-06 
0.0 0.9374 0 2.0 1e-06 
0.0 0.9375 0 2.0 1e-06 
0.0 0.9376 0 2.0 1e-06 
0.0 0.9377 0 2.0 1e-06 
0.0 0.9378 0 2.0 1e-06 
0.0 0.9379 0 2.0 1e-06 
0.0 0.938 0 2.0 1e-06 
0.0 0.9381 0 2.0 1e-06 
0.0 0.9382 0 2.0 1e-06 
0.0 0.9383 0 2.0 1e-06 
0.0 0.9384 0 2.0 1e-06 
0.0 0.9385 0 2.0 1e-06 
0.0 0.9386 0 2.0 1e-06 
0.0 0.9387 0 2.0 1e-06 
0.0 0.9388 0 2.0 1e-06 
0.0 0.9389 0 2.0 1e-06 
0.0 0.939 0 2.0 1e-06 
0.0 0.9391 0 2.0 1e-06 
0.0 0.9392 0 2.0 1e-06 
0.0 0.9393 0 2.0 1e-06 
0.0 0.9394 0 2.0 1e-06 
0.0 0.9395 0 2.0 1e-06 
0.0 0.9396 0 2.0 1e-06 
0.0 0.9397 0 2.0 1e-06 
0.0 0.9398 0 2.0 1e-06 
0.0 0.9399 0 2.0 1e-06 
0.0 0.94 0 2.0 1e-06 
0.0 0.9401 0 2.0 1e-06 
0.0 0.9402 0 2.0 1e-06 
0.0 0.9403 0 2.0 1e-06 
0.0 0.9404 0 2.0 1e-06 
0.0 0.9405 0 2.0 1e-06 
0.0 0.9406 0 2.0 1e-06 
0.0 0.9407 0 2.0 1e-06 
0.0 0.9408 0 2.0 1e-06 
0.0 0.9409 0 2.0 1e-06 
0.0 0.941 0 2.0 1e-06 
0.0 0.9411 0 2.0 1e-06 
0.0 0.9412 0 2.0 1e-06 
0.0 0.9413 0 2.0 1e-06 
0.0 0.9414 0 2.0 1e-06 
0.0 0.9415 0 2.0 1e-06 
0.0 0.9416 0 2.0 1e-06 
0.0 0.9417 0 2.0 1e-06 
0.0 0.9418 0 2.0 1e-06 
0.0 0.9419 0 2.0 1e-06 
0.0 0.942 0 2.0 1e-06 
0.0 0.9421 0 2.0 1e-06 
0.0 0.9422 0 2.0 1e-06 
0.0 0.9423 0 2.0 1e-06 
0.0 0.9424 0 2.0 1e-06 
0.0 0.9425 0 2.0 1e-06 
0.0 0.9426 0 2.0 1e-06 
0.0 0.9427 0 2.0 1e-06 
0.0 0.9428 0 2.0 1e-06 
0.0 0.9429 0 2.0 1e-06 
0.0 0.943 0 2.0 1e-06 
0.0 0.9431 0 2.0 1e-06 
0.0 0.9432 0 2.0 1e-06 
0.0 0.9433 0 2.0 1e-06 
0.0 0.9434 0 2.0 1e-06 
0.0 0.9435 0 2.0 1e-06 
0.0 0.9436 0 2.0 1e-06 
0.0 0.9437 0 2.0 1e-06 
0.0 0.9438 0 2.0 1e-06 
0.0 0.9439 0 2.0 1e-06 
0.0 0.944 0 2.0 1e-06 
0.0 0.9441 0 2.0 1e-06 
0.0 0.9442 0 2.0 1e-06 
0.0 0.9443 0 2.0 1e-06 
0.0 0.9444 0 2.0 1e-06 
0.0 0.9445 0 2.0 1e-06 
0.0 0.9446 0 2.0 1e-06 
0.0 0.9447 0 2.0 1e-06 
0.0 0.9448 0 2.0 1e-06 
0.0 0.9449 0 2.0 1e-06 
0.0 0.945 0 2.0 1e-06 
0.0 0.9451 0 2.0 1e-06 
0.0 0.9452 0 2.0 1e-06 
0.0 0.9453 0 2.0 1e-06 
0.0 0.9454 0 2.0 1e-06 
0.0 0.9455 0 2.0 1e-06 
0.0 0.9456 0 2.0 1e-06 
0.0 0.9457 0 2.0 1e-06 
0.0 0.9458 0 2.0 1e-06 
0.0 0.9459 0 2.0 1e-06 
0.0 0.946 0 2.0 1e-06 
0.0 0.9461 0 2.0 1e-06 
0.0 0.9462 0 2.0 1e-06 
0.0 0.9463 0 2.0 1e-06 
0.0 0.9464 0 2.0 1e-06 
0.0 0.9465 0 2.0 1e-06 
0.0 0.9466 0 2.0 1e-06 
0.0 0.9467 0 2.0 1e-06 
0.0 0.9468 0 2.0 1e-06 
0.0 0.9469 0 2.0 1e-06 
0.0 0.947 0 2.0 1e-06 
0.0 0.9471 0 2.0 1e-06 
0.0 0.9472 0 2.0 1e-06 
0.0 0.9473 0 2.0 1e-06 
0.0 0.9474 0 2.0 1e-06 
0.0 0.9475 0 2.0 1e-06 
0.0 0.9476 0 2.0 1e-06 
0.0 0.9477 0 2.0 1e-06 
0.0 0.9478 0 2.0 1e-06 
0.0 0.9479 0 2.0 1e-06 
0.0 0.948 0 2.0 1e-06 
0.0 0.9481 0 2.0 1e-06 
0.0 0.9482 0 2.0 1e-06 
0.0 0.9483 0 2.0 1e-06 
0.0 0.9484 0 2.0 1e-06 
0.0 0.9485 0 2.0 1e-06 
0.0 0.9486 0 2.0 1e-06 
0.0 0.9487 0 2.0 1e-06 
0.0 0.9488 0 2.0 1e-06 
0.0 0.9489 0 2.0 1e-06 
0.0 0.949 0 2.0 1e-06 
0.0 0.9491 0 2.0 1e-06 
0.0 0.9492 0 2.0 1e-06 
0.0 0.9493 0 2.0 1e-06 
0.0 0.9494 0 2.0 1e-06 
0.0 0.9495 0 2.0 1e-06 
0.0 0.9496 0 2.0 1e-06 
0.0 0.9497 0 2.0 1e-06 
0.0 0.9498 0 2.0 1e-06 
0.0 0.9499 0 2.0 1e-06 
0.0 0.95 0 2.0 1e-06 
0.0 0.9501 0 2.0 1e-06 
0.0 0.9502 0 2.0 1e-06 
0.0 0.9503 0 2.0 1e-06 
0.0 0.9504 0 2.0 1e-06 
0.0 0.9505 0 2.0 1e-06 
0.0 0.9506 0 2.0 1e-06 
0.0 0.9507 0 2.0 1e-06 
0.0 0.9508 0 2.0 1e-06 
0.0 0.9509 0 2.0 1e-06 
0.0 0.951 0 2.0 1e-06 
0.0 0.9511 0 2.0 1e-06 
0.0 0.9512 0 2.0 1e-06 
0.0 0.9513 0 2.0 1e-06 
0.0 0.9514 0 2.0 1e-06 
0.0 0.9515 0 2.0 1e-06 
0.0 0.9516 0 2.0 1e-06 
0.0 0.9517 0 2.0 1e-06 
0.0 0.9518 0 2.0 1e-06 
0.0 0.9519 0 2.0 1e-06 
0.0 0.952 0 2.0 1e-06 
0.0 0.9521 0 2.0 1e-06 
0.0 0.9522 0 2.0 1e-06 
0.0 0.9523 0 2.0 1e-06 
0.0 0.9524 0 2.0 1e-06 
0.0 0.9525 0 2.0 1e-06 
0.0 0.9526 0 2.0 1e-06 
0.0 0.9527 0 2.0 1e-06 
0.0 0.9528 0 2.0 1e-06 
0.0 0.9529 0 2.0 1e-06 
0.0 0.953 0 2.0 1e-06 
0.0 0.9531 0 2.0 1e-06 
0.0 0.9532 0 2.0 1e-06 
0.0 0.9533 0 2.0 1e-06 
0.0 0.9534 0 2.0 1e-06 
0.0 0.9535 0 2.0 1e-06 
0.0 0.9536 0 2.0 1e-06 
0.0 0.9537 0 2.0 1e-06 
0.0 0.9538 0 2.0 1e-06 
0.0 0.9539 0 2.0 1e-06 
0.0 0.954 0 2.0 1e-06 
0.0 0.9541 0 2.0 1e-06 
0.0 0.9542 0 2.0 1e-06 
0.0 0.9543 0 2.0 1e-06 
0.0 0.9544 0 2.0 1e-06 
0.0 0.9545 0 2.0 1e-06 
0.0 0.9546 0 2.0 1e-06 
0.0 0.9547 0 2.0 1e-06 
0.0 0.9548 0 2.0 1e-06 
0.0 0.9549 0 2.0 1e-06 
0.0 0.955 0 2.0 1e-06 
0.0 0.9551 0 2.0 1e-06 
0.0 0.9552 0 2.0 1e-06 
0.0 0.9553 0 2.0 1e-06 
0.0 0.9554 0 2.0 1e-06 
0.0 0.9555 0 2.0 1e-06 
0.0 0.9556 0 2.0 1e-06 
0.0 0.9557 0 2.0 1e-06 
0.0 0.9558 0 2.0 1e-06 
0.0 0.9559 0 2.0 1e-06 
0.0 0.956 0 2.0 1e-06 
0.0 0.9561 0 2.0 1e-06 
0.0 0.9562 0 2.0 1e-06 
0.0 0.9563 0 2.0 1e-06 
0.0 0.9564 0 2.0 1e-06 
0.0 0.9565 0 2.0 1e-06 
0.0 0.9566 0 2.0 1e-06 
0.0 0.9567 0 2.0 1e-06 
0.0 0.9568 0 2.0 1e-06 
0.0 0.9569 0 2.0 1e-06 
0.0 0.957 0 2.0 1e-06 
0.0 0.9571 0 2.0 1e-06 
0.0 0.9572 0 2.0 1e-06 
0.0 0.9573 0 2.0 1e-06 
0.0 0.9574 0 2.0 1e-06 
0.0 0.9575 0 2.0 1e-06 
0.0 0.9576 0 2.0 1e-06 
0.0 0.9577 0 2.0 1e-06 
0.0 0.9578 0 2.0 1e-06 
0.0 0.9579 0 2.0 1e-06 
0.0 0.958 0 2.0 1e-06 
0.0 0.9581 0 2.0 1e-06 
0.0 0.9582 0 2.0 1e-06 
0.0 0.9583 0 2.0 1e-06 
0.0 0.9584 0 2.0 1e-06 
0.0 0.9585 0 2.0 1e-06 
0.0 0.9586 0 2.0 1e-06 
0.0 0.9587 0 2.0 1e-06 
0.0 0.9588 0 2.0 1e-06 
0.0 0.9589 0 2.0 1e-06 
0.0 0.959 0 2.0 1e-06 
0.0 0.9591 0 2.0 1e-06 
0.0 0.9592 0 2.0 1e-06 
0.0 0.9593 0 2.0 1e-06 
0.0 0.9594 0 2.0 1e-06 
0.0 0.9595 0 2.0 1e-06 
0.0 0.9596 0 2.0 1e-06 
0.0 0.9597 0 2.0 1e-06 
0.0 0.9598 0 2.0 1e-06 
0.0 0.9599 0 2.0 1e-06 
0.0 0.96 0 2.0 1e-06 
0.0 0.9601 0 2.0 1e-06 
0.0 0.9602 0 2.0 1e-06 
0.0 0.9603 0 2.0 1e-06 
0.0 0.9604 0 2.0 1e-06 
0.0 0.9605 0 2.0 1e-06 
0.0 0.9606 0 2.0 1e-06 
0.0 0.9607 0 2.0 1e-06 
0.0 0.9608 0 2.0 1e-06 
0.0 0.9609 0 2.0 1e-06 
0.0 0.961 0 2.0 1e-06 
0.0 0.9611 0 2.0 1e-06 
0.0 0.9612 0 2.0 1e-06 
0.0 0.9613 0 2.0 1e-06 
0.0 0.9614 0 2.0 1e-06 
0.0 0.9615 0 2.0 1e-06 
0.0 0.9616 0 2.0 1e-06 
0.0 0.9617 0 2.0 1e-06 
0.0 0.9618 0 2.0 1e-06 
0.0 0.9619 0 2.0 1e-06 
0.0 0.962 0 2.0 1e-06 
0.0 0.9621 0 2.0 1e-06 
0.0 0.9622 0 2.0 1e-06 
0.0 0.9623 0 2.0 1e-06 
0.0 0.9624 0 2.0 1e-06 
0.0 0.9625 0 2.0 1e-06 
0.0 0.9626 0 2.0 1e-06 
0.0 0.9627 0 2.0 1e-06 
0.0 0.9628 0 2.0 1e-06 
0.0 0.9629 0 2.0 1e-06 
0.0 0.963 0 2.0 1e-06 
0.0 0.9631 0 2.0 1e-06 
0.0 0.9632 0 2.0 1e-06 
0.0 0.9633 0 2.0 1e-06 
0.0 0.9634 0 2.0 1e-06 
0.0 0.9635 0 2.0 1e-06 
0.0 0.9636 0 2.0 1e-06 
0.0 0.9637 0 2.0 1e-06 
0.0 0.9638 0 2.0 1e-06 
0.0 0.9639 0 2.0 1e-06 
0.0 0.964 0 2.0 1e-06 
0.0 0.9641 0 2.0 1e-06 
0.0 0.9642 0 2.0 1e-06 
0.0 0.9643 0 2.0 1e-06 
0.0 0.9644 0 2.0 1e-06 
0.0 0.9645 0 2.0 1e-06 
0.0 0.9646 0 2.0 1e-06 
0.0 0.9647 0 2.0 1e-06 
0.0 0.9648 0 2.0 1e-06 
0.0 0.9649 0 2.0 1e-06 
0.0 0.965 0 2.0 1e-06 
0.0 0.9651 0 2.0 1e-06 
0.0 0.9652 0 2.0 1e-06 
0.0 0.9653 0 2.0 1e-06 
0.0 0.9654 0 2.0 1e-06 
0.0 0.9655 0 2.0 1e-06 
0.0 0.9656 0 2.0 1e-06 
0.0 0.9657 0 2.0 1e-06 
0.0 0.9658 0 2.0 1e-06 
0.0 0.9659 0 2.0 1e-06 
0.0 0.966 0 2.0 1e-06 
0.0 0.9661 0 2.0 1e-06 
0.0 0.9662 0 2.0 1e-06 
0.0 0.9663 0 2.0 1e-06 
0.0 0.9664 0 2.0 1e-06 
0.0 0.9665 0 2.0 1e-06 
0.0 0.9666 0 2.0 1e-06 
0.0 0.9667 0 2.0 1e-06 
0.0 0.9668 0 2.0 1e-06 
0.0 0.9669 0 2.0 1e-06 
0.0 0.967 0 2.0 1e-06 
0.0 0.9671 0 2.0 1e-06 
0.0 0.9672 0 2.0 1e-06 
0.0 0.9673 0 2.0 1e-06 
0.0 0.9674 0 2.0 1e-06 
0.0 0.9675 0 2.0 1e-06 
0.0 0.9676 0 2.0 1e-06 
0.0 0.9677 0 2.0 1e-06 
0.0 0.9678 0 2.0 1e-06 
0.0 0.9679 0 2.0 1e-06 
0.0 0.968 0 2.0 1e-06 
0.0 0.9681 0 2.0 1e-06 
0.0 0.9682 0 2.0 1e-06 
0.0 0.9683 0 2.0 1e-06 
0.0 0.9684 0 2.0 1e-06 
0.0 0.9685 0 2.0 1e-06 
0.0 0.9686 0 2.0 1e-06 
0.0 0.9687 0 2.0 1e-06 
0.0 0.9688 0 2.0 1e-06 
0.0 0.9689 0 2.0 1e-06 
0.0 0.969 0 2.0 1e-06 
0.0 0.9691 0 2.0 1e-06 
0.0 0.9692 0 2.0 1e-06 
0.0 0.9693 0 2.0 1e-06 
0.0 0.9694 0 2.0 1e-06 
0.0 0.9695 0 2.0 1e-06 
0.0 0.9696 0 2.0 1e-06 
0.0 0.9697 0 2.0 1e-06 
0.0 0.9698 0 2.0 1e-06 
0.0 0.9699 0 2.0 1e-06 
0.0 0.97 0 2.0 1e-06 
0.0 0.9701 0 2.0 1e-06 
0.0 0.9702 0 2.0 1e-06 
0.0 0.9703 0 2.0 1e-06 
0.0 0.9704 0 2.0 1e-06 
0.0 0.9705 0 2.0 1e-06 
0.0 0.9706 0 2.0 1e-06 
0.0 0.9707 0 2.0 1e-06 
0.0 0.9708 0 2.0 1e-06 
0.0 0.9709 0 2.0 1e-06 
0.0 0.971 0 2.0 1e-06 
0.0 0.9711 0 2.0 1e-06 
0.0 0.9712 0 2.0 1e-06 
0.0 0.9713 0 2.0 1e-06 
0.0 0.9714 0 2.0 1e-06 
0.0 0.9715 0 2.0 1e-06 
0.0 0.9716 0 2.0 1e-06 
0.0 0.9717 0 2.0 1e-06 
0.0 0.9718 0 2.0 1e-06 
0.0 0.9719 0 2.0 1e-06 
0.0 0.972 0 2.0 1e-06 
0.0 0.9721 0 2.0 1e-06 
0.0 0.9722 0 2.0 1e-06 
0.0 0.9723 0 2.0 1e-06 
0.0 0.9724 0 2.0 1e-06 
0.0 0.9725 0 2.0 1e-06 
0.0 0.9726 0 2.0 1e-06 
0.0 0.9727 0 2.0 1e-06 
0.0 0.9728 0 2.0 1e-06 
0.0 0.9729 0 2.0 1e-06 
0.0 0.973 0 2.0 1e-06 
0.0 0.9731 0 2.0 1e-06 
0.0 0.9732 0 2.0 1e-06 
0.0 0.9733 0 2.0 1e-06 
0.0 0.9734 0 2.0 1e-06 
0.0 0.9735 0 2.0 1e-06 
0.0 0.9736 0 2.0 1e-06 
0.0 0.9737 0 2.0 1e-06 
0.0 0.9738 0 2.0 1e-06 
0.0 0.9739 0 2.0 1e-06 
0.0 0.974 0 2.0 1e-06 
0.0 0.9741 0 2.0 1e-06 
0.0 0.9742 0 2.0 1e-06 
0.0 0.9743 0 2.0 1e-06 
0.0 0.9744 0 2.0 1e-06 
0.0 0.9745 0 2.0 1e-06 
0.0 0.9746 0 2.0 1e-06 
0.0 0.9747 0 2.0 1e-06 
0.0 0.9748 0 2.0 1e-06 
0.0 0.9749 0 2.0 1e-06 
0.0 0.975 0 2.0 1e-06 
0.0 0.9751 0 2.0 1e-06 
0.0 0.9752 0 2.0 1e-06 
0.0 0.9753 0 2.0 1e-06 
0.0 0.9754 0 2.0 1e-06 
0.0 0.9755 0 2.0 1e-06 
0.0 0.9756 0 2.0 1e-06 
0.0 0.9757 0 2.0 1e-06 
0.0 0.9758 0 2.0 1e-06 
0.0 0.9759 0 2.0 1e-06 
0.0 0.976 0 2.0 1e-06 
0.0 0.9761 0 2.0 1e-06 
0.0 0.9762 0 2.0 1e-06 
0.0 0.9763 0 2.0 1e-06 
0.0 0.9764 0 2.0 1e-06 
0.0 0.9765 0 2.0 1e-06 
0.0 0.9766 0 2.0 1e-06 
0.0 0.9767 0 2.0 1e-06 
0.0 0.9768 0 2.0 1e-06 
0.0 0.9769 0 2.0 1e-06 
0.0 0.977 0 2.0 1e-06 
0.0 0.9771 0 2.0 1e-06 
0.0 0.9772 0 2.0 1e-06 
0.0 0.9773 0 2.0 1e-06 
0.0 0.9774 0 2.0 1e-06 
0.0 0.9775 0 2.0 1e-06 
0.0 0.9776 0 2.0 1e-06 
0.0 0.9777 0 2.0 1e-06 
0.0 0.9778 0 2.0 1e-06 
0.0 0.9779 0 2.0 1e-06 
0.0 0.978 0 2.0 1e-06 
0.0 0.9781 0 2.0 1e-06 
0.0 0.9782 0 2.0 1e-06 
0.0 0.9783 0 2.0 1e-06 
0.0 0.9784 0 2.0 1e-06 
0.0 0.9785 0 2.0 1e-06 
0.0 0.9786 0 2.0 1e-06 
0.0 0.9787 0 2.0 1e-06 
0.0 0.9788 0 2.0 1e-06 
0.0 0.9789 0 2.0 1e-06 
0.0 0.979 0 2.0 1e-06 
0.0 0.9791 0 2.0 1e-06 
0.0 0.9792 0 2.0 1e-06 
0.0 0.9793 0 2.0 1e-06 
0.0 0.9794 0 2.0 1e-06 
0.0 0.9795 0 2.0 1e-06 
0.0 0.9796 0 2.0 1e-06 
0.0 0.9797 0 2.0 1e-06 
0.0 0.9798 0 2.0 1e-06 
0.0 0.9799 0 2.0 1e-06 
0.0 0.98 0 2.0 1e-06 
0.0 0.9801 0 2.0 1e-06 
0.0 0.9802 0 2.0 1e-06 
0.0 0.9803 0 2.0 1e-06 
0.0 0.9804 0 2.0 1e-06 
0.0 0.9805 0 2.0 1e-06 
0.0 0.9806 0 2.0 1e-06 
0.0 0.9807 0 2.0 1e-06 
0.0 0.9808 0 2.0 1e-06 
0.0 0.9809 0 2.0 1e-06 
0.0 0.981 0 2.0 1e-06 
0.0 0.9811 0 2.0 1e-06 
0.0 0.9812 0 2.0 1e-06 
0.0 0.9813 0 2.0 1e-06 
0.0 0.9814 0 2.0 1e-06 
0.0 0.9815 0 2.0 1e-06 
0.0 0.9816 0 2.0 1e-06 
0.0 0.9817 0 2.0 1e-06 
0.0 0.9818 0 2.0 1e-06 
0.0 0.9819 0 2.0 1e-06 
0.0 0.982 0 2.0 1e-06 
0.0 0.9821 0 2.0 1e-06 
0.0 0.9822 0 2.0 1e-06 
0.0 0.9823 0 2.0 1e-06 
0.0 0.9824 0 2.0 1e-06 
0.0 0.9825 0 2.0 1e-06 
0.0 0.9826 0 2.0 1e-06 
0.0 0.9827 0 2.0 1e-06 
0.0 0.9828 0 2.0 1e-06 
0.0 0.9829 0 2.0 1e-06 
0.0 0.983 0 2.0 1e-06 
0.0 0.9831 0 2.0 1e-06 
0.0 0.9832 0 2.0 1e-06 
0.0 0.9833 0 2.0 1e-06 
0.0 0.9834 0 2.0 1e-06 
0.0 0.9835 0 2.0 1e-06 
0.0 0.9836 0 2.0 1e-06 
0.0 0.9837 0 2.0 1e-06 
0.0 0.9838 0 2.0 1e-06 
0.0 0.9839 0 2.0 1e-06 
0.0 0.984 0 2.0 1e-06 
0.0 0.9841 0 2.0 1e-06 
0.0 0.9842 0 2.0 1e-06 
0.0 0.9843 0 2.0 1e-06 
0.0 0.9844 0 2.0 1e-06 
0.0 0.9845 0 2.0 1e-06 
0.0 0.9846 0 2.0 1e-06 
0.0 0.9847 0 2.0 1e-06 
0.0 0.9848 0 2.0 1e-06 
0.0 0.9849 0 2.0 1e-06 
0.0 0.985 0 2.0 1e-06 
0.0 0.9851 0 2.0 1e-06 
0.0 0.9852 0 2.0 1e-06 
0.0 0.9853 0 2.0 1e-06 
0.0 0.9854 0 2.0 1e-06 
0.0 0.9855 0 2.0 1e-06 
0.0 0.9856 0 2.0 1e-06 
0.0 0.9857 0 2.0 1e-06 
0.0 0.9858 0 2.0 1e-06 
0.0 0.9859 0 2.0 1e-06 
0.0 0.986 0 2.0 1e-06 
0.0 0.9861 0 2.0 1e-06 
0.0 0.9862 0 2.0 1e-06 
0.0 0.9863 0 2.0 1e-06 
0.0 0.9864 0 2.0 1e-06 
0.0 0.9865 0 2.0 1e-06 
0.0 0.9866 0 2.0 1e-06 
0.0 0.9867 0 2.0 1e-06 
0.0 0.9868 0 2.0 1e-06 
0.0 0.9869 0 2.0 1e-06 
0.0 0.987 0 2.0 1e-06 
0.0 0.9871 0 2.0 1e-06 
0.0 0.9872 0 2.0 1e-06 
0.0 0.9873 0 2.0 1e-06 
0.0 0.9874 0 2.0 1e-06 
0.0 0.9875 0 2.0 1e-06 
0.0 0.9876 0 2.0 1e-06 
0.0 0.9877 0 2.0 1e-06 
0.0 0.9878 0 2.0 1e-06 
0.0 0.9879 0 2.0 1e-06 
0.0 0.988 0 2.0 1e-06 
0.0 0.9881 0 2.0 1e-06 
0.0 0.9882 0 2.0 1e-06 
0.0 0.9883 0 2.0 1e-06 
0.0 0.9884 0 2.0 1e-06 
0.0 0.9885 0 2.0 1e-06 
0.0 0.9886 0 2.0 1e-06 
0.0 0.9887 0 2.0 1e-06 
0.0 0.9888 0 2.0 1e-06 
0.0 0.9889 0 2.0 1e-06 
0.0 0.989 0 2.0 1e-06 
0.0 0.9891 0 2.0 1e-06 
0.0 0.9892 0 2.0 1e-06 
0.0 0.9893 0 2.0 1e-06 
0.0 0.9894 0 2.0 1e-06 
0.0 0.9895 0 2.0 1e-06 
0.0 0.9896 0 2.0 1e-06 
0.0 0.9897 0 2.0 1e-06 
0.0 0.9898 0 2.0 1e-06 
0.0 0.9899 0 2.0 1e-06 
0.0 0.99 0 2.0 1e-06 
0.0 0.9901 0 2.0 1e-06 
0.0 0.9902 0 2.0 1e-06 
0.0 0.9903 0 2.0 1e-06 
0.0 0.9904 0 2.0 1e-06 
0.0 0.9905 0 2.0 1e-06 
0.0 0.9906 0 2.0 1e-06 
0.0 0.9907 0 2.0 1e-06 
0.0 0.9908 0 2.0 1e-06 
0.0 0.9909 0 2.0 1e-06 
0.0 0.991 0 2.0 1e-06 
0.0 0.9911 0 2.0 1e-06 
0.0 0.9912 0 2.0 1e-06 
0.0 0.9913 0 2.0 1e-06 
0.0 0.9914 0 2.0 1e-06 
0.0 0.9915 0 2.0 1e-06 
0.0 0.9916 0 2.0 1e-06 
0.0 0.9917 0 2.0 1e-06 
0.0 0.9918 0 2.0 1e-06 
0.0 0.9919 0 2.0 1e-06 
0.0 0.992 0 2.0 1e-06 
0.0 0.9921 0 2.0 1e-06 
0.0 0.9922 0 2.0 1e-06 
0.0 0.9923 0 2.0 1e-06 
0.0 0.9924 0 2.0 1e-06 
0.0 0.9925 0 2.0 1e-06 
0.0 0.9926 0 2.0 1e-06 
0.0 0.9927 0 2.0 1e-06 
0.0 0.9928 0 2.0 1e-06 
0.0 0.9929 0 2.0 1e-06 
0.0 0.993 0 2.0 1e-06 
0.0 0.9931 0 2.0 1e-06 
0.0 0.9932 0 2.0 1e-06 
0.0 0.9933 0 2.0 1e-06 
0.0 0.9934 0 2.0 1e-06 
0.0 0.9935 0 2.0 1e-06 
0.0 0.9936 0 2.0 1e-06 
0.0 0.9937 0 2.0 1e-06 
0.0 0.9938 0 2.0 1e-06 
0.0 0.9939 0 2.0 1e-06 
0.0 0.994 0 2.0 1e-06 
0.0 0.9941 0 2.0 1e-06 
0.0 0.9942 0 2.0 1e-06 
0.0 0.9943 0 2.0 1e-06 
0.0 0.9944 0 2.0 1e-06 
0.0 0.9945 0 2.0 1e-06 
0.0 0.9946 0 2.0 1e-06 
0.0 0.9947 0 2.0 1e-06 
0.0 0.9948 0 2.0 1e-06 
0.0 0.9949 0 2.0 1e-06 
0.0 0.995 0 2.0 1e-06 
0.0 0.9951 0 2.0 1e-06 
0.0 0.9952 0 2.0 1e-06 
0.0 0.9953 0 2.0 1e-06 
0.0 0.9954 0 2.0 1e-06 
0.0 0.9955 0 2.0 1e-06 
0.0 0.9956 0 2.0 1e-06 
0.0 0.9957 0 2.0 1e-06 
0.0 0.9958 0 2.0 1e-06 
0.0 0.9959 0 2.0 1e-06 
0.0 0.996 0 2.0 1e-06 
0.0 0.9961 0 2.0 1e-06 
0.0 0.9962 0 2.0 1e-06 
0.0 0.9963 0 2.0 1e-06 
0.0 0.9964 0 2.0 1e-06 
0.0 0.9965 0 2.0 1e-06 
0.0 0.9966 0 2.0 1e-06 
0.0 0.9967 0 2.0 1e-06 
0.0 0.9968 0 2.0 1e-06 
0.0 0.9969 0 2.0 1e-06 
0.0 0.997 0 2.0 1e-06 
0.0 0.9971 0 2.0 1e-06 
0.0 0.9972 0 2.0 1e-06 
0.0 0.9973 0 2.0 1e-06 
0.0 0.9974 0 2.0 1e-06 
0.0 0.9975 0 2.0 1e-06 
0.0 0.9976 0 2.0 1e-06 
0.0 0.9977 0 2.0 1e-06 
0.0 0.9978 0 2.0 1e-06 
0.0 0.9979 0 2.0 1e-06 
0.0 0.998 0 2.0 1e-06 
0.0 0.9981 0 2.0 1e-06 
0.0 0.9982 0 2.0 1e-06 
0.0 0.9983 0 2.0 1e-06 
0.0 0.9984 0 2.0 1e-06 
0.0 0.9985 0 2.0 1e-06 
0.0 0.9986 0 2.0 1e-06 
0.0 0.9987 0 2.0 1e-06 
0.0 0.9988 0 2.0 1e-06 
0.0 0.9989 0 2.0 1e-06 
0.0 0.999 0 2.0 1e-06 
0.0 0.9991 0 2.0 1e-06 
0.0 0.9992 0 2.0 1e-06 
0.0 0.9993 0 2.0 1e-06 
0.0 0.9994 0 2.0 1e-06 
0.0 0.9995 0 2.0 1e-06 
0.0 0.9996 0 2.0 1e-06 
0.0 0.9997 0 2.0 1e-06 
0.0 0.9998 0 2.0 1e-06 
0.0 0.9999 0 2.0 1e-06 
0.0 1.0 0 2.0 1e-06 
0.0 1.0001 0 2.0 1e-06 
0.0 1.0002 0 2.0 1e-06 
0.0 1.0003 0 2.0 1e-06 
0.0 1.0004 0 2.0 1e-06 
0.0 1.0005 0 2.0 1e-06 
0.0 1.0006 0 2.0 1e-06 
0.0 1.0007 0 2.0 1e-06 
0.0 1.0008 0 2.0 1e-06 
0.0 1.0009 0 2.0 1e-06 
0.0 1.001 0 2.0 1e-06 
0.0 1.0011 0 2.0 1e-06 
0.0 1.0012 0 2.0 1e-06 
0.0 1.0013 0 2.0 1e-06 
0.0 1.0014 0 2.0 1e-06 
0.0 1.0015 0 2.0 1e-06 
0.0 1.0016 0 2.0 1e-06 
0.0 1.0017 0 2.0 1e-06 
0.0 1.0018 0 2.0 1e-06 
0.0 1.0019 0 2.0 1e-06 
0.0 1.002 0 2.0 1e-06 
0.0 1.0021 0 2.0 1e-06 
0.0 1.0022 0 2.0 1e-06 
0.0 1.0023 0 2.0 1e-06 
0.0 1.0024 0 2.0 1e-06 
0.0 1.0025 0 2.0 1e-06 
0.0 1.0026 0 2.0 1e-06 
0.0 1.0027 0 2.0 1e-06 
0.0 1.0028 0 2.0 1e-06 
0.0 1.0029 0 2.0 1e-06 
0.0 1.003 0 2.0 1e-06 
0.0 1.0031 0 2.0 1e-06 
0.0 1.0032 0 2.0 1e-06 
0.0 1.0033 0 2.0 1e-06 
0.0 1.0034 0 2.0 1e-06 
0.0 1.0035 0 2.0 1e-06 
0.0 1.0036 0 2.0 1e-06 
0.0 1.0037 0 2.0 1e-06 
0.0 1.0038 0 2.0 1e-06 
0.0 1.0039 0 2.0 1e-06 
0.0 1.004 0 2.0 1e-06 
0.0 1.0041 0 2.0 1e-06 
0.0 1.0042 0 2.0 1e-06 
0.0 1.0043 0 2.0 1e-06 
0.0 1.0044 0 2.0 1e-06 
0.0 1.0045 0 2.0 1e-06 
0.0 1.0046 0 2.0 1e-06 
0.0 1.0047 0 2.0 1e-06 
0.0 1.0048 0 2.0 1e-06 
0.0 1.0049 0 2.0 1e-06 
0.0 1.005 0 2.0 1e-06 
0.0 1.0051 0 2.0 1e-06 
0.0 1.0052 0 2.0 1e-06 
0.0 1.0053 0 2.0 1e-06 
0.0 1.0054 0 2.0 1e-06 
0.0 1.0055 0 2.0 1e-06 
0.0 1.0056 0 2.0 1e-06 
0.0 1.0057 0 2.0 1e-06 
0.0 1.0058 0 2.0 1e-06 
0.0 1.0059 0 2.0 1e-06 
0.0 1.006 0 2.0 1e-06 
0.0 1.0061 0 2.0 1e-06 
0.0 1.0062 0 2.0 1e-06 
0.0 1.0063 0 2.0 1e-06 
0.0 1.0064 0 2.0 1e-06 
0.0 1.0065 0 2.0 1e-06 
0.0 1.0066 0 2.0 1e-06 
0.0 1.0067 0 2.0 1e-06 
0.0 1.0068 0 2.0 1e-06 
0.0 1.0069 0 2.0 1e-06 
0.0 1.007 0 2.0 1e-06 
0.0 1.0071 0 2.0 1e-06 
0.0 1.0072 0 2.0 1e-06 
0.0 1.0073 0 2.0 1e-06 
0.0 1.0074 0 2.0 1e-06 
0.0 1.0075 0 2.0 1e-06 
0.0 1.0076 0 2.0 1e-06 
0.0 1.0077 0 2.0 1e-06 
0.0 1.0078 0 2.0 1e-06 
0.0 1.0079 0 2.0 1e-06 
0.0 1.008 0 2.0 1e-06 
0.0 1.0081 0 2.0 1e-06 
0.0 1.0082 0 2.0 1e-06 
0.0 1.0083 0 2.0 1e-06 
0.0 1.0084 0 2.0 1e-06 
0.0 1.0085 0 2.0 1e-06 
0.0 1.0086 0 2.0 1e-06 
0.0 1.0087 0 2.0 1e-06 
0.0 1.0088 0 2.0 1e-06 
0.0 1.0089 0 2.0 1e-06 
0.0 1.009 0 2.0 1e-06 
0.0 1.0091 0 2.0 1e-06 
0.0 1.0092 0 2.0 1e-06 
0.0 1.0093 0 2.0 1e-06 
0.0 1.0094 0 2.0 1e-06 
0.0 1.0095 0 2.0 1e-06 
0.0 1.0096 0 2.0 1e-06 
0.0 1.0097 0 2.0 1e-06 
0.0 1.0098 0 2.0 1e-06 
0.0 1.0099 0 2.0 1e-06 
0.0 1.01 0 2.0 1e-06 
0.0 1.0101 0 2.0 1e-06 
0.0 1.0102 0 2.0 1e-06 
0.0 1.0103 0 2.0 1e-06 
0.0 1.0104 0 2.0 1e-06 
0.0 1.0105 0 2.0 1e-06 
0.0 1.0106 0 2.0 1e-06 
0.0 1.0107 0 2.0 1e-06 
0.0 1.0108 0 2.0 1e-06 
0.0 1.0109 0 2.0 1e-06 
0.0 1.011 0 2.0 1e-06 
0.0 1.0111 0 2.0 1e-06 
0.0 1.0112 0 2.0 1e-06 
0.0 1.0113 0 2.0 1e-06 
0.0 1.0114 0 2.0 1e-06 
0.0 1.0115 0 2.0 1e-06 
0.0 1.0116 0 2.0 1e-06 
0.0 1.0117 0 2.0 1e-06 
0.0 1.0118 0 2.0 1e-06 
0.0 1.0119 0 2.0 1e-06 
0.0 1.012 0 2.0 1e-06 
0.0 1.0121 0 2.0 1e-06 
0.0 1.0122 0 2.0 1e-06 
0.0 1.0123 0 2.0 1e-06 
0.0 1.0124 0 2.0 1e-06 
0.0 1.0125 0 2.0 1e-06 
0.0 1.0126 0 2.0 1e-06 
0.0 1.0127 0 2.0 1e-06 
0.0 1.0128 0 2.0 1e-06 
0.0 1.0129 0 2.0 1e-06 
0.0 1.013 0 2.0 1e-06 
0.0 1.0131 0 2.0 1e-06 
0.0 1.0132 0 2.0 1e-06 
0.0 1.0133 0 2.0 1e-06 
0.0 1.0134 0 2.0 1e-06 
0.0 1.0135 0 2.0 1e-06 
0.0 1.0136 0 2.0 1e-06 
0.0 1.0137 0 2.0 1e-06 
0.0 1.0138 0 2.0 1e-06 
0.0 1.0139 0 2.0 1e-06 
0.0 1.014 0 2.0 1e-06 
0.0 1.0141 0 2.0 1e-06 
0.0 1.0142 0 2.0 1e-06 
0.0 1.0143 0 2.0 1e-06 
0.0 1.0144 0 2.0 1e-06 
0.0 1.0145 0 2.0 1e-06 
0.0 1.0146 0 2.0 1e-06 
0.0 1.0147 0 2.0 1e-06 
0.0 1.0148 0 2.0 1e-06 
0.0 1.0149 0 2.0 1e-06 
0.0 1.015 0 2.0 1e-06 
0.0 1.0151 0 2.0 1e-06 
0.0 1.0152 0 2.0 1e-06 
0.0 1.0153 0 2.0 1e-06 
0.0 1.0154 0 2.0 1e-06 
0.0 1.0155 0 2.0 1e-06 
0.0 1.0156 0 2.0 1e-06 
0.0 1.0157 0 2.0 1e-06 
0.0 1.0158 0 2.0 1e-06 
0.0 1.0159 0 2.0 1e-06 
0.0 1.016 0 2.0 1e-06 
0.0 1.0161 0 2.0 1e-06 
0.0 1.0162 0 2.0 1e-06 
0.0 1.0163 0 2.0 1e-06 
0.0 1.0164 0 2.0 1e-06 
0.0 1.0165 0 2.0 1e-06 
0.0 1.0166 0 2.0 1e-06 
0.0 1.0167 0 2.0 1e-06 
0.0 1.0168 0 2.0 1e-06 
0.0 1.0169 0 2.0 1e-06 
0.0 1.017 0 2.0 1e-06 
0.0 1.0171 0 2.0 1e-06 
0.0 1.0172 0 2.0 1e-06 
0.0 1.0173 0 2.0 1e-06 
0.0 1.0174 0 2.0 1e-06 
0.0 1.0175 0 2.0 1e-06 
0.0 1.0176 0 2.0 1e-06 
0.0 1.0177 0 2.0 1e-06 
0.0 1.0178 0 2.0 1e-06 
0.0 1.0179 0 2.0 1e-06 
0.0 1.018 0 2.0 1e-06 
0.0 1.0181 0 2.0 1e-06 
0.0 1.0182 0 2.0 1e-06 
0.0 1.0183 0 2.0 1e-06 
0.0 1.0184 0 2.0 1e-06 
0.0 1.0185 0 2.0 1e-06 
0.0 1.0186 0 2.0 1e-06 
0.0 1.0187 0 2.0 1e-06 
0.0 1.0188 0 2.0 1e-06 
0.0 1.0189 0 2.0 1e-06 
0.0 1.019 0 2.0 1e-06 
0.0 1.0191 0 2.0 1e-06 
0.0 1.0192 0 2.0 1e-06 
0.0 1.0193 0 2.0 1e-06 
0.0 1.0194 0 2.0 1e-06 
0.0 1.0195 0 2.0 1e-06 
0.0 1.0196 0 2.0 1e-06 
0.0 1.0197 0 2.0 1e-06 
0.0 1.0198 0 2.0 1e-06 
0.0 1.0199 0 2.0 1e-06 
0.0 1.02 0 2.0 1e-06 
0.0 1.0201 0 2.0 1e-06 
0.0 1.0202 0 2.0 1e-06 
0.0 1.0203 0 2.0 1e-06 
0.0 1.0204 0 2.0 1e-06 
0.0 1.0205 0 2.0 1e-06 
0.0 1.0206 0 2.0 1e-06 
0.0 1.0207 0 2.0 1e-06 
0.0 1.0208 0 2.0 1e-06 
0.0 1.0209 0 2.0 1e-06 
0.0 1.021 0 2.0 1e-06 
0.0 1.0211 0 2.0 1e-06 
0.0 1.0212 0 2.0 1e-06 
0.0 1.0213 0 2.0 1e-06 
0.0 1.0214 0 2.0 1e-06 
0.0 1.0215 0 2.0 1e-06 
0.0 1.0216 0 2.0 1e-06 
0.0 1.0217 0 2.0 1e-06 
0.0 1.0218 0 2.0 1e-06 
0.0 1.0219 0 2.0 1e-06 
0.0 1.022 0 2.0 1e-06 
0.0 1.0221 0 2.0 1e-06 
0.0 1.0222 0 2.0 1e-06 
0.0 1.0223 0 2.0 1e-06 
0.0 1.0224 0 2.0 1e-06 
0.0 1.0225 0 2.0 1e-06 
0.0 1.0226 0 2.0 1e-06 
0.0 1.0227 0 2.0 1e-06 
0.0 1.0228 0 2.0 1e-06 
0.0 1.0229 0 2.0 1e-06 
0.0 1.023 0 2.0 1e-06 
0.0 1.0231 0 2.0 1e-06 
0.0 1.0232 0 2.0 1e-06 
0.0 1.0233 0 2.0 1e-06 
0.0 1.0234 0 2.0 1e-06 
0.0 1.0235 0 2.0 1e-06 
0.0 1.0236 0 2.0 1e-06 
0.0 1.0237 0 2.0 1e-06 
0.0 1.0238 0 2.0 1e-06 
0.0 1.0239 0 2.0 1e-06 
0.0 1.024 0 2.0 1e-06 
0.0 1.0241 0 2.0 1e-06 
0.0 1.0242 0 2.0 1e-06 
0.0 1.0243 0 2.0 1e-06 
0.0 1.0244 0 2.0 1e-06 
0.0 1.0245 0 2.0 1e-06 
0.0 1.0246 0 2.0 1e-06 
0.0 1.0247 0 2.0 1e-06 
0.0 1.0248 0 2.0 1e-06 
0.0 1.0249 0 2.0 1e-06 
0.0 1.025 0 2.0 1e-06 
0.0 1.0251 0 2.0 1e-06 
0.0 1.0252 0 2.0 1e-06 
0.0 1.0253 0 2.0 1e-06 
0.0 1.0254 0 2.0 1e-06 
0.0 1.0255 0 2.0 1e-06 
0.0 1.0256 0 2.0 1e-06 
0.0 1.0257 0 2.0 1e-06 
0.0 1.0258 0 2.0 1e-06 
0.0 1.0259 0 2.0 1e-06 
0.0 1.026 0 2.0 1e-06 
0.0 1.0261 0 2.0 1e-06 
0.0 1.0262 0 2.0 1e-06 
0.0 1.0263 0 2.0 1e-06 
0.0 1.0264 0 2.0 1e-06 
0.0 1.0265 0 2.0 1e-06 
0.0 1.0266 0 2.0 1e-06 
0.0 1.0267 0 2.0 1e-06 
0.0 1.0268 0 2.0 1e-06 
0.0 1.0269 0 2.0 1e-06 
0.0 1.027 0 2.0 1e-06 
0.0 1.0271 0 2.0 1e-06 
0.0 1.0272 0 2.0 1e-06 
0.0 1.0273 0 2.0 1e-06 
0.0 1.0274 0 2.0 1e-06 
0.0 1.0275 0 2.0 1e-06 
0.0 1.0276 0 2.0 1e-06 
0.0 1.0277 0 2.0 1e-06 
0.0 1.0278 0 2.0 1e-06 
0.0 1.0279 0 2.0 1e-06 
0.0 1.028 0 2.0 1e-06 
0.0 1.0281 0 2.0 1e-06 
0.0 1.0282 0 2.0 1e-06 
0.0 1.0283 0 2.0 1e-06 
0.0 1.0284 0 2.0 1e-06 
0.0 1.0285 0 2.0 1e-06 
0.0 1.0286 0 2.0 1e-06 
0.0 1.0287 0 2.0 1e-06 
0.0 1.0288 0 2.0 1e-06 
0.0 1.0289 0 2.0 1e-06 
0.0 1.029 0 2.0 1e-06 
0.0 1.0291 0 2.0 1e-06 
0.0 1.0292 0 2.0 1e-06 
0.0 1.0293 0 2.0 1e-06 
0.0 1.0294 0 2.0 1e-06 
0.0 1.0295 0 2.0 1e-06 
0.0 1.0296 0 2.0 1e-06 
0.0 1.0297 0 2.0 1e-06 
0.0 1.0298 0 2.0 1e-06 
0.0 1.0299 0 2.0 1e-06 
0.0 1.03 0 2.0 1e-06 
0.0 1.0301 0 2.0 1e-06 
0.0 1.0302 0 2.0 1e-06 
0.0 1.0303 0 2.0 1e-06 
0.0 1.0304 0 2.0 1e-06 
0.0 1.0305 0 2.0 1e-06 
0.0 1.0306 0 2.0 1e-06 
0.0 1.0307 0 2.0 1e-06 
0.0 1.0308 0 2.0 1e-06 
0.0 1.0309 0 2.0 1e-06 
0.0 1.031 0 2.0 1e-06 
0.0 1.0311 0 2.0 1e-06 
0.0 1.0312 0 2.0 1e-06 
0.0 1.0313 0 2.0 1e-06 
0.0 1.0314 0 2.0 1e-06 
0.0 1.0315 0 2.0 1e-06 
0.0 1.0316 0 2.0 1e-06 
0.0 1.0317 0 2.0 1e-06 
0.0 1.0318 0 2.0 1e-06 
0.0 1.0319 0 2.0 1e-06 
0.0 1.032 0 2.0 1e-06 
0.0 1.0321 0 2.0 1e-06 
0.0 1.0322 0 2.0 1e-06 
0.0 1.0323 0 2.0 1e-06 
0.0 1.0324 0 2.0 1e-06 
0.0 1.0325 0 2.0 1e-06 
0.0 1.0326 0 2.0 1e-06 
0.0 1.0327 0 2.0 1e-06 
0.0 1.0328 0 2.0 1e-06 
0.0 1.0329 0 2.0 1e-06 
0.0 1.033 0 2.0 1e-06 
0.0 1.0331 0 2.0 1e-06 
0.0 1.0332 0 2.0 1e-06 
0.0 1.0333 0 2.0 1e-06 
0.0 1.0334 0 2.0 1e-06 
0.0 1.0335 0 2.0 1e-06 
0.0 1.0336 0 2.0 1e-06 
0.0 1.0337 0 2.0 1e-06 
0.0 1.0338 0 2.0 1e-06 
0.0 1.0339 0 2.0 1e-06 
0.0 1.034 0 2.0 1e-06 
0.0 1.0341 0 2.0 1e-06 
0.0 1.0342 0 2.0 1e-06 
0.0 1.0343 0 2.0 1e-06 
0.0 1.0344 0 2.0 1e-06 
0.0 1.0345 0 2.0 1e-06 
0.0 1.0346 0 2.0 1e-06 
0.0 1.0347 0 2.0 1e-06 
0.0 1.0348 0 2.0 1e-06 
0.0 1.0349 0 2.0 1e-06 
0.0 1.035 0 2.0 1e-06 
0.0 1.0351 0 2.0 1e-06 
0.0 1.0352 0 2.0 1e-06 
0.0 1.0353 0 2.0 1e-06 
0.0 1.0354 0 2.0 1e-06 
0.0 1.0355 0 2.0 1e-06 
0.0 1.0356 0 2.0 1e-06 
0.0 1.0357 0 2.0 1e-06 
0.0 1.0358 0 2.0 1e-06 
0.0 1.0359 0 2.0 1e-06 
0.0 1.036 0 2.0 1e-06 
0.0 1.0361 0 2.0 1e-06 
0.0 1.0362 0 2.0 1e-06 
0.0 1.0363 0 2.0 1e-06 
0.0 1.0364 0 2.0 1e-06 
0.0 1.0365 0 2.0 1e-06 
0.0 1.0366 0 2.0 1e-06 
0.0 1.0367 0 2.0 1e-06 
0.0 1.0368 0 2.0 1e-06 
0.0 1.0369 0 2.0 1e-06 
0.0 1.037 0 2.0 1e-06 
0.0 1.0371 0 2.0 1e-06 
0.0 1.0372 0 2.0 1e-06 
0.0 1.0373 0 2.0 1e-06 
0.0 1.0374 0 2.0 1e-06 
0.0 1.0375 0 2.0 1e-06 
0.0 1.0376 0 2.0 1e-06 
0.0 1.0377 0 2.0 1e-06 
0.0 1.0378 0 2.0 1e-06 
0.0 1.0379 0 2.0 1e-06 
0.0 1.038 0 2.0 1e-06 
0.0 1.0381 0 2.0 1e-06 
0.0 1.0382 0 2.0 1e-06 
0.0 1.0383 0 2.0 1e-06 
0.0 1.0384 0 2.0 1e-06 
0.0 1.0385 0 2.0 1e-06 
0.0 1.0386 0 2.0 1e-06 
0.0 1.0387 0 2.0 1e-06 
0.0 1.0388 0 2.0 1e-06 
0.0 1.0389 0 2.0 1e-06 
0.0 1.039 0 2.0 1e-06 
0.0 1.0391 0 2.0 1e-06 
0.0 1.0392 0 2.0 1e-06 
0.0 1.0393 0 2.0 1e-06 
0.0 1.0394 0 2.0 1e-06 
0.0 1.0395 0 2.0 1e-06 
0.0 1.0396 0 2.0 1e-06 
0.0 1.0397 0 2.0 1e-06 
0.0 1.0398 0 2.0 1e-06 
0.0 1.0399 0 2.0 1e-06 
0.0 1.04 0 2.0 1e-06 
0.0 1.0401 0 2.0 1e-06 
0.0 1.0402 0 2.0 1e-06 
0.0 1.0403 0 2.0 1e-06 
0.0 1.0404 0 2.0 1e-06 
0.0 1.0405 0 2.0 1e-06 
0.0 1.0406 0 2.0 1e-06 
0.0 1.0407 0 2.0 1e-06 
0.0 1.0408 0 2.0 1e-06 
0.0 1.0409 0 2.0 1e-06 
0.0 1.041 0 2.0 1e-06 
0.0 1.0411 0 2.0 1e-06 
0.0 1.0412 0 2.0 1e-06 
0.0 1.0413 0 2.0 1e-06 
0.0 1.0414 0 2.0 1e-06 
0.0 1.0415 0 2.0 1e-06 
0.0 1.0416 0 2.0 1e-06 
0.0 1.0417 0 2.0 1e-06 
0.0 1.0418 0 2.0 1e-06 
0.0 1.0419 0 2.0 1e-06 
0.0 1.042 0 2.0 1e-06 
0.0 1.0421 0 2.0 1e-06 
0.0 1.0422 0 2.0 1e-06 
0.0 1.0423 0 2.0 1e-06 
0.0 1.0424 0 2.0 1e-06 
0.0 1.0425 0 2.0 1e-06 
0.0 1.0426 0 2.0 1e-06 
0.0 1.0427 0 2.0 1e-06 
0.0 1.0428 0 2.0 1e-06 
0.0 1.0429 0 2.0 1e-06 
0.0 1.043 0 2.0 1e-06 
0.0 1.0431 0 2.0 1e-06 
0.0 1.0432 0 2.0 1e-06 
0.0 1.0433 0 2.0 1e-06 
0.0 1.0434 0 2.0 1e-06 
0.0 1.0435 0 2.0 1e-06 
0.0 1.0436 0 2.0 1e-06 
0.0 1.0437 0 2.0 1e-06 
0.0 1.0438 0 2.0 1e-06 
0.0 1.0439 0 2.0 1e-06 
0.0 1.044 0 2.0 1e-06 
0.0 1.0441 0 2.0 1e-06 
0.0 1.0442 0 2.0 1e-06 
0.0 1.0443 0 2.0 1e-06 
0.0 1.0444 0 2.0 1e-06 
0.0 1.0445 0 2.0 1e-06 
0.0 1.0446 0 2.0 1e-06 
0.0 1.0447 0 2.0 1e-06 
0.0 1.0448 0 2.0 1e-06 
0.0 1.0449 0 2.0 1e-06 
0.0 1.045 0 2.0 1e-06 
0.0 1.0451 0 2.0 1e-06 
0.0 1.0452 0 2.0 1e-06 
0.0 1.0453 0 2.0 1e-06 
0.0 1.0454 0 2.0 1e-06 
0.0 1.0455 0 2.0 1e-06 
0.0 1.0456 0 2.0 1e-06 
0.0 1.0457 0 2.0 1e-06 
0.0 1.0458 0 2.0 1e-06 
0.0 1.0459 0 2.0 1e-06 
0.0 1.046 0 2.0 1e-06 
0.0 1.0461 0 2.0 1e-06 
0.0 1.0462 0 2.0 1e-06 
0.0 1.0463 0 2.0 1e-06 
0.0 1.0464 0 2.0 1e-06 
0.0 1.0465 0 2.0 1e-06 
0.0 1.0466 0 2.0 1e-06 
0.0 1.0467 0 2.0 1e-06 
0.0 1.0468 0 2.0 1e-06 
0.0 1.0469 0 2.0 1e-06 
0.0 1.047 0 2.0 1e-06 
0.0 1.0471 0 2.0 1e-06 
0.0 1.0472 0 2.0 1e-06 
0.0 1.0473 0 2.0 1e-06 
0.0 1.0474 0 2.0 1e-06 
0.0 1.0475 0 2.0 1e-06 
0.0 1.0476 0 2.0 1e-06 
0.0 1.0477 0 2.0 1e-06 
0.0 1.0478 0 2.0 1e-06 
0.0 1.0479 0 2.0 1e-06 
0.0 1.048 0 2.0 1e-06 
0.0 1.0481 0 2.0 1e-06 
0.0 1.0482 0 2.0 1e-06 
0.0 1.0483 0 2.0 1e-06 
0.0 1.0484 0 2.0 1e-06 
0.0 1.0485 0 2.0 1e-06 
0.0 1.0486 0 2.0 1e-06 
0.0 1.0487 0 2.0 1e-06 
0.0 1.0488 0 2.0 1e-06 
0.0 1.0489 0 2.0 1e-06 
0.0 1.049 0 2.0 1e-06 
0.0 1.0491 0 2.0 1e-06 
0.0 1.0492 0 2.0 1e-06 
0.0 1.0493 0 2.0 1e-06 
0.0 1.0494 0 2.0 1e-06 
0.0 1.0495 0 2.0 1e-06 
0.0 1.0496 0 2.0 1e-06 
0.0 1.0497 0 2.0 1e-06 
0.0 1.0498 0 2.0 1e-06 
0.0 1.0499 0 2.0 1e-06 
0.0 1.05 0 2.0 1e-06 
0.0 1.0501 0 2.0 1e-06 
0.0 1.0502 0 2.0 1e-06 
0.0 1.0503 0 2.0 1e-06 
0.0 1.0504 0 2.0 1e-06 
0.0 1.0505 0 2.0 1e-06 
0.0 1.0506 0 2.0 1e-06 
0.0 1.0507 0 2.0 1e-06 
0.0 1.0508 0 2.0 1e-06 
0.0 1.0509 0 2.0 1e-06 
0.0 1.051 0 2.0 1e-06 
0.0 1.0511 0 2.0 1e-06 
0.0 1.0512 0 2.0 1e-06 
0.0 1.0513 0 2.0 1e-06 
0.0 1.0514 0 2.0 1e-06 
0.0 1.0515 0 2.0 1e-06 
0.0 1.0516 0 2.0 1e-06 
0.0 1.0517 0 2.0 1e-06 
0.0 1.0518 0 2.0 1e-06 
0.0 1.0519 0 2.0 1e-06 
0.0 1.052 0 2.0 1e-06 
0.0 1.0521 0 2.0 1e-06 
0.0 1.0522 0 2.0 1e-06 
0.0 1.0523 0 2.0 1e-06 
0.0 1.0524 0 2.0 1e-06 
0.0 1.0525 0 2.0 1e-06 
0.0 1.0526 0 2.0 1e-06 
0.0 1.0527 0 2.0 1e-06 
0.0 1.0528 0 2.0 1e-06 
0.0 1.0529 0 2.0 1e-06 
0.0 1.053 0 2.0 1e-06 
0.0 1.0531 0 2.0 1e-06 
0.0 1.0532 0 2.0 1e-06 
0.0 1.0533 0 2.0 1e-06 
0.0 1.0534 0 2.0 1e-06 
0.0 1.0535 0 2.0 1e-06 
0.0 1.0536 0 2.0 1e-06 
0.0 1.0537 0 2.0 1e-06 
0.0 1.0538 0 2.0 1e-06 
0.0 1.0539 0 2.0 1e-06 
0.0 1.054 0 2.0 1e-06 
0.0 1.0541 0 2.0 1e-06 
0.0 1.0542 0 2.0 1e-06 
0.0 1.0543 0 2.0 1e-06 
0.0 1.0544 0 2.0 1e-06 
0.0 1.0545 0 2.0 1e-06 
0.0 1.0546 0 2.0 1e-06 
0.0 1.0547 0 2.0 1e-06 
0.0 1.0548 0 2.0 1e-06 
0.0 1.0549 0 2.0 1e-06 
0.0 1.055 0 2.0 1e-06 
0.0 1.0551 0 2.0 1e-06 
0.0 1.0552 0 2.0 1e-06 
0.0 1.0553 0 2.0 1e-06 
0.0 1.0554 0 2.0 1e-06 
0.0 1.0555 0 2.0 1e-06 
0.0 1.0556 0 2.0 1e-06 
0.0 1.0557 0 2.0 1e-06 
0.0 1.0558 0 2.0 1e-06 
0.0 1.0559 0 2.0 1e-06 
0.0 1.056 0 2.0 1e-06 
0.0 1.0561 0 2.0 1e-06 
0.0 1.0562 0 2.0 1e-06 
0.0 1.0563 0 2.0 1e-06 
0.0 1.0564 0 2.0 1e-06 
0.0 1.0565 0 2.0 1e-06 
0.0 1.0566 0 2.0 1e-06 
0.0 1.0567 0 2.0 1e-06 
0.0 1.0568 0 2.0 1e-06 
0.0 1.0569 0 2.0 1e-06 
0.0 1.057 0 2.0 1e-06 
0.0 1.0571 0 2.0 1e-06 
0.0 1.0572 0 2.0 1e-06 
0.0 1.0573 0 2.0 1e-06 
0.0 1.0574 0 2.0 1e-06 
0.0 1.0575 0 2.0 1e-06 
0.0 1.0576 0 2.0 1e-06 
0.0 1.0577 0 2.0 1e-06 
0.0 1.0578 0 2.0 1e-06 
0.0 1.0579 0 2.0 1e-06 
0.0 1.058 0 2.0 1e-06 
0.0 1.0581 0 2.0 1e-06 
0.0 1.0582 0 2.0 1e-06 
0.0 1.0583 0 2.0 1e-06 
0.0 1.0584 0 2.0 1e-06 
0.0 1.0585 0 2.0 1e-06 
0.0 1.0586 0 2.0 1e-06 
0.0 1.0587 0 2.0 1e-06 
0.0 1.0588 0 2.0 1e-06 
0.0 1.0589 0 2.0 1e-06 
0.0 1.059 0 2.0 1e-06 
0.0 1.0591 0 2.0 1e-06 
0.0 1.0592 0 2.0 1e-06 
0.0 1.0593 0 2.0 1e-06 
0.0 1.0594 0 2.0 1e-06 
0.0 1.0595 0 2.0 1e-06 
0.0 1.0596 0 2.0 1e-06 
0.0 1.0597 0 2.0 1e-06 
0.0 1.0598 0 2.0 1e-06 
0.0 1.0599 0 2.0 1e-06 
0.0 1.06 0 2.0 1e-06 
0.0 1.0601 0 2.0 1e-06 
0.0 1.0602 0 2.0 1e-06 
0.0 1.0603 0 2.0 1e-06 
0.0 1.0604 0 2.0 1e-06 
0.0 1.0605 0 2.0 1e-06 
0.0 1.0606 0 2.0 1e-06 
0.0 1.0607 0 2.0 1e-06 
0.0 1.0608 0 2.0 1e-06 
0.0 1.0609 0 2.0 1e-06 
0.0 1.061 0 2.0 1e-06 
0.0 1.0611 0 2.0 1e-06 
0.0 1.0612 0 2.0 1e-06 
0.0 1.0613 0 2.0 1e-06 
0.0 1.0614 0 2.0 1e-06 
0.0 1.0615 0 2.0 1e-06 
0.0 1.0616 0 2.0 1e-06 
0.0 1.0617 0 2.0 1e-06 
0.0 1.0618 0 2.0 1e-06 
0.0 1.0619 0 2.0 1e-06 
0.0 1.062 0 2.0 1e-06 
0.0 1.0621 0 2.0 1e-06 
0.0 1.0622 0 2.0 1e-06 
0.0 1.0623 0 2.0 1e-06 
0.0 1.0624 0 2.0 1e-06 
0.0 1.0625 0 2.0 1e-06 
0.0 1.0626 0 2.0 1e-06 
0.0 1.0627 0 2.0 1e-06 
0.0 1.0628 0 2.0 1e-06 
0.0 1.0629 0 2.0 1e-06 
0.0 1.063 0 2.0 1e-06 
0.0 1.0631 0 2.0 1e-06 
0.0 1.0632 0 2.0 1e-06 
0.0 1.0633 0 2.0 1e-06 
0.0 1.0634 0 2.0 1e-06 
0.0 1.0635 0 2.0 1e-06 
0.0 1.0636 0 2.0 1e-06 
0.0 1.0637 0 2.0 1e-06 
0.0 1.0638 0 2.0 1e-06 
0.0 1.0639 0 2.0 1e-06 
0.0 1.064 0 2.0 1e-06 
0.0 1.0641 0 2.0 1e-06 
0.0 1.0642 0 2.0 1e-06 
0.0 1.0643 0 2.0 1e-06 
0.0 1.0644 0 2.0 1e-06 
0.0 1.0645 0 2.0 1e-06 
0.0 1.0646 0 2.0 1e-06 
0.0 1.0647 0 2.0 1e-06 
0.0 1.0648 0 2.0 1e-06 
0.0 1.0649 0 2.0 1e-06 
0.0 1.065 0 2.0 1e-06 
0.0 1.0651 0 2.0 1e-06 
0.0 1.0652 0 2.0 1e-06 
0.0 1.0653 0 2.0 1e-06 
0.0 1.0654 0 2.0 1e-06 
0.0 1.0655 0 2.0 1e-06 
0.0 1.0656 0 2.0 1e-06 
0.0 1.0657 0 2.0 1e-06 
0.0 1.0658 0 2.0 1e-06 
0.0 1.0659 0 2.0 1e-06 
0.0 1.066 0 2.0 1e-06 
0.0 1.0661 0 2.0 1e-06 
0.0 1.0662 0 2.0 1e-06 
0.0 1.0663 0 2.0 1e-06 
0.0 1.0664 0 2.0 1e-06 
0.0 1.0665 0 2.0 1e-06 
0.0 1.0666 0 2.0 1e-06 
0.0 1.0667 0 2.0 1e-06 
0.0 1.0668 0 2.0 1e-06 
0.0 1.0669 0 2.0 1e-06 
0.0 1.067 0 2.0 1e-06 
0.0 1.0671 0 2.0 1e-06 
0.0 1.0672 0 2.0 1e-06 
0.0 1.0673 0 2.0 1e-06 
0.0 1.0674 0 2.0 1e-06 
0.0 1.0675 0 2.0 1e-06 
0.0 1.0676 0 2.0 1e-06 
0.0 1.0677 0 2.0 1e-06 
0.0 1.0678 0 2.0 1e-06 
0.0 1.0679 0 2.0 1e-06 
0.0 1.068 0 2.0 1e-06 
0.0 1.0681 0 2.0 1e-06 
0.0 1.0682 0 2.0 1e-06 
0.0 1.0683 0 2.0 1e-06 
0.0 1.0684 0 2.0 1e-06 
0.0 1.0685 0 2.0 1e-06 
0.0 1.0686 0 2.0 1e-06 
0.0 1.0687 0 2.0 1e-06 
0.0 1.0688 0 2.0 1e-06 
0.0 1.0689 0 2.0 1e-06 
0.0 1.069 0 2.0 1e-06 
0.0 1.0691 0 2.0 1e-06 
0.0 1.0692 0 2.0 1e-06 
0.0 1.0693 0 2.0 1e-06 
0.0 1.0694 0 2.0 1e-06 
0.0 1.0695 0 2.0 1e-06 
0.0 1.0696 0 2.0 1e-06 
0.0 1.0697 0 2.0 1e-06 
0.0 1.0698 0 2.0 1e-06 
0.0 1.0699 0 2.0 1e-06 
0.0 1.07 0 2.0 1e-06 
0.0 1.0701 0 2.0 1e-06 
0.0 1.0702 0 2.0 1e-06 
0.0 1.0703 0 2.0 1e-06 
0.0 1.0704 0 2.0 1e-06 
0.0 1.0705 0 2.0 1e-06 
0.0 1.0706 0 2.0 1e-06 
0.0 1.0707 0 2.0 1e-06 
0.0 1.0708 0 2.0 1e-06 
0.0 1.0709 0 2.0 1e-06 
0.0 1.071 0 2.0 1e-06 
0.0 1.0711 0 2.0 1e-06 
0.0 1.0712 0 2.0 1e-06 
0.0 1.0713 0 2.0 1e-06 
0.0 1.0714 0 2.0 1e-06 
0.0 1.0715 0 2.0 1e-06 
0.0 1.0716 0 2.0 1e-06 
0.0 1.0717 0 2.0 1e-06 
0.0 1.0718 0 2.0 1e-06 
0.0 1.0719 0 2.0 1e-06 
0.0 1.072 0 2.0 1e-06 
0.0 1.0721 0 2.0 1e-06 
0.0 1.0722 0 2.0 1e-06 
0.0 1.0723 0 2.0 1e-06 
0.0 1.0724 0 2.0 1e-06 
0.0 1.0725 0 2.0 1e-06 
0.0 1.0726 0 2.0 1e-06 
0.0 1.0727 0 2.0 1e-06 
0.0 1.0728 0 2.0 1e-06 
0.0 1.0729 0 2.0 1e-06 
0.0 1.073 0 2.0 1e-06 
0.0 1.0731 0 2.0 1e-06 
0.0 1.0732 0 2.0 1e-06 
0.0 1.0733 0 2.0 1e-06 
0.0 1.0734 0 2.0 1e-06 
0.0 1.0735 0 2.0 1e-06 
0.0 1.0736 0 2.0 1e-06 
0.0 1.0737 0 2.0 1e-06 
0.0 1.0738 0 2.0 1e-06 
0.0 1.0739 0 2.0 1e-06 
0.0 1.074 0 2.0 1e-06 
0.0 1.0741 0 2.0 1e-06 
0.0 1.0742 0 2.0 1e-06 
0.0 1.0743 0 2.0 1e-06 
0.0 1.0744 0 2.0 1e-06 
0.0 1.0745 0 2.0 1e-06 
0.0 1.0746 0 2.0 1e-06 
0.0 1.0747 0 2.0 1e-06 
0.0 1.0748 0 2.0 1e-06 
0.0 1.0749 0 2.0 1e-06 
0.0 1.075 0 2.0 1e-06 
0.0 1.0751 0 2.0 1e-06 
0.0 1.0752 0 2.0 1e-06 
0.0 1.0753 0 2.0 1e-06 
0.0 1.0754 0 2.0 1e-06 
0.0 1.0755 0 2.0 1e-06 
0.0 1.0756 0 2.0 1e-06 
0.0 1.0757 0 2.0 1e-06 
0.0 1.0758 0 2.0 1e-06 
0.0 1.0759 0 2.0 1e-06 
0.0 1.076 0 2.0 1e-06 
0.0 1.0761 0 2.0 1e-06 
0.0 1.0762 0 2.0 1e-06 
0.0 1.0763 0 2.0 1e-06 
0.0 1.0764 0 2.0 1e-06 
0.0 1.0765 0 2.0 1e-06 
0.0 1.0766 0 2.0 1e-06 
0.0 1.0767 0 2.0 1e-06 
0.0 1.0768 0 2.0 1e-06 
0.0 1.0769 0 2.0 1e-06 
0.0 1.077 0 2.0 1e-06 
0.0 1.0771 0 2.0 1e-06 
0.0 1.0772 0 2.0 1e-06 
0.0 1.0773 0 2.0 1e-06 
0.0 1.0774 0 2.0 1e-06 
0.0 1.0775 0 2.0 1e-06 
0.0 1.0776 0 2.0 1e-06 
0.0 1.0777 0 2.0 1e-06 
0.0 1.0778 0 2.0 1e-06 
0.0 1.0779 0 2.0 1e-06 
0.0 1.078 0 2.0 1e-06 
0.0 1.0781 0 2.0 1e-06 
0.0 1.0782 0 2.0 1e-06 
0.0 1.0783 0 2.0 1e-06 
0.0 1.0784 0 2.0 1e-06 
0.0 1.0785 0 2.0 1e-06 
0.0 1.0786 0 2.0 1e-06 
0.0 1.0787 0 2.0 1e-06 
0.0 1.0788 0 2.0 1e-06 
0.0 1.0789 0 2.0 1e-06 
0.0 1.079 0 2.0 1e-06 
0.0 1.0791 0 2.0 1e-06 
0.0 1.0792 0 2.0 1e-06 
0.0 1.0793 0 2.0 1e-06 
0.0 1.0794 0 2.0 1e-06 
0.0 1.0795 0 2.0 1e-06 
0.0 1.0796 0 2.0 1e-06 
0.0 1.0797 0 2.0 1e-06 
0.0 1.0798 0 2.0 1e-06 
0.0 1.0799 0 2.0 1e-06 
0.0 1.08 0 2.0 1e-06 
0.0 1.0801 0 2.0 1e-06 
0.0 1.0802 0 2.0 1e-06 
0.0 1.0803 0 2.0 1e-06 
0.0 1.0804 0 2.0 1e-06 
0.0 1.0805 0 2.0 1e-06 
0.0 1.0806 0 2.0 1e-06 
0.0 1.0807 0 2.0 1e-06 
0.0 1.0808 0 2.0 1e-06 
0.0 1.0809 0 2.0 1e-06 
0.0 1.081 0 2.0 1e-06 
0.0 1.0811 0 2.0 1e-06 
0.0 1.0812 0 2.0 1e-06 
0.0 1.0813 0 2.0 1e-06 
0.0 1.0814 0 2.0 1e-06 
0.0 1.0815 0 2.0 1e-06 
0.0 1.0816 0 2.0 1e-06 
0.0 1.0817 0 2.0 1e-06 
0.0 1.0818 0 2.0 1e-06 
0.0 1.0819 0 2.0 1e-06 
0.0 1.082 0 2.0 1e-06 
0.0 1.0821 0 2.0 1e-06 
0.0 1.0822 0 2.0 1e-06 
0.0 1.0823 0 2.0 1e-06 
0.0 1.0824 0 2.0 1e-06 
0.0 1.0825 0 2.0 1e-06 
0.0 1.0826 0 2.0 1e-06 
0.0 1.0827 0 2.0 1e-06 
0.0 1.0828 0 2.0 1e-06 
0.0 1.0829 0 2.0 1e-06 
0.0 1.083 0 2.0 1e-06 
0.0 1.0831 0 2.0 1e-06 
0.0 1.0832 0 2.0 1e-06 
0.0 1.0833 0 2.0 1e-06 
0.0 1.0834 0 2.0 1e-06 
0.0 1.0835 0 2.0 1e-06 
0.0 1.0836 0 2.0 1e-06 
0.0 1.0837 0 2.0 1e-06 
0.0 1.0838 0 2.0 1e-06 
0.0 1.0839 0 2.0 1e-06 
0.0 1.084 0 2.0 1e-06 
0.0 1.0841 0 2.0 1e-06 
0.0 1.0842 0 2.0 1e-06 
0.0 1.0843 0 2.0 1e-06 
0.0 1.0844 0 2.0 1e-06 
0.0 1.0845 0 2.0 1e-06 
0.0 1.0846 0 2.0 1e-06 
0.0 1.0847 0 2.0 1e-06 
0.0 1.0848 0 2.0 1e-06 
0.0 1.0849 0 2.0 1e-06 
0.0 1.085 0 2.0 1e-06 
0.0 1.0851 0 2.0 1e-06 
0.0 1.0852 0 2.0 1e-06 
0.0 1.0853 0 2.0 1e-06 
0.0 1.0854 0 2.0 1e-06 
0.0 1.0855 0 2.0 1e-06 
0.0 1.0856 0 2.0 1e-06 
0.0 1.0857 0 2.0 1e-06 
0.0 1.0858 0 2.0 1e-06 
0.0 1.0859 0 2.0 1e-06 
0.0 1.086 0 2.0 1e-06 
0.0 1.0861 0 2.0 1e-06 
0.0 1.0862 0 2.0 1e-06 
0.0 1.0863 0 2.0 1e-06 
0.0 1.0864 0 2.0 1e-06 
0.0 1.0865 0 2.0 1e-06 
0.0 1.0866 0 2.0 1e-06 
0.0 1.0867 0 2.0 1e-06 
0.0 1.0868 0 2.0 1e-06 
0.0 1.0869 0 2.0 1e-06 
0.0 1.087 0 2.0 1e-06 
0.0 1.0871 0 2.0 1e-06 
0.0 1.0872 0 2.0 1e-06 
0.0 1.0873 0 2.0 1e-06 
0.0 1.0874 0 2.0 1e-06 
0.0 1.0875 0 2.0 1e-06 
0.0 1.0876 0 2.0 1e-06 
0.0 1.0877 0 2.0 1e-06 
0.0 1.0878 0 2.0 1e-06 
0.0 1.0879 0 2.0 1e-06 
0.0 1.088 0 2.0 1e-06 
0.0 1.0881 0 2.0 1e-06 
0.0 1.0882 0 2.0 1e-06 
0.0 1.0883 0 2.0 1e-06 
0.0 1.0884 0 2.0 1e-06 
0.0 1.0885 0 2.0 1e-06 
0.0 1.0886 0 2.0 1e-06 
0.0 1.0887 0 2.0 1e-06 
0.0 1.0888 0 2.0 1e-06 
0.0 1.0889 0 2.0 1e-06 
0.0 1.089 0 2.0 1e-06 
0.0 1.0891 0 2.0 1e-06 
0.0 1.0892 0 2.0 1e-06 
0.0 1.0893 0 2.0 1e-06 
0.0 1.0894 0 2.0 1e-06 
0.0 1.0895 0 2.0 1e-06 
0.0 1.0896 0 2.0 1e-06 
0.0 1.0897 0 2.0 1e-06 
0.0 1.0898 0 2.0 1e-06 
0.0 1.0899 0 2.0 1e-06 
0.0 1.09 0 2.0 1e-06 
0.0 1.0901 0 2.0 1e-06 
0.0 1.0902 0 2.0 1e-06 
0.0 1.0903 0 2.0 1e-06 
0.0 1.0904 0 2.0 1e-06 
0.0 1.0905 0 2.0 1e-06 
0.0 1.0906 0 2.0 1e-06 
0.0 1.0907 0 2.0 1e-06 
0.0 1.0908 0 2.0 1e-06 
0.0 1.0909 0 2.0 1e-06 
0.0 1.091 0 2.0 1e-06 
0.0 1.0911 0 2.0 1e-06 
0.0 1.0912 0 2.0 1e-06 
0.0 1.0913 0 2.0 1e-06 
0.0 1.0914 0 2.0 1e-06 
0.0 1.0915 0 2.0 1e-06 
0.0 1.0916 0 2.0 1e-06 
0.0 1.0917 0 2.0 1e-06 
0.0 1.0918 0 2.0 1e-06 
0.0 1.0919 0 2.0 1e-06 
0.0 1.092 0 2.0 1e-06 
0.0 1.0921 0 2.0 1e-06 
0.0 1.0922 0 2.0 1e-06 
0.0 1.0923 0 2.0 1e-06 
0.0 1.0924 0 2.0 1e-06 
0.0 1.0925 0 2.0 1e-06 
0.0 1.0926 0 2.0 1e-06 
0.0 1.0927 0 2.0 1e-06 
0.0 1.0928 0 2.0 1e-06 
0.0 1.0929 0 2.0 1e-06 
0.0 1.093 0 2.0 1e-06 
0.0 1.0931 0 2.0 1e-06 
0.0 1.0932 0 2.0 1e-06 
0.0 1.0933 0 2.0 1e-06 
0.0 1.0934 0 2.0 1e-06 
0.0 1.0935 0 2.0 1e-06 
0.0 1.0936 0 2.0 1e-06 
0.0 1.0937 0 2.0 1e-06 
0.0 1.0938 0 2.0 1e-06 
0.0 1.0939 0 2.0 1e-06 
0.0 1.094 0 2.0 1e-06 
0.0 1.0941 0 2.0 1e-06 
0.0 1.0942 0 2.0 1e-06 
0.0 1.0943 0 2.0 1e-06 
0.0 1.0944 0 2.0 1e-06 
0.0 1.0945 0 2.0 1e-06 
0.0 1.0946 0 2.0 1e-06 
0.0 1.0947 0 2.0 1e-06 
0.0 1.0948 0 2.0 1e-06 
0.0 1.0949 0 2.0 1e-06 
0.0 1.095 0 2.0 1e-06 
0.0 1.0951 0 2.0 1e-06 
0.0 1.0952 0 2.0 1e-06 
0.0 1.0953 0 2.0 1e-06 
0.0 1.0954 0 2.0 1e-06 
0.0 1.0955 0 2.0 1e-06 
0.0 1.0956 0 2.0 1e-06 
0.0 1.0957 0 2.0 1e-06 
0.0 1.0958 0 2.0 1e-06 
0.0 1.0959 0 2.0 1e-06 
0.0 1.096 0 2.0 1e-06 
0.0 1.0961 0 2.0 1e-06 
0.0 1.0962 0 2.0 1e-06 
0.0 1.0963 0 2.0 1e-06 
0.0 1.0964 0 2.0 1e-06 
0.0 1.0965 0 2.0 1e-06 
0.0 1.0966 0 2.0 1e-06 
0.0 1.0967 0 2.0 1e-06 
0.0 1.0968 0 2.0 1e-06 
0.0 1.0969 0 2.0 1e-06 
0.0 1.097 0 2.0 1e-06 
0.0 1.0971 0 2.0 1e-06 
0.0 1.0972 0 2.0 1e-06 
0.0 1.0973 0 2.0 1e-06 
0.0 1.0974 0 2.0 1e-06 
0.0 1.0975 0 2.0 1e-06 
0.0 1.0976 0 2.0 1e-06 
0.0 1.0977 0 2.0 1e-06 
0.0 1.0978 0 2.0 1e-06 
0.0 1.0979 0 2.0 1e-06 
0.0 1.098 0 2.0 1e-06 
0.0 1.0981 0 2.0 1e-06 
0.0 1.0982 0 2.0 1e-06 
0.0 1.0983 0 2.0 1e-06 
0.0 1.0984 0 2.0 1e-06 
0.0 1.0985 0 2.0 1e-06 
0.0 1.0986 0 2.0 1e-06 
0.0 1.0987 0 2.0 1e-06 
0.0 1.0988 0 2.0 1e-06 
0.0 1.0989 0 2.0 1e-06 
0.0 1.099 0 2.0 1e-06 
0.0 1.0991 0 2.0 1e-06 
0.0 1.0992 0 2.0 1e-06 
0.0 1.0993 0 2.0 1e-06 
0.0 1.0994 0 2.0 1e-06 
0.0 1.0995 0 2.0 1e-06 
0.0 1.0996 0 2.0 1e-06 
0.0 1.0997 0 2.0 1e-06 
0.0 1.0998 0 2.0 1e-06 
0.0 1.0999 0 2.0 1e-06 
0.0 1.1 0 2.0 1e-06 
0.0 1.1001 0 2.0 1e-06 
0.0 1.1002 0 2.0 1e-06 
0.0 1.1003 0 2.0 1e-06 
0.0 1.1004 0 2.0 1e-06 
0.0 1.1005 0 2.0 1e-06 
0.0 1.1006 0 2.0 1e-06 
0.0 1.1007 0 2.0 1e-06 
0.0 1.1008 0 2.0 1e-06 
0.0 1.1009 0 2.0 1e-06 
0.0 1.101 0 2.0 1e-06 
0.0 1.1011 0 2.0 1e-06 
0.0 1.1012 0 2.0 1e-06 
0.0 1.1013 0 2.0 1e-06 
0.0 1.1014 0 2.0 1e-06 
0.0 1.1015 0 2.0 1e-06 
0.0 1.1016 0 2.0 1e-06 
0.0 1.1017 0 2.0 1e-06 
0.0 1.1018 0 2.0 1e-06 
0.0 1.1019 0 2.0 1e-06 
0.0 1.102 0 2.0 1e-06 
0.0 1.1021 0 2.0 1e-06 
0.0 1.1022 0 2.0 1e-06 
0.0 1.1023 0 2.0 1e-06 
0.0 1.1024 0 2.0 1e-06 
0.0 1.1025 0 2.0 1e-06 
0.0 1.1026 0 2.0 1e-06 
0.0 1.1027 0 2.0 1e-06 
0.0 1.1028 0 2.0 1e-06 
0.0 1.1029 0 2.0 1e-06 
0.0 1.103 0 2.0 1e-06 
0.0 1.1031 0 2.0 1e-06 
0.0 1.1032 0 2.0 1e-06 
0.0 1.1033 0 2.0 1e-06 
0.0 1.1034 0 2.0 1e-06 
0.0 1.1035 0 2.0 1e-06 
0.0 1.1036 0 2.0 1e-06 
0.0 1.1037 0 2.0 1e-06 
0.0 1.1038 0 2.0 1e-06 
0.0 1.1039 0 2.0 1e-06 
0.0 1.104 0 2.0 1e-06 
0.0 1.1041 0 2.0 1e-06 
0.0 1.1042 0 2.0 1e-06 
0.0 1.1043 0 2.0 1e-06 
0.0 1.1044 0 2.0 1e-06 
0.0 1.1045 0 2.0 1e-06 
0.0 1.1046 0 2.0 1e-06 
0.0 1.1047 0 2.0 1e-06 
0.0 1.1048 0 2.0 1e-06 
0.0 1.1049 0 2.0 1e-06 
0.0 1.105 0 2.0 1e-06 
0.0 1.1051 0 2.0 1e-06 
0.0 1.1052 0 2.0 1e-06 
0.0 1.1053 0 2.0 1e-06 
0.0 1.1054 0 2.0 1e-06 
0.0 1.1055 0 2.0 1e-06 
0.0 1.1056 0 2.0 1e-06 
0.0 1.1057 0 2.0 1e-06 
0.0 1.1058 0 2.0 1e-06 
0.0 1.1059 0 2.0 1e-06 
0.0 1.106 0 2.0 1e-06 
0.0 1.1061 0 2.0 1e-06 
0.0 1.1062 0 2.0 1e-06 
0.0 1.1063 0 2.0 1e-06 
0.0 1.1064 0 2.0 1e-06 
0.0 1.1065 0 2.0 1e-06 
0.0 1.1066 0 2.0 1e-06 
0.0 1.1067 0 2.0 1e-06 
0.0 1.1068 0 2.0 1e-06 
0.0 1.1069 0 2.0 1e-06 
0.0 1.107 0 2.0 1e-06 
0.0 1.1071 0 2.0 1e-06 
0.0 1.1072 0 2.0 1e-06 
0.0 1.1073 0 2.0 1e-06 
0.0 1.1074 0 2.0 1e-06 
0.0 1.1075 0 2.0 1e-06 
0.0 1.1076 0 2.0 1e-06 
0.0 1.1077 0 2.0 1e-06 
0.0 1.1078 0 2.0 1e-06 
0.0 1.1079 0 2.0 1e-06 
0.0 1.108 0 2.0 1e-06 
0.0 1.1081 0 2.0 1e-06 
0.0 1.1082 0 2.0 1e-06 
0.0 1.1083 0 2.0 1e-06 
0.0 1.1084 0 2.0 1e-06 
0.0 1.1085 0 2.0 1e-06 
0.0 1.1086 0 2.0 1e-06 
0.0 1.1087 0 2.0 1e-06 
0.0 1.1088 0 2.0 1e-06 
0.0 1.1089 0 2.0 1e-06 
0.0 1.109 0 2.0 1e-06 
0.0 1.1091 0 2.0 1e-06 
0.0 1.1092 0 2.0 1e-06 
0.0 1.1093 0 2.0 1e-06 
0.0 1.1094 0 2.0 1e-06 
0.0 1.1095 0 2.0 1e-06 
0.0 1.1096 0 2.0 1e-06 
0.0 1.1097 0 2.0 1e-06 
0.0 1.1098 0 2.0 1e-06 
0.0 1.1099 0 2.0 1e-06 
0.0 1.11 0 2.0 1e-06 
0.0 1.1101 0 2.0 1e-06 
0.0 1.1102 0 2.0 1e-06 
0.0 1.1103 0 2.0 1e-06 
0.0 1.1104 0 2.0 1e-06 
0.0 1.1105 0 2.0 1e-06 
0.0 1.1106 0 2.0 1e-06 
0.0 1.1107 0 2.0 1e-06 
0.0 1.1108 0 2.0 1e-06 
0.0 1.1109 0 2.0 1e-06 
0.0 1.111 0 2.0 1e-06 
0.0 1.1111 0 2.0 1e-06 
0.0 1.1112 0 2.0 1e-06 
0.0 1.1113 0 2.0 1e-06 
0.0 1.1114 0 2.0 1e-06 
0.0 1.1115 0 2.0 1e-06 
0.0 1.1116 0 2.0 1e-06 
0.0 1.1117 0 2.0 1e-06 
0.0 1.1118 0 2.0 1e-06 
0.0 1.1119 0 2.0 1e-06 
0.0 1.112 0 2.0 1e-06 
0.0 1.1121 0 2.0 1e-06 
0.0 1.1122 0 2.0 1e-06 
0.0 1.1123 0 2.0 1e-06 
0.0 1.1124 0 2.0 1e-06 
0.0 1.1125 0 2.0 1e-06 
0.0 1.1126 0 2.0 1e-06 
0.0 1.1127 0 2.0 1e-06 
0.0 1.1128 0 2.0 1e-06 
0.0 1.1129 0 2.0 1e-06 
0.0 1.113 0 2.0 1e-06 
0.0 1.1131 0 2.0 1e-06 
0.0 1.1132 0 2.0 1e-06 
0.0 1.1133 0 2.0 1e-06 
0.0 1.1134 0 2.0 1e-06 
0.0 1.1135 0 2.0 1e-06 
0.0 1.1136 0 2.0 1e-06 
0.0 1.1137 0 2.0 1e-06 
0.0 1.1138 0 2.0 1e-06 
0.0 1.1139 0 2.0 1e-06 
0.0 1.114 0 2.0 1e-06 
0.0 1.1141 0 2.0 1e-06 
0.0 1.1142 0 2.0 1e-06 
0.0 1.1143 0 2.0 1e-06 
0.0 1.1144 0 2.0 1e-06 
0.0 1.1145 0 2.0 1e-06 
0.0 1.1146 0 2.0 1e-06 
0.0 1.1147 0 2.0 1e-06 
0.0 1.1148 0 2.0 1e-06 
0.0 1.1149 0 2.0 1e-06 
0.0 1.115 0 2.0 1e-06 
0.0 1.1151 0 2.0 1e-06 
0.0 1.1152 0 2.0 1e-06 
0.0 1.1153 0 2.0 1e-06 
0.0 1.1154 0 2.0 1e-06 
0.0 1.1155 0 2.0 1e-06 
0.0 1.1156 0 2.0 1e-06 
0.0 1.1157 0 2.0 1e-06 
0.0 1.1158 0 2.0 1e-06 
0.0 1.1159 0 2.0 1e-06 
0.0 1.116 0 2.0 1e-06 
0.0 1.1161 0 2.0 1e-06 
0.0 1.1162 0 2.0 1e-06 
0.0 1.1163 0 2.0 1e-06 
0.0 1.1164 0 2.0 1e-06 
0.0 1.1165 0 2.0 1e-06 
0.0 1.1166 0 2.0 1e-06 
0.0 1.1167 0 2.0 1e-06 
0.0 1.1168 0 2.0 1e-06 
0.0 1.1169 0 2.0 1e-06 
0.0 1.117 0 2.0 1e-06 
0.0 1.1171 0 2.0 1e-06 
0.0 1.1172 0 2.0 1e-06 
0.0 1.1173 0 2.0 1e-06 
0.0 1.1174 0 2.0 1e-06 
0.0 1.1175 0 2.0 1e-06 
0.0 1.1176 0 2.0 1e-06 
0.0 1.1177 0 2.0 1e-06 
0.0 1.1178 0 2.0 1e-06 
0.0 1.1179 0 2.0 1e-06 
0.0 1.118 0 2.0 1e-06 
0.0 1.1181 0 2.0 1e-06 
0.0 1.1182 0 2.0 1e-06 
0.0 1.1183 0 2.0 1e-06 
0.0 1.1184 0 2.0 1e-06 
0.0 1.1185 0 2.0 1e-06 
0.0 1.1186 0 2.0 1e-06 
0.0 1.1187 0 2.0 1e-06 
0.0 1.1188 0 2.0 1e-06 
0.0 1.1189 0 2.0 1e-06 
0.0 1.119 0 2.0 1e-06 
0.0 1.1191 0 2.0 1e-06 
0.0 1.1192 0 2.0 1e-06 
0.0 1.1193 0 2.0 1e-06 
0.0 1.1194 0 2.0 1e-06 
0.0 1.1195 0 2.0 1e-06 
0.0 1.1196 0 2.0 1e-06 
0.0 1.1197 0 2.0 1e-06 
0.0 1.1198 0 2.0 1e-06 
0.0 1.1199 0 2.0 1e-06 
0.0 1.12 0 2.0 1e-06 
0.0 1.1201 0 2.0 1e-06 
0.0 1.1202 0 2.0 1e-06 
0.0 1.1203 0 2.0 1e-06 
0.0 1.1204 0 2.0 1e-06 
0.0 1.1205 0 2.0 1e-06 
0.0 1.1206 0 2.0 1e-06 
0.0 1.1207 0 2.0 1e-06 
0.0 1.1208 0 2.0 1e-06 
0.0 1.1209 0 2.0 1e-06 
0.0 1.121 0 2.0 1e-06 
0.0 1.1211 0 2.0 1e-06 
0.0 1.1212 0 2.0 1e-06 
0.0 1.1213 0 2.0 1e-06 
0.0 1.1214 0 2.0 1e-06 
0.0 1.1215 0 2.0 1e-06 
0.0 1.1216 0 2.0 1e-06 
0.0 1.1217 0 2.0 1e-06 
0.0 1.1218 0 2.0 1e-06 
0.0 1.1219 0 2.0 1e-06 
0.0 1.122 0 2.0 1e-06 
0.0 1.1221 0 2.0 1e-06 
0.0 1.1222 0 2.0 1e-06 
0.0 1.1223 0 2.0 1e-06 
0.0 1.1224 0 2.0 1e-06 
0.0 1.1225 0 2.0 1e-06 
0.0 1.1226 0 2.0 1e-06 
0.0 1.1227 0 2.0 1e-06 
0.0 1.1228 0 2.0 1e-06 
0.0 1.1229 0 2.0 1e-06 
0.0 1.123 0 2.0 1e-06 
0.0 1.1231 0 2.0 1e-06 
0.0 1.1232 0 2.0 1e-06 
0.0 1.1233 0 2.0 1e-06 
0.0 1.1234 0 2.0 1e-06 
0.0 1.1235 0 2.0 1e-06 
0.0 1.1236 0 2.0 1e-06 
0.0 1.1237 0 2.0 1e-06 
0.0 1.1238 0 2.0 1e-06 
0.0 1.1239 0 2.0 1e-06 
0.0 1.124 0 2.0 1e-06 
0.0 1.1241 0 2.0 1e-06 
0.0 1.1242 0 2.0 1e-06 
0.0 1.1243 0 2.0 1e-06 
0.0 1.1244 0 2.0 1e-06 
0.0 1.1245 0 2.0 1e-06 
0.0 1.1246 0 2.0 1e-06 
0.0 1.1247 0 2.0 1e-06 
0.0 1.1248 0 2.0 1e-06 
0.0 1.1249 0 2.0 1e-06 
0.0 1.125 0 2.0 1e-06 
0.0 1.1251 0 2.0 1e-06 
0.0 1.1252 0 2.0 1e-06 
0.0 1.1253 0 2.0 1e-06 
0.0 1.1254 0 2.0 1e-06 
0.0 1.1255 0 2.0 1e-06 
0.0 1.1256 0 2.0 1e-06 
0.0 1.1257 0 2.0 1e-06 
0.0 1.1258 0 2.0 1e-06 
0.0 1.1259 0 2.0 1e-06 
0.0 1.126 0 2.0 1e-06 
0.0 1.1261 0 2.0 1e-06 
0.0 1.1262 0 2.0 1e-06 
0.0 1.1263 0 2.0 1e-06 
0.0 1.1264 0 2.0 1e-06 
0.0 1.1265 0 2.0 1e-06 
0.0 1.1266 0 2.0 1e-06 
0.0 1.1267 0 2.0 1e-06 
0.0 1.1268 0 2.0 1e-06 
0.0 1.1269 0 2.0 1e-06 
0.0 1.127 0 2.0 1e-06 
0.0 1.1271 0 2.0 1e-06 
0.0 1.1272 0 2.0 1e-06 
0.0 1.1273 0 2.0 1e-06 
0.0 1.1274 0 2.0 1e-06 
0.0 1.1275 0 2.0 1e-06 
0.0 1.1276 0 2.0 1e-06 
0.0 1.1277 0 2.0 1e-06 
0.0 1.1278 0 2.0 1e-06 
0.0 1.1279 0 2.0 1e-06 
0.0 1.128 0 2.0 1e-06 
0.0 1.1281 0 2.0 1e-06 
0.0 1.1282 0 2.0 1e-06 
0.0 1.1283 0 2.0 1e-06 
0.0 1.1284 0 2.0 1e-06 
0.0 1.1285 0 2.0 1e-06 
0.0 1.1286 0 2.0 1e-06 
0.0 1.1287 0 2.0 1e-06 
0.0 1.1288 0 2.0 1e-06 
0.0 1.1289 0 2.0 1e-06 
0.0 1.129 0 2.0 1e-06 
0.0 1.1291 0 2.0 1e-06 
0.0 1.1292 0 2.0 1e-06 
0.0 1.1293 0 2.0 1e-06 
0.0 1.1294 0 2.0 1e-06 
0.0 1.1295 0 2.0 1e-06 
0.0 1.1296 0 2.0 1e-06 
0.0 1.1297 0 2.0 1e-06 
0.0 1.1298 0 2.0 1e-06 
0.0 1.1299 0 2.0 1e-06 
0.0 1.13 0 2.0 1e-06 
0.0 1.1301 0 2.0 1e-06 
0.0 1.1302 0 2.0 1e-06 
0.0 1.1303 0 2.0 1e-06 
0.0 1.1304 0 2.0 1e-06 
0.0 1.1305 0 2.0 1e-06 
0.0 1.1306 0 2.0 1e-06 
0.0 1.1307 0 2.0 1e-06 
0.0 1.1308 0 2.0 1e-06 
0.0 1.1309 0 2.0 1e-06 
0.0 1.131 0 2.0 1e-06 
0.0 1.1311 0 2.0 1e-06 
0.0 1.1312 0 2.0 1e-06 
0.0 1.1313 0 2.0 1e-06 
0.0 1.1314 0 2.0 1e-06 
0.0 1.1315 0 2.0 1e-06 
0.0 1.1316 0 2.0 1e-06 
0.0 1.1317 0 2.0 1e-06 
0.0 1.1318 0 2.0 1e-06 
0.0 1.1319 0 2.0 1e-06 
0.0 1.132 0 2.0 1e-06 
0.0 1.1321 0 2.0 1e-06 
0.0 1.1322 0 2.0 1e-06 
0.0 1.1323 0 2.0 1e-06 
0.0 1.1324 0 2.0 1e-06 
0.0 1.1325 0 2.0 1e-06 
0.0 1.1326 0 2.0 1e-06 
0.0 1.1327 0 2.0 1e-06 
0.0 1.1328 0 2.0 1e-06 
0.0 1.1329 0 2.0 1e-06 
0.0 1.133 0 2.0 1e-06 
0.0 1.1331 0 2.0 1e-06 
0.0 1.1332 0 2.0 1e-06 
0.0 1.1333 0 2.0 1e-06 
0.0 1.1334 0 2.0 1e-06 
0.0 1.1335 0 2.0 1e-06 
0.0 1.1336 0 2.0 1e-06 
0.0 1.1337 0 2.0 1e-06 
0.0 1.1338 0 2.0 1e-06 
0.0 1.1339 0 2.0 1e-06 
0.0 1.134 0 2.0 1e-06 
0.0 1.1341 0 2.0 1e-06 
0.0 1.1342 0 2.0 1e-06 
0.0 1.1343 0 2.0 1e-06 
0.0 1.1344 0 2.0 1e-06 
0.0 1.1345 0 2.0 1e-06 
0.0 1.1346 0 2.0 1e-06 
0.0 1.1347 0 2.0 1e-06 
0.0 1.1348 0 2.0 1e-06 
0.0 1.1349 0 2.0 1e-06 
0.0 1.135 0 2.0 1e-06 
0.0 1.1351 0 2.0 1e-06 
0.0 1.1352 0 2.0 1e-06 
0.0 1.1353 0 2.0 1e-06 
0.0 1.1354 0 2.0 1e-06 
0.0 1.1355 0 2.0 1e-06 
0.0 1.1356 0 2.0 1e-06 
0.0 1.1357 0 2.0 1e-06 
0.0 1.1358 0 2.0 1e-06 
0.0 1.1359 0 2.0 1e-06 
0.0 1.136 0 2.0 1e-06 
0.0 1.1361 0 2.0 1e-06 
0.0 1.1362 0 2.0 1e-06 
0.0 1.1363 0 2.0 1e-06 
0.0 1.1364 0 2.0 1e-06 
0.0 1.1365 0 2.0 1e-06 
0.0 1.1366 0 2.0 1e-06 
0.0 1.1367 0 2.0 1e-06 
0.0 1.1368 0 2.0 1e-06 
0.0 1.1369 0 2.0 1e-06 
0.0 1.137 0 2.0 1e-06 
0.0 1.1371 0 2.0 1e-06 
0.0 1.1372 0 2.0 1e-06 
0.0 1.1373 0 2.0 1e-06 
0.0 1.1374 0 2.0 1e-06 
0.0 1.1375 0 2.0 1e-06 
0.0 1.1376 0 2.0 1e-06 
0.0 1.1377 0 2.0 1e-06 
0.0 1.1378 0 2.0 1e-06 
0.0 1.1379 0 2.0 1e-06 
0.0 1.138 0 2.0 1e-06 
0.0 1.1381 0 2.0 1e-06 
0.0 1.1382 0 2.0 1e-06 
0.0 1.1383 0 2.0 1e-06 
0.0 1.1384 0 2.0 1e-06 
0.0 1.1385 0 2.0 1e-06 
0.0 1.1386 0 2.0 1e-06 
0.0 1.1387 0 2.0 1e-06 
0.0 1.1388 0 2.0 1e-06 
0.0 1.1389 0 2.0 1e-06 
0.0 1.139 0 2.0 1e-06 
0.0 1.1391 0 2.0 1e-06 
0.0 1.1392 0 2.0 1e-06 
0.0 1.1393 0 2.0 1e-06 
0.0 1.1394 0 2.0 1e-06 
0.0 1.1395 0 2.0 1e-06 
0.0 1.1396 0 2.0 1e-06 
0.0 1.1397 0 2.0 1e-06 
0.0 1.1398 0 2.0 1e-06 
0.0 1.1399 0 2.0 1e-06 
0.0 1.14 0 2.0 1e-06 
0.0 1.1401 0 2.0 1e-06 
0.0 1.1402 0 2.0 1e-06 
0.0 1.1403 0 2.0 1e-06 
0.0 1.1404 0 2.0 1e-06 
0.0 1.1405 0 2.0 1e-06 
0.0 1.1406 0 2.0 1e-06 
0.0 1.1407 0 2.0 1e-06 
0.0 1.1408 0 2.0 1e-06 
0.0 1.1409 0 2.0 1e-06 
0.0 1.141 0 2.0 1e-06 
0.0 1.1411 0 2.0 1e-06 
0.0 1.1412 0 2.0 1e-06 
0.0 1.1413 0 2.0 1e-06 
0.0 1.1414 0 2.0 1e-06 
0.0 1.1415 0 2.0 1e-06 
0.0 1.1416 0 2.0 1e-06 
0.0 1.1417 0 2.0 1e-06 
0.0 1.1418 0 2.0 1e-06 
0.0 1.1419 0 2.0 1e-06 
0.0 1.142 0 2.0 1e-06 
0.0 1.1421 0 2.0 1e-06 
0.0 1.1422 0 2.0 1e-06 
0.0 1.1423 0 2.0 1e-06 
0.0 1.1424 0 2.0 1e-06 
0.0 1.1425 0 2.0 1e-06 
0.0 1.1426 0 2.0 1e-06 
0.0 1.1427 0 2.0 1e-06 
0.0 1.1428 0 2.0 1e-06 
0.0 1.1429 0 2.0 1e-06 
0.0 1.143 0 2.0 1e-06 
0.0 1.1431 0 2.0 1e-06 
0.0 1.1432 0 2.0 1e-06 
0.0 1.1433 0 2.0 1e-06 
0.0 1.1434 0 2.0 1e-06 
0.0 1.1435 0 2.0 1e-06 
0.0 1.1436 0 2.0 1e-06 
0.0 1.1437 0 2.0 1e-06 
0.0 1.1438 0 2.0 1e-06 
0.0 1.1439 0 2.0 1e-06 
0.0 1.144 0 2.0 1e-06 
0.0 1.1441 0 2.0 1e-06 
0.0 1.1442 0 2.0 1e-06 
0.0 1.1443 0 2.0 1e-06 
0.0 1.1444 0 2.0 1e-06 
0.0 1.1445 0 2.0 1e-06 
0.0 1.1446 0 2.0 1e-06 
0.0 1.1447 0 2.0 1e-06 
0.0 1.1448 0 2.0 1e-06 
0.0 1.1449 0 2.0 1e-06 
0.0 1.145 0 2.0 1e-06 
0.0 1.1451 0 2.0 1e-06 
0.0 1.1452 0 2.0 1e-06 
0.0 1.1453 0 2.0 1e-06 
0.0 1.1454 0 2.0 1e-06 
0.0 1.1455 0 2.0 1e-06 
0.0 1.1456 0 2.0 1e-06 
0.0 1.1457 0 2.0 1e-06 
0.0 1.1458 0 2.0 1e-06 
0.0 1.1459 0 2.0 1e-06 
0.0 1.146 0 2.0 1e-06 
0.0 1.1461 0 2.0 1e-06 
0.0 1.1462 0 2.0 1e-06 
0.0 1.1463 0 2.0 1e-06 
0.0 1.1464 0 2.0 1e-06 
0.0 1.1465 0 2.0 1e-06 
0.0 1.1466 0 2.0 1e-06 
0.0 1.1467 0 2.0 1e-06 
0.0 1.1468 0 2.0 1e-06 
0.0 1.1469 0 2.0 1e-06 
0.0 1.147 0 2.0 1e-06 
0.0 1.1471 0 2.0 1e-06 
0.0 1.1472 0 2.0 1e-06 
0.0 1.1473 0 2.0 1e-06 
0.0 1.1474 0 2.0 1e-06 
0.0 1.1475 0 2.0 1e-06 
0.0 1.1476 0 2.0 1e-06 
0.0 1.1477 0 2.0 1e-06 
0.0 1.1478 0 2.0 1e-06 
0.0 1.1479 0 2.0 1e-06 
0.0 1.148 0 2.0 1e-06 
0.0 1.1481 0 2.0 1e-06 
0.0 1.1482 0 2.0 1e-06 
0.0 1.1483 0 2.0 1e-06 
0.0 1.1484 0 2.0 1e-06 
0.0 1.1485 0 2.0 1e-06 
0.0 1.1486 0 2.0 1e-06 
0.0 1.1487 0 2.0 1e-06 
0.0 1.1488 0 2.0 1e-06 
0.0 1.1489 0 2.0 1e-06 
0.0 1.149 0 2.0 1e-06 
0.0 1.1491 0 2.0 1e-06 
0.0 1.1492 0 2.0 1e-06 
0.0 1.1493 0 2.0 1e-06 
0.0 1.1494 0 2.0 1e-06 
0.0 1.1495 0 2.0 1e-06 
0.0 1.1496 0 2.0 1e-06 
0.0 1.1497 0 2.0 1e-06 
0.0 1.1498 0 2.0 1e-06 
0.0 1.1499 0 2.0 1e-06 
0.0 1.15 0 2.0 1e-06 
0.0 1.1501 0 2.0 1e-06 
0.0 1.1502 0 2.0 1e-06 
0.0 1.1503 0 2.0 1e-06 
0.0 1.1504 0 2.0 1e-06 
0.0 1.1505 0 2.0 1e-06 
0.0 1.1506 0 2.0 1e-06 
0.0 1.1507 0 2.0 1e-06 
0.0 1.1508 0 2.0 1e-06 
0.0 1.1509 0 2.0 1e-06 
0.0 1.151 0 2.0 1e-06 
0.0 1.1511 0 2.0 1e-06 
0.0 1.1512 0 2.0 1e-06 
0.0 1.1513 0 2.0 1e-06 
0.0 1.1514 0 2.0 1e-06 
0.0 1.1515 0 2.0 1e-06 
0.0 1.1516 0 2.0 1e-06 
0.0 1.1517 0 2.0 1e-06 
0.0 1.1518 0 2.0 1e-06 
0.0 1.1519 0 2.0 1e-06 
0.0 1.152 0 2.0 1e-06 
0.0 1.1521 0 2.0 1e-06 
0.0 1.1522 0 2.0 1e-06 
0.0 1.1523 0 2.0 1e-06 
0.0 1.1524 0 2.0 1e-06 
0.0 1.1525 0 2.0 1e-06 
0.0 1.1526 0 2.0 1e-06 
0.0 1.1527 0 2.0 1e-06 
0.0 1.1528 0 2.0 1e-06 
0.0 1.1529 0 2.0 1e-06 
0.0 1.153 0 2.0 1e-06 
0.0 1.1531 0 2.0 1e-06 
0.0 1.1532 0 2.0 1e-06 
0.0 1.1533 0 2.0 1e-06 
0.0 1.1534 0 2.0 1e-06 
0.0 1.1535 0 2.0 1e-06 
0.0 1.1536 0 2.0 1e-06 
0.0 1.1537 0 2.0 1e-06 
0.0 1.1538 0 2.0 1e-06 
0.0 1.1539 0 2.0 1e-06 
0.0 1.154 0 2.0 1e-06 
0.0 1.1541 0 2.0 1e-06 
0.0 1.1542 0 2.0 1e-06 
0.0 1.1543 0 2.0 1e-06 
0.0 1.1544 0 2.0 1e-06 
0.0 1.1545 0 2.0 1e-06 
0.0 1.1546 0 2.0 1e-06 
0.0 1.1547 0 2.0 1e-06 
0.0 1.1548 0 2.0 1e-06 
0.0 1.1549 0 2.0 1e-06 
0.0 1.155 0 2.0 1e-06 
0.0 1.1551 0 2.0 1e-06 
0.0 1.1552 0 2.0 1e-06 
0.0 1.1553 0 2.0 1e-06 
0.0 1.1554 0 2.0 1e-06 
0.0 1.1555 0 2.0 1e-06 
0.0 1.1556 0 2.0 1e-06 
0.0 1.1557 0 2.0 1e-06 
0.0 1.1558 0 2.0 1e-06 
0.0 1.1559 0 2.0 1e-06 
0.0 1.156 0 2.0 1e-06 
0.0 1.1561 0 2.0 1e-06 
0.0 1.1562 0 2.0 1e-06 
0.0 1.1563 0 2.0 1e-06 
0.0 1.1564 0 2.0 1e-06 
0.0 1.1565 0 2.0 1e-06 
0.0 1.1566 0 2.0 1e-06 
0.0 1.1567 0 2.0 1e-06 
0.0 1.1568 0 2.0 1e-06 
0.0 1.1569 0 2.0 1e-06 
0.0 1.157 0 2.0 1e-06 
0.0 1.1571 0 2.0 1e-06 
0.0 1.1572 0 2.0 1e-06 
0.0 1.1573 0 2.0 1e-06 
0.0 1.1574 0 2.0 1e-06 
0.0 1.1575 0 2.0 1e-06 
0.0 1.1576 0 2.0 1e-06 
0.0 1.1577 0 2.0 1e-06 
0.0 1.1578 0 2.0 1e-06 
0.0 1.1579 0 2.0 1e-06 
0.0 1.158 0 2.0 1e-06 
0.0 1.1581 0 2.0 1e-06 
0.0 1.1582 0 2.0 1e-06 
0.0 1.1583 0 2.0 1e-06 
0.0 1.1584 0 2.0 1e-06 
0.0 1.1585 0 2.0 1e-06 
0.0 1.1586 0 2.0 1e-06 
0.0 1.1587 0 2.0 1e-06 
0.0 1.1588 0 2.0 1e-06 
0.0 1.1589 0 2.0 1e-06 
0.0 1.159 0 2.0 1e-06 
0.0 1.1591 0 2.0 1e-06 
0.0 1.1592 0 2.0 1e-06 
0.0 1.1593 0 2.0 1e-06 
0.0 1.1594 0 2.0 1e-06 
0.0 1.1595 0 2.0 1e-06 
0.0 1.1596 0 2.0 1e-06 
0.0 1.1597 0 2.0 1e-06 
0.0 1.1598 0 2.0 1e-06 
0.0 1.1599 0 2.0 1e-06 
0.0 1.16 0 2.0 1e-06 
0.0 1.1601 0 2.0 1e-06 
0.0 1.1602 0 2.0 1e-06 
0.0 1.1603 0 2.0 1e-06 
0.0 1.1604 0 2.0 1e-06 
0.0 1.1605 0 2.0 1e-06 
0.0 1.1606 0 2.0 1e-06 
0.0 1.1607 0 2.0 1e-06 
0.0 1.1608 0 2.0 1e-06 
0.0 1.1609 0 2.0 1e-06 
0.0 1.161 0 2.0 1e-06 
0.0 1.1611 0 2.0 1e-06 
0.0 1.1612 0 2.0 1e-06 
0.0 1.1613 0 2.0 1e-06 
0.0 1.1614 0 2.0 1e-06 
0.0 1.1615 0 2.0 1e-06 
0.0 1.1616 0 2.0 1e-06 
0.0 1.1617 0 2.0 1e-06 
0.0 1.1618 0 2.0 1e-06 
0.0 1.1619 0 2.0 1e-06 
0.0 1.162 0 2.0 1e-06 
0.0 1.1621 0 2.0 1e-06 
0.0 1.1622 0 2.0 1e-06 
0.0 1.1623 0 2.0 1e-06 
0.0 1.1624 0 2.0 1e-06 
0.0 1.1625 0 2.0 1e-06 
0.0 1.1626 0 2.0 1e-06 
0.0 1.1627 0 2.0 1e-06 
0.0 1.1628 0 2.0 1e-06 
0.0 1.1629 0 2.0 1e-06 
0.0 1.163 0 2.0 1e-06 
0.0 1.1631 0 2.0 1e-06 
0.0 1.1632 0 2.0 1e-06 
0.0 1.1633 0 2.0 1e-06 
0.0 1.1634 0 2.0 1e-06 
0.0 1.1635 0 2.0 1e-06 
0.0 1.1636 0 2.0 1e-06 
0.0 1.1637 0 2.0 1e-06 
0.0 1.1638 0 2.0 1e-06 
0.0 1.1639 0 2.0 1e-06 
0.0 1.164 0 2.0 1e-06 
0.0 1.1641 0 2.0 1e-06 
0.0 1.1642 0 2.0 1e-06 
0.0 1.1643 0 2.0 1e-06 
0.0 1.1644 0 2.0 1e-06 
0.0 1.1645 0 2.0 1e-06 
0.0 1.1646 0 2.0 1e-06 
0.0 1.1647 0 2.0 1e-06 
0.0 1.1648 0 2.0 1e-06 
0.0 1.1649 0 2.0 1e-06 
0.0 1.165 0 2.0 1e-06 
0.0 1.1651 0 2.0 1e-06 
0.0 1.1652 0 2.0 1e-06 
0.0 1.1653 0 2.0 1e-06 
0.0 1.1654 0 2.0 1e-06 
0.0 1.1655 0 2.0 1e-06 
0.0 1.1656 0 2.0 1e-06 
0.0 1.1657 0 2.0 1e-06 
0.0 1.1658 0 2.0 1e-06 
0.0 1.1659 0 2.0 1e-06 
0.0 1.166 0 2.0 1e-06 
0.0 1.1661 0 2.0 1e-06 
0.0 1.1662 0 2.0 1e-06 
0.0 1.1663 0 2.0 1e-06 
0.0 1.1664 0 2.0 1e-06 
0.0 1.1665 0 2.0 1e-06 
0.0 1.1666 0 2.0 1e-06 
0.0 1.1667 0 2.0 1e-06 
0.0 1.1668 0 2.0 1e-06 
0.0 1.1669 0 2.0 1e-06 
0.0 1.167 0 2.0 1e-06 
0.0 1.1671 0 2.0 1e-06 
0.0 1.1672 0 2.0 1e-06 
0.0 1.1673 0 2.0 1e-06 
0.0 1.1674 0 2.0 1e-06 
0.0 1.1675 0 2.0 1e-06 
0.0 1.1676 0 2.0 1e-06 
0.0 1.1677 0 2.0 1e-06 
0.0 1.1678 0 2.0 1e-06 
0.0 1.1679 0 2.0 1e-06 
0.0 1.168 0 2.0 1e-06 
0.0 1.1681 0 2.0 1e-06 
0.0 1.1682 0 2.0 1e-06 
0.0 1.1683 0 2.0 1e-06 
0.0 1.1684 0 2.0 1e-06 
0.0 1.1685 0 2.0 1e-06 
0.0 1.1686 0 2.0 1e-06 
0.0 1.1687 0 2.0 1e-06 
0.0 1.1688 0 2.0 1e-06 
0.0 1.1689 0 2.0 1e-06 
0.0 1.169 0 2.0 1e-06 
0.0 1.1691 0 2.0 1e-06 
0.0 1.1692 0 2.0 1e-06 
0.0 1.1693 0 2.0 1e-06 
0.0 1.1694 0 2.0 1e-06 
0.0 1.1695 0 2.0 1e-06 
0.0 1.1696 0 2.0 1e-06 
0.0 1.1697 0 2.0 1e-06 
0.0 1.1698 0 2.0 1e-06 
0.0 1.1699 0 2.0 1e-06 
0.0 1.17 0 2.0 1e-06 
0.0 1.1701 0 2.0 1e-06 
0.0 1.1702 0 2.0 1e-06 
0.0 1.1703 0 2.0 1e-06 
0.0 1.1704 0 2.0 1e-06 
0.0 1.1705 0 2.0 1e-06 
0.0 1.1706 0 2.0 1e-06 
0.0 1.1707 0 2.0 1e-06 
0.0 1.1708 0 2.0 1e-06 
0.0 1.1709 0 2.0 1e-06 
0.0 1.171 0 2.0 1e-06 
0.0 1.1711 0 2.0 1e-06 
0.0 1.1712 0 2.0 1e-06 
0.0 1.1713 0 2.0 1e-06 
0.0 1.1714 0 2.0 1e-06 
0.0 1.1715 0 2.0 1e-06 
0.0 1.1716 0 2.0 1e-06 
0.0 1.1717 0 2.0 1e-06 
0.0 1.1718 0 2.0 1e-06 
0.0 1.1719 0 2.0 1e-06 
0.0 1.172 0 2.0 1e-06 
0.0 1.1721 0 2.0 1e-06 
0.0 1.1722 0 2.0 1e-06 
0.0 1.1723 0 2.0 1e-06 
0.0 1.1724 0 2.0 1e-06 
0.0 1.1725 0 2.0 1e-06 
0.0 1.1726 0 2.0 1e-06 
0.0 1.1727 0 2.0 1e-06 
0.0 1.1728 0 2.0 1e-06 
0.0 1.1729 0 2.0 1e-06 
0.0 1.173 0 2.0 1e-06 
0.0 1.1731 0 2.0 1e-06 
0.0 1.1732 0 2.0 1e-06 
0.0 1.1733 0 2.0 1e-06 
0.0 1.1734 0 2.0 1e-06 
0.0 1.1735 0 2.0 1e-06 
0.0 1.1736 0 2.0 1e-06 
0.0 1.1737 0 2.0 1e-06 
0.0 1.1738 0 2.0 1e-06 
0.0 1.1739 0 2.0 1e-06 
0.0 1.174 0 2.0 1e-06 
0.0 1.1741 0 2.0 1e-06 
0.0 1.1742 0 2.0 1e-06 
0.0 1.1743 0 2.0 1e-06 
0.0 1.1744 0 2.0 1e-06 
0.0 1.1745 0 2.0 1e-06 
0.0 1.1746 0 2.0 1e-06 
0.0 1.1747 0 2.0 1e-06 
0.0 1.1748 0 2.0 1e-06 
0.0 1.1749 0 2.0 1e-06 
0.0 1.175 0 2.0 1e-06 
0.0 1.1751 0 2.0 1e-06 
0.0 1.1752 0 2.0 1e-06 
0.0 1.1753 0 2.0 1e-06 
0.0 1.1754 0 2.0 1e-06 
0.0 1.1755 0 2.0 1e-06 
0.0 1.1756 0 2.0 1e-06 
0.0 1.1757 0 2.0 1e-06 
0.0 1.1758 0 2.0 1e-06 
0.0 1.1759 0 2.0 1e-06 
0.0 1.176 0 2.0 1e-06 
0.0 1.1761 0 2.0 1e-06 
0.0 1.1762 0 2.0 1e-06 
0.0 1.1763 0 2.0 1e-06 
0.0 1.1764 0 2.0 1e-06 
0.0 1.1765 0 2.0 1e-06 
0.0 1.1766 0 2.0 1e-06 
0.0 1.1767 0 2.0 1e-06 
0.0 1.1768 0 2.0 1e-06 
0.0 1.1769 0 2.0 1e-06 
0.0 1.177 0 2.0 1e-06 
0.0 1.1771 0 2.0 1e-06 
0.0 1.1772 0 2.0 1e-06 
0.0 1.1773 0 2.0 1e-06 
0.0 1.1774 0 2.0 1e-06 
0.0 1.1775 0 2.0 1e-06 
0.0 1.1776 0 2.0 1e-06 
0.0 1.1777 0 2.0 1e-06 
0.0 1.1778 0 2.0 1e-06 
0.0 1.1779 0 2.0 1e-06 
0.0 1.178 0 2.0 1e-06 
0.0 1.1781 0 2.0 1e-06 
0.0 1.1782 0 2.0 1e-06 
0.0 1.1783 0 2.0 1e-06 
0.0 1.1784 0 2.0 1e-06 
0.0 1.1785 0 2.0 1e-06 
0.0 1.1786 0 2.0 1e-06 
0.0 1.1787 0 2.0 1e-06 
0.0 1.1788 0 2.0 1e-06 
0.0 1.1789 0 2.0 1e-06 
0.0 1.179 0 2.0 1e-06 
0.0 1.1791 0 2.0 1e-06 
0.0 1.1792 0 2.0 1e-06 
0.0 1.1793 0 2.0 1e-06 
0.0 1.1794 0 2.0 1e-06 
0.0 1.1795 0 2.0 1e-06 
0.0 1.1796 0 2.0 1e-06 
0.0 1.1797 0 2.0 1e-06 
0.0 1.1798 0 2.0 1e-06 
0.0 1.1799 0 2.0 1e-06 
0.0 1.18 0 2.0 1e-06 
0.0 1.1801 0 2.0 1e-06 
0.0 1.1802 0 2.0 1e-06 
0.0 1.1803 0 2.0 1e-06 
0.0 1.1804 0 2.0 1e-06 
0.0 1.1805 0 2.0 1e-06 
0.0 1.1806 0 2.0 1e-06 
0.0 1.1807 0 2.0 1e-06 
0.0 1.1808 0 2.0 1e-06 
0.0 1.1809 0 2.0 1e-06 
0.0 1.181 0 2.0 1e-06 
0.0 1.1811 0 2.0 1e-06 
0.0 1.1812 0 2.0 1e-06 
0.0 1.1813 0 2.0 1e-06 
0.0 1.1814 0 2.0 1e-06 
0.0 1.1815 0 2.0 1e-06 
0.0 1.1816 0 2.0 1e-06 
0.0 1.1817 0 2.0 1e-06 
0.0 1.1818 0 2.0 1e-06 
0.0 1.1819 0 2.0 1e-06 
0.0 1.182 0 2.0 1e-06 
0.0 1.1821 0 2.0 1e-06 
0.0 1.1822 0 2.0 1e-06 
0.0 1.1823 0 2.0 1e-06 
0.0 1.1824 0 2.0 1e-06 
0.0 1.1825 0 2.0 1e-06 
0.0 1.1826 0 2.0 1e-06 
0.0 1.1827 0 2.0 1e-06 
0.0 1.1828 0 2.0 1e-06 
0.0 1.1829 0 2.0 1e-06 
0.0 1.183 0 2.0 1e-06 
0.0 1.1831 0 2.0 1e-06 
0.0 1.1832 0 2.0 1e-06 
0.0 1.1833 0 2.0 1e-06 
0.0 1.1834 0 2.0 1e-06 
0.0 1.1835 0 2.0 1e-06 
0.0 1.1836 0 2.0 1e-06 
0.0 1.1837 0 2.0 1e-06 
0.0 1.1838 0 2.0 1e-06 
0.0 1.1839 0 2.0 1e-06 
0.0 1.184 0 2.0 1e-06 
0.0 1.1841 0 2.0 1e-06 
0.0 1.1842 0 2.0 1e-06 
0.0 1.1843 0 2.0 1e-06 
0.0 1.1844 0 2.0 1e-06 
0.0 1.1845 0 2.0 1e-06 
0.0 1.1846 0 2.0 1e-06 
0.0 1.1847 0 2.0 1e-06 
0.0 1.1848 0 2.0 1e-06 
0.0 1.1849 0 2.0 1e-06 
0.0 1.185 0 2.0 1e-06 
0.0 1.1851 0 2.0 1e-06 
0.0 1.1852 0 2.0 1e-06 
0.0 1.1853 0 2.0 1e-06 
0.0 1.1854 0 2.0 1e-06 
0.0 1.1855 0 2.0 1e-06 
0.0 1.1856 0 2.0 1e-06 
0.0 1.1857 0 2.0 1e-06 
0.0 1.1858 0 2.0 1e-06 
0.0 1.1859 0 2.0 1e-06 
0.0 1.186 0 2.0 1e-06 
0.0 1.1861 0 2.0 1e-06 
0.0 1.1862 0 2.0 1e-06 
0.0 1.1863 0 2.0 1e-06 
0.0 1.1864 0 2.0 1e-06 
0.0 1.1865 0 2.0 1e-06 
0.0 1.1866 0 2.0 1e-06 
0.0 1.1867 0 2.0 1e-06 
0.0 1.1868 0 2.0 1e-06 
0.0 1.1869 0 2.0 1e-06 
0.0 1.187 0 2.0 1e-06 
0.0 1.1871 0 2.0 1e-06 
0.0 1.1872 0 2.0 1e-06 
0.0 1.1873 0 2.0 1e-06 
0.0 1.1874 0 2.0 1e-06 
0.0 1.1875 0 2.0 1e-06 
0.0 1.1876 0 2.0 1e-06 
0.0 1.1877 0 2.0 1e-06 
0.0 1.1878 0 2.0 1e-06 
0.0 1.1879 0 2.0 1e-06 
0.0 1.188 0 2.0 1e-06 
0.0 1.1881 0 2.0 1e-06 
0.0 1.1882 0 2.0 1e-06 
0.0 1.1883 0 2.0 1e-06 
0.0 1.1884 0 2.0 1e-06 
0.0 1.1885 0 2.0 1e-06 
0.0 1.1886 0 2.0 1e-06 
0.0 1.1887 0 2.0 1e-06 
0.0 1.1888 0 2.0 1e-06 
0.0 1.1889 0 2.0 1e-06 
0.0 1.189 0 2.0 1e-06 
0.0 1.1891 0 2.0 1e-06 
0.0 1.1892 0 2.0 1e-06 
0.0 1.1893 0 2.0 1e-06 
0.0 1.1894 0 2.0 1e-06 
0.0 1.1895 0 2.0 1e-06 
0.0 1.1896 0 2.0 1e-06 
0.0 1.1897 0 2.0 1e-06 
0.0 1.1898 0 2.0 1e-06 
0.0 1.1899 0 2.0 1e-06 
0.0 1.19 0 2.0 1e-06 
0.0 1.1901 0 2.0 1e-06 
0.0 1.1902 0 2.0 1e-06 
0.0 1.1903 0 2.0 1e-06 
0.0 1.1904 0 2.0 1e-06 
0.0 1.1905 0 2.0 1e-06 
0.0 1.1906 0 2.0 1e-06 
0.0 1.1907 0 2.0 1e-06 
0.0 1.1908 0 2.0 1e-06 
0.0 1.1909 0 2.0 1e-06 
0.0 1.191 0 2.0 1e-06 
0.0 1.1911 0 2.0 1e-06 
0.0 1.1912 0 2.0 1e-06 
0.0 1.1913 0 2.0 1e-06 
0.0 1.1914 0 2.0 1e-06 
0.0 1.1915 0 2.0 1e-06 
0.0 1.1916 0 2.0 1e-06 
0.0 1.1917 0 2.0 1e-06 
0.0 1.1918 0 2.0 1e-06 
0.0 1.1919 0 2.0 1e-06 
0.0 1.192 0 2.0 1e-06 
0.0 1.1921 0 2.0 1e-06 
0.0 1.1922 0 2.0 1e-06 
0.0 1.1923 0 2.0 1e-06 
0.0 1.1924 0 2.0 1e-06 
0.0 1.1925 0 2.0 1e-06 
0.0 1.1926 0 2.0 1e-06 
0.0 1.1927 0 2.0 1e-06 
0.0 1.1928 0 2.0 1e-06 
0.0 1.1929 0 2.0 1e-06 
0.0 1.193 0 2.0 1e-06 
0.0 1.1931 0 2.0 1e-06 
0.0 1.1932 0 2.0 1e-06 
0.0 1.1933 0 2.0 1e-06 
0.0 1.1934 0 2.0 1e-06 
0.0 1.1935 0 2.0 1e-06 
0.0 1.1936 0 2.0 1e-06 
0.0 1.1937 0 2.0 1e-06 
0.0 1.1938 0 2.0 1e-06 
0.0 1.1939 0 2.0 1e-06 
0.0 1.194 0 2.0 1e-06 
0.0 1.1941 0 2.0 1e-06 
0.0 1.1942 0 2.0 1e-06 
0.0 1.1943 0 2.0 1e-06 
0.0 1.1944 0 2.0 1e-06 
0.0 1.1945 0 2.0 1e-06 
0.0 1.1946 0 2.0 1e-06 
0.0 1.1947 0 2.0 1e-06 
0.0 1.1948 0 2.0 1e-06 
0.0 1.1949 0 2.0 1e-06 
0.0 1.195 0 2.0 1e-06 
0.0 1.1951 0 2.0 1e-06 
0.0 1.1952 0 2.0 1e-06 
0.0 1.1953 0 2.0 1e-06 
0.0 1.1954 0 2.0 1e-06 
0.0 1.1955 0 2.0 1e-06 
0.0 1.1956 0 2.0 1e-06 
0.0 1.1957 0 2.0 1e-06 
0.0 1.1958 0 2.0 1e-06 
0.0 1.1959 0 2.0 1e-06 
0.0 1.196 0 2.0 1e-06 
0.0 1.1961 0 2.0 1e-06 
0.0 1.1962 0 2.0 1e-06 
0.0 1.1963 0 2.0 1e-06 
0.0 1.1964 0 2.0 1e-06 
0.0 1.1965 0 2.0 1e-06 
0.0 1.1966 0 2.0 1e-06 
0.0 1.1967 0 2.0 1e-06 
0.0 1.1968 0 2.0 1e-06 
0.0 1.1969 0 2.0 1e-06 
0.0 1.197 0 2.0 1e-06 
0.0 1.1971 0 2.0 1e-06 
0.0 1.1972 0 2.0 1e-06 
0.0 1.1973 0 2.0 1e-06 
0.0 1.1974 0 2.0 1e-06 
0.0 1.1975 0 2.0 1e-06 
0.0 1.1976 0 2.0 1e-06 
0.0 1.1977 0 2.0 1e-06 
0.0 1.1978 0 2.0 1e-06 
0.0 1.1979 0 2.0 1e-06 
0.0 1.198 0 2.0 1e-06 
0.0 1.1981 0 2.0 1e-06 
0.0 1.1982 0 2.0 1e-06 
0.0 1.1983 0 2.0 1e-06 
0.0 1.1984 0 2.0 1e-06 
0.0 1.1985 0 2.0 1e-06 
0.0 1.1986 0 2.0 1e-06 
0.0 1.1987 0 2.0 1e-06 
0.0 1.1988 0 2.0 1e-06 
0.0 1.1989 0 2.0 1e-06 
0.0 1.199 0 2.0 1e-06 
0.0 1.1991 0 2.0 1e-06 
0.0 1.1992 0 2.0 1e-06 
0.0 1.1993 0 2.0 1e-06 
0.0 1.1994 0 2.0 1e-06 
0.0 1.1995 0 2.0 1e-06 
0.0 1.1996 0 2.0 1e-06 
0.0 1.1997 0 2.0 1e-06 
0.0 1.1998 0 2.0 1e-06 
0.0 1.1999 0 2.0 1e-06 
0.0 1.2 0 2.0 1e-06 
0.0 1.2001 0 2.0 1e-06 
0.0 1.2002 0 2.0 1e-06 
0.0 1.2003 0 2.0 1e-06 
0.0 1.2004 0 2.0 1e-06 
0.0 1.2005 0 2.0 1e-06 
0.0 1.2006 0 2.0 1e-06 
0.0 1.2007 0 2.0 1e-06 
0.0 1.2008 0 2.0 1e-06 
0.0 1.2009 0 2.0 1e-06 
0.0 1.201 0 2.0 1e-06 
0.0 1.2011 0 2.0 1e-06 
0.0 1.2012 0 2.0 1e-06 
0.0 1.2013 0 2.0 1e-06 
0.0 1.2014 0 2.0 1e-06 
0.0 1.2015 0 2.0 1e-06 
0.0 1.2016 0 2.0 1e-06 
0.0 1.2017 0 2.0 1e-06 
0.0 1.2018 0 2.0 1e-06 
0.0 1.2019 0 2.0 1e-06 
0.0 1.202 0 2.0 1e-06 
0.0 1.2021 0 2.0 1e-06 
0.0 1.2022 0 2.0 1e-06 
0.0 1.2023 0 2.0 1e-06 
0.0 1.2024 0 2.0 1e-06 
0.0 1.2025 0 2.0 1e-06 
0.0 1.2026 0 2.0 1e-06 
0.0 1.2027 0 2.0 1e-06 
0.0 1.2028 0 2.0 1e-06 
0.0 1.2029 0 2.0 1e-06 
0.0 1.203 0 2.0 1e-06 
0.0 1.2031 0 2.0 1e-06 
0.0 1.2032 0 2.0 1e-06 
0.0 1.2033 0 2.0 1e-06 
0.0 1.2034 0 2.0 1e-06 
0.0 1.2035 0 2.0 1e-06 
0.0 1.2036 0 2.0 1e-06 
0.0 1.2037 0 2.0 1e-06 
0.0 1.2038 0 2.0 1e-06 
0.0 1.2039 0 2.0 1e-06 
0.0 1.204 0 2.0 1e-06 
0.0 1.2041 0 2.0 1e-06 
0.0 1.2042 0 2.0 1e-06 
0.0 1.2043 0 2.0 1e-06 
0.0 1.2044 0 2.0 1e-06 
0.0 1.2045 0 2.0 1e-06 
0.0 1.2046 0 2.0 1e-06 
0.0 1.2047 0 2.0 1e-06 
0.0 1.2048 0 2.0 1e-06 
0.0 1.2049 0 2.0 1e-06 
0.0 1.205 0 2.0 1e-06 
0.0 1.2051 0 2.0 1e-06 
0.0 1.2052 0 2.0 1e-06 
0.0 1.2053 0 2.0 1e-06 
0.0 1.2054 0 2.0 1e-06 
0.0 1.2055 0 2.0 1e-06 
0.0 1.2056 0 2.0 1e-06 
0.0 1.2057 0 2.0 1e-06 
0.0 1.2058 0 2.0 1e-06 
0.0 1.2059 0 2.0 1e-06 
0.0 1.206 0 2.0 1e-06 
0.0 1.2061 0 2.0 1e-06 
0.0 1.2062 0 2.0 1e-06 
0.0 1.2063 0 2.0 1e-06 
0.0 1.2064 0 2.0 1e-06 
0.0 1.2065 0 2.0 1e-06 
0.0 1.2066 0 2.0 1e-06 
0.0 1.2067 0 2.0 1e-06 
0.0 1.2068 0 2.0 1e-06 
0.0 1.2069 0 2.0 1e-06 
0.0 1.207 0 2.0 1e-06 
0.0 1.2071 0 2.0 1e-06 
0.0 1.2072 0 2.0 1e-06 
0.0 1.2073 0 2.0 1e-06 
0.0 1.2074 0 2.0 1e-06 
0.0 1.2075 0 2.0 1e-06 
0.0 1.2076 0 2.0 1e-06 
0.0 1.2077 0 2.0 1e-06 
0.0 1.2078 0 2.0 1e-06 
0.0 1.2079 0 2.0 1e-06 
0.0 1.208 0 2.0 1e-06 
0.0 1.2081 0 2.0 1e-06 
0.0 1.2082 0 2.0 1e-06 
0.0 1.2083 0 2.0 1e-06 
0.0 1.2084 0 2.0 1e-06 
0.0 1.2085 0 2.0 1e-06 
0.0 1.2086 0 2.0 1e-06 
0.0 1.2087 0 2.0 1e-06 
0.0 1.2088 0 2.0 1e-06 
0.0 1.2089 0 2.0 1e-06 
0.0 1.209 0 2.0 1e-06 
0.0 1.2091 0 2.0 1e-06 
0.0 1.2092 0 2.0 1e-06 
0.0 1.2093 0 2.0 1e-06 
0.0 1.2094 0 2.0 1e-06 
0.0 1.2095 0 2.0 1e-06 
0.0 1.2096 0 2.0 1e-06 
0.0 1.2097 0 2.0 1e-06 
0.0 1.2098 0 2.0 1e-06 
0.0 1.2099 0 2.0 1e-06 
0.0 1.21 0 2.0 1e-06 
0.0 1.2101 0 2.0 1e-06 
0.0 1.2102 0 2.0 1e-06 
0.0 1.2103 0 2.0 1e-06 
0.0 1.2104 0 2.0 1e-06 
0.0 1.2105 0 2.0 1e-06 
0.0 1.2106 0 2.0 1e-06 
0.0 1.2107 0 2.0 1e-06 
0.0 1.2108 0 2.0 1e-06 
0.0 1.2109 0 2.0 1e-06 
0.0 1.211 0 2.0 1e-06 
0.0 1.2111 0 2.0 1e-06 
0.0 1.2112 0 2.0 1e-06 
0.0 1.2113 0 2.0 1e-06 
0.0 1.2114 0 2.0 1e-06 
0.0 1.2115 0 2.0 1e-06 
0.0 1.2116 0 2.0 1e-06 
0.0 1.2117 0 2.0 1e-06 
0.0 1.2118 0 2.0 1e-06 
0.0 1.2119 0 2.0 1e-06 
0.0 1.212 0 2.0 1e-06 
0.0 1.2121 0 2.0 1e-06 
0.0 1.2122 0 2.0 1e-06 
0.0 1.2123 0 2.0 1e-06 
0.0 1.2124 0 2.0 1e-06 
0.0 1.2125 0 2.0 1e-06 
0.0 1.2126 0 2.0 1e-06 
0.0 1.2127 0 2.0 1e-06 
0.0 1.2128 0 2.0 1e-06 
0.0 1.2129 0 2.0 1e-06 
0.0 1.213 0 2.0 1e-06 
0.0 1.2131 0 2.0 1e-06 
0.0 1.2132 0 2.0 1e-06 
0.0 1.2133 0 2.0 1e-06 
0.0 1.2134 0 2.0 1e-06 
0.0 1.2135 0 2.0 1e-06 
0.0 1.2136 0 2.0 1e-06 
0.0 1.2137 0 2.0 1e-06 
0.0 1.2138 0 2.0 1e-06 
0.0 1.2139 0 2.0 1e-06 
0.0 1.214 0 2.0 1e-06 
0.0 1.2141 0 2.0 1e-06 
0.0 1.2142 0 2.0 1e-06 
0.0 1.2143 0 2.0 1e-06 
0.0 1.2144 0 2.0 1e-06 
0.0 1.2145 0 2.0 1e-06 
0.0 1.2146 0 2.0 1e-06 
0.0 1.2147 0 2.0 1e-06 
0.0 1.2148 0 2.0 1e-06 
0.0 1.2149 0 2.0 1e-06 
0.0 1.215 0 2.0 1e-06 
0.0 1.2151 0 2.0 1e-06 
0.0 1.2152 0 2.0 1e-06 
0.0 1.2153 0 2.0 1e-06 
0.0 1.2154 0 2.0 1e-06 
0.0 1.2155 0 2.0 1e-06 
0.0 1.2156 0 2.0 1e-06 
0.0 1.2157 0 2.0 1e-06 
0.0 1.2158 0 2.0 1e-06 
0.0 1.2159 0 2.0 1e-06 
0.0 1.216 0 2.0 1e-06 
0.0 1.2161 0 2.0 1e-06 
0.0 1.2162 0 2.0 1e-06 
0.0 1.2163 0 2.0 1e-06 
0.0 1.2164 0 2.0 1e-06 
0.0 1.2165 0 2.0 1e-06 
0.0 1.2166 0 2.0 1e-06 
0.0 1.2167 0 2.0 1e-06 
0.0 1.2168 0 2.0 1e-06 
0.0 1.2169 0 2.0 1e-06 
0.0 1.217 0 2.0 1e-06 
0.0 1.2171 0 2.0 1e-06 
0.0 1.2172 0 2.0 1e-06 
0.0 1.2173 0 2.0 1e-06 
0.0 1.2174 0 2.0 1e-06 
0.0 1.2175 0 2.0 1e-06 
0.0 1.2176 0 2.0 1e-06 
0.0 1.2177 0 2.0 1e-06 
0.0 1.2178 0 2.0 1e-06 
0.0 1.2179 0 2.0 1e-06 
0.0 1.218 0 2.0 1e-06 
0.0 1.2181 0 2.0 1e-06 
0.0 1.2182 0 2.0 1e-06 
0.0 1.2183 0 2.0 1e-06 
0.0 1.2184 0 2.0 1e-06 
0.0 1.2185 0 2.0 1e-06 
0.0 1.2186 0 2.0 1e-06 
0.0 1.2187 0 2.0 1e-06 
0.0 1.2188 0 2.0 1e-06 
0.0 1.2189 0 2.0 1e-06 
0.0 1.219 0 2.0 1e-06 
0.0 1.2191 0 2.0 1e-06 
0.0 1.2192 0 2.0 1e-06 
0.0 1.2193 0 2.0 1e-06 
0.0 1.2194 0 2.0 1e-06 
0.0 1.2195 0 2.0 1e-06 
0.0 1.2196 0 2.0 1e-06 
0.0 1.2197 0 2.0 1e-06 
0.0 1.2198 0 2.0 1e-06 
0.0 1.2199 0 2.0 1e-06 
0.0 1.22 0 2.0 1e-06 
0.0 1.2201 0 2.0 1e-06 
0.0 1.2202 0 2.0 1e-06 
0.0 1.2203 0 2.0 1e-06 
0.0 1.2204 0 2.0 1e-06 
0.0 1.2205 0 2.0 1e-06 
0.0 1.2206 0 2.0 1e-06 
0.0 1.2207 0 2.0 1e-06 
0.0 1.2208 0 2.0 1e-06 
0.0 1.2209 0 2.0 1e-06 
0.0 1.221 0 2.0 1e-06 
0.0 1.2211 0 2.0 1e-06 
0.0 1.2212 0 2.0 1e-06 
0.0 1.2213 0 2.0 1e-06 
0.0 1.2214 0 2.0 1e-06 
0.0 1.2215 0 2.0 1e-06 
0.0 1.2216 0 2.0 1e-06 
0.0 1.2217 0 2.0 1e-06 
0.0 1.2218 0 2.0 1e-06 
0.0 1.2219 0 2.0 1e-06 
0.0 1.222 0 2.0 1e-06 
0.0 1.2221 0 2.0 1e-06 
0.0 1.2222 0 2.0 1e-06 
0.0 1.2223 0 2.0 1e-06 
0.0 1.2224 0 2.0 1e-06 
0.0 1.2225 0 2.0 1e-06 
0.0 1.2226 0 2.0 1e-06 
0.0 1.2227 0 2.0 1e-06 
0.0 1.2228 0 2.0 1e-06 
0.0 1.2229 0 2.0 1e-06 
0.0 1.223 0 2.0 1e-06 
0.0 1.2231 0 2.0 1e-06 
0.0 1.2232 0 2.0 1e-06 
0.0 1.2233 0 2.0 1e-06 
0.0 1.2234 0 2.0 1e-06 
0.0 1.2235 0 2.0 1e-06 
0.0 1.2236 0 2.0 1e-06 
0.0 1.2237 0 2.0 1e-06 
0.0 1.2238 0 2.0 1e-06 
0.0 1.2239 0 2.0 1e-06 
0.0 1.224 0 2.0 1e-06 
0.0 1.2241 0 2.0 1e-06 
0.0 1.2242 0 2.0 1e-06 
0.0 1.2243 0 2.0 1e-06 
0.0 1.2244 0 2.0 1e-06 
0.0 1.2245 0 2.0 1e-06 
0.0 1.2246 0 2.0 1e-06 
0.0 1.2247 0 2.0 1e-06 
0.0 1.2248 0 2.0 1e-06 
0.0 1.2249 0 2.0 1e-06 
0.0 1.225 0 2.0 1e-06 
0.0 1.2251 0 2.0 1e-06 
0.0 1.2252 0 2.0 1e-06 
0.0 1.2253 0 2.0 1e-06 
0.0 1.2254 0 2.0 1e-06 
0.0 1.2255 0 2.0 1e-06 
0.0 1.2256 0 2.0 1e-06 
0.0 1.2257 0 2.0 1e-06 
0.0 1.2258 0 2.0 1e-06 
0.0 1.2259 0 2.0 1e-06 
0.0 1.226 0 2.0 1e-06 
0.0 1.2261 0 2.0 1e-06 
0.0 1.2262 0 2.0 1e-06 
0.0 1.2263 0 2.0 1e-06 
0.0 1.2264 0 2.0 1e-06 
0.0 1.2265 0 2.0 1e-06 
0.0 1.2266 0 2.0 1e-06 
0.0 1.2267 0 2.0 1e-06 
0.0 1.2268 0 2.0 1e-06 
0.0 1.2269 0 2.0 1e-06 
0.0 1.227 0 2.0 1e-06 
0.0 1.2271 0 2.0 1e-06 
0.0 1.2272 0 2.0 1e-06 
0.0 1.2273 0 2.0 1e-06 
0.0 1.2274 0 2.0 1e-06 
0.0 1.2275 0 2.0 1e-06 
0.0 1.2276 0 2.0 1e-06 
0.0 1.2277 0 2.0 1e-06 
0.0 1.2278 0 2.0 1e-06 
0.0 1.2279 0 2.0 1e-06 
0.0 1.228 0 2.0 1e-06 
0.0 1.2281 0 2.0 1e-06 
0.0 1.2282 0 2.0 1e-06 
0.0 1.2283 0 2.0 1e-06 
0.0 1.2284 0 2.0 1e-06 
0.0 1.2285 0 2.0 1e-06 
0.0 1.2286 0 2.0 1e-06 
0.0 1.2287 0 2.0 1e-06 
0.0 1.2288 0 2.0 1e-06 
0.0 1.2289 0 2.0 1e-06 
0.0 1.229 0 2.0 1e-06 
0.0 1.2291 0 2.0 1e-06 
0.0 1.2292 0 2.0 1e-06 
0.0 1.2293 0 2.0 1e-06 
0.0 1.2294 0 2.0 1e-06 
0.0 1.2295 0 2.0 1e-06 
0.0 1.2296 0 2.0 1e-06 
0.0 1.2297 0 2.0 1e-06 
0.0 1.2298 0 2.0 1e-06 
0.0 1.2299 0 2.0 1e-06 
0.0 1.23 0 2.0 1e-06 
0.0 1.2301 0 2.0 1e-06 
0.0 1.2302 0 2.0 1e-06 
0.0 1.2303 0 2.0 1e-06 
0.0 1.2304 0 2.0 1e-06 
0.0 1.2305 0 2.0 1e-06 
0.0 1.2306 0 2.0 1e-06 
0.0 1.2307 0 2.0 1e-06 
0.0 1.2308 0 2.0 1e-06 
0.0 1.2309 0 2.0 1e-06 
0.0 1.231 0 2.0 1e-06 
0.0 1.2311 0 2.0 1e-06 
0.0 1.2312 0 2.0 1e-06 
0.0 1.2313 0 2.0 1e-06 
0.0 1.2314 0 2.0 1e-06 
0.0 1.2315 0 2.0 1e-06 
0.0 1.2316 0 2.0 1e-06 
0.0 1.2317 0 2.0 1e-06 
0.0 1.2318 0 2.0 1e-06 
0.0 1.2319 0 2.0 1e-06 
0.0 1.232 0 2.0 1e-06 
0.0 1.2321 0 2.0 1e-06 
0.0 1.2322 0 2.0 1e-06 
0.0 1.2323 0 2.0 1e-06 
0.0 1.2324 0 2.0 1e-06 
0.0 1.2325 0 2.0 1e-06 
0.0 1.2326 0 2.0 1e-06 
0.0 1.2327 0 2.0 1e-06 
0.0 1.2328 0 2.0 1e-06 
0.0 1.2329 0 2.0 1e-06 
0.0 1.233 0 2.0 1e-06 
0.0 1.2331 0 2.0 1e-06 
0.0 1.2332 0 2.0 1e-06 
0.0 1.2333 0 2.0 1e-06 
0.0 1.2334 0 2.0 1e-06 
0.0 1.2335 0 2.0 1e-06 
0.0 1.2336 0 2.0 1e-06 
0.0 1.2337 0 2.0 1e-06 
0.0 1.2338 0 2.0 1e-06 
0.0 1.2339 0 2.0 1e-06 
0.0 1.234 0 2.0 1e-06 
0.0 1.2341 0 2.0 1e-06 
0.0 1.2342 0 2.0 1e-06 
0.0 1.2343 0 2.0 1e-06 
0.0 1.2344 0 2.0 1e-06 
0.0 1.2345 0 2.0 1e-06 
0.0 1.2346 0 2.0 1e-06 
0.0 1.2347 0 2.0 1e-06 
0.0 1.2348 0 2.0 1e-06 
0.0 1.2349 0 2.0 1e-06 
0.0 1.235 0 2.0 1e-06 
0.0 1.2351 0 2.0 1e-06 
0.0 1.2352 0 2.0 1e-06 
0.0 1.2353 0 2.0 1e-06 
0.0 1.2354 0 2.0 1e-06 
0.0 1.2355 0 2.0 1e-06 
0.0 1.2356 0 2.0 1e-06 
0.0 1.2357 0 2.0 1e-06 
0.0 1.2358 0 2.0 1e-06 
0.0 1.2359 0 2.0 1e-06 
0.0 1.236 0 2.0 1e-06 
0.0 1.2361 0 2.0 1e-06 
0.0 1.2362 0 2.0 1e-06 
0.0 1.2363 0 2.0 1e-06 
0.0 1.2364 0 2.0 1e-06 
0.0 1.2365 0 2.0 1e-06 
0.0 1.2366 0 2.0 1e-06 
0.0 1.2367 0 2.0 1e-06 
0.0 1.2368 0 2.0 1e-06 
0.0 1.2369 0 2.0 1e-06 
0.0 1.237 0 2.0 1e-06 
0.0 1.2371 0 2.0 1e-06 
0.0 1.2372 0 2.0 1e-06 
0.0 1.2373 0 2.0 1e-06 
0.0 1.2374 0 2.0 1e-06 
0.0 1.2375 0 2.0 1e-06 
0.0 1.2376 0 2.0 1e-06 
0.0 1.2377 0 2.0 1e-06 
0.0 1.2378 0 2.0 1e-06 
0.0 1.2379 0 2.0 1e-06 
0.0 1.238 0 2.0 1e-06 
0.0 1.2381 0 2.0 1e-06 
0.0 1.2382 0 2.0 1e-06 
0.0 1.2383 0 2.0 1e-06 
0.0 1.2384 0 2.0 1e-06 
0.0 1.2385 0 2.0 1e-06 
0.0 1.2386 0 2.0 1e-06 
0.0 1.2387 0 2.0 1e-06 
0.0 1.2388 0 2.0 1e-06 
0.0 1.2389 0 2.0 1e-06 
0.0 1.239 0 2.0 1e-06 
0.0 1.2391 0 2.0 1e-06 
0.0 1.2392 0 2.0 1e-06 
0.0 1.2393 0 2.0 1e-06 
0.0 1.2394 0 2.0 1e-06 
0.0 1.2395 0 2.0 1e-06 
0.0 1.2396 0 2.0 1e-06 
0.0 1.2397 0 2.0 1e-06 
0.0 1.2398 0 2.0 1e-06 
0.0 1.2399 0 2.0 1e-06 
0.0 1.24 0 2.0 1e-06 
0.0 1.2401 0 2.0 1e-06 
0.0 1.2402 0 2.0 1e-06 
0.0 1.2403 0 2.0 1e-06 
0.0 1.2404 0 2.0 1e-06 
0.0 1.2405 0 2.0 1e-06 
0.0 1.2406 0 2.0 1e-06 
0.0 1.2407 0 2.0 1e-06 
0.0 1.2408 0 2.0 1e-06 
0.0 1.2409 0 2.0 1e-06 
0.0 1.241 0 2.0 1e-06 
0.0 1.2411 0 2.0 1e-06 
0.0 1.2412 0 2.0 1e-06 
0.0 1.2413 0 2.0 1e-06 
0.0 1.2414 0 2.0 1e-06 
0.0 1.2415 0 2.0 1e-06 
0.0 1.2416 0 2.0 1e-06 
0.0 1.2417 0 2.0 1e-06 
0.0 1.2418 0 2.0 1e-06 
0.0 1.2419 0 2.0 1e-06 
0.0 1.242 0 2.0 1e-06 
0.0 1.2421 0 2.0 1e-06 
0.0 1.2422 0 2.0 1e-06 
0.0 1.2423 0 2.0 1e-06 
0.0 1.2424 0 2.0 1e-06 
0.0 1.2425 0 2.0 1e-06 
0.0 1.2426 0 2.0 1e-06 
0.0 1.2427 0 2.0 1e-06 
0.0 1.2428 0 2.0 1e-06 
0.0 1.2429 0 2.0 1e-06 
0.0 1.243 0 2.0 1e-06 
0.0 1.2431 0 2.0 1e-06 
0.0 1.2432 0 2.0 1e-06 
0.0 1.2433 0 2.0 1e-06 
0.0 1.2434 0 2.0 1e-06 
0.0 1.2435 0 2.0 1e-06 
0.0 1.2436 0 2.0 1e-06 
0.0 1.2437 0 2.0 1e-06 
0.0 1.2438 0 2.0 1e-06 
0.0 1.2439 0 2.0 1e-06 
0.0 1.244 0 2.0 1e-06 
0.0 1.2441 0 2.0 1e-06 
0.0 1.2442 0 2.0 1e-06 
0.0 1.2443 0 2.0 1e-06 
0.0 1.2444 0 2.0 1e-06 
0.0 1.2445 0 2.0 1e-06 
0.0 1.2446 0 2.0 1e-06 
0.0 1.2447 0 2.0 1e-06 
0.0 1.2448 0 2.0 1e-06 
0.0 1.2449 0 2.0 1e-06 
0.0 1.245 0 2.0 1e-06 
0.0 1.2451 0 2.0 1e-06 
0.0 1.2452 0 2.0 1e-06 
0.0 1.2453 0 2.0 1e-06 
0.0 1.2454 0 2.0 1e-06 
0.0 1.2455 0 2.0 1e-06 
0.0 1.2456 0 2.0 1e-06 
0.0 1.2457 0 2.0 1e-06 
0.0 1.2458 0 2.0 1e-06 
0.0 1.2459 0 2.0 1e-06 
0.0 1.246 0 2.0 1e-06 
0.0 1.2461 0 2.0 1e-06 
0.0 1.2462 0 2.0 1e-06 
0.0 1.2463 0 2.0 1e-06 
0.0 1.2464 0 2.0 1e-06 
0.0 1.2465 0 2.0 1e-06 
0.0 1.2466 0 2.0 1e-06 
0.0 1.2467 0 2.0 1e-06 
0.0 1.2468 0 2.0 1e-06 
0.0 1.2469 0 2.0 1e-06 
0.0 1.247 0 2.0 1e-06 
0.0 1.2471 0 2.0 1e-06 
0.0 1.2472 0 2.0 1e-06 
0.0 1.2473 0 2.0 1e-06 
0.0 1.2474 0 2.0 1e-06 
0.0 1.2475 0 2.0 1e-06 
0.0 1.2476 0 2.0 1e-06 
0.0 1.2477 0 2.0 1e-06 
0.0 1.2478 0 2.0 1e-06 
0.0 1.2479 0 2.0 1e-06 
0.0 1.248 0 2.0 1e-06 
0.0 1.2481 0 2.0 1e-06 
0.0 1.2482 0 2.0 1e-06 
0.0 1.2483 0 2.0 1e-06 
0.0 1.2484 0 2.0 1e-06 
0.0 1.2485 0 2.0 1e-06 
0.0 1.2486 0 2.0 1e-06 
0.0 1.2487 0 2.0 1e-06 
0.0 1.2488 0 2.0 1e-06 
0.0 1.2489 0 2.0 1e-06 
0.0 1.249 0 2.0 1e-06 
0.0 1.2491 0 2.0 1e-06 
0.0 1.2492 0 2.0 1e-06 
0.0 1.2493 0 2.0 1e-06 
0.0 1.2494 0 2.0 1e-06 
0.0 1.2495 0 2.0 1e-06 
0.0 1.2496 0 2.0 1e-06 
0.0 1.2497 0 2.0 1e-06 
0.0 1.2498 0 2.0 1e-06 
0.0 1.2499 0 2.0 1e-06 
0.0 1.25 0 2.0 1e-06 
0.0 1.2501 0 2.0 1e-06 
0.0 1.2502 0 2.0 1e-06 
0.0 1.2503 0 2.0 1e-06 
0.0 1.2504 0 2.0 1e-06 
0.0 1.2505 0 2.0 1e-06 
0.0 1.2506 0 2.0 1e-06 
0.0 1.2507 0 2.0 1e-06 
0.0 1.2508 0 2.0 1e-06 
0.0 1.2509 0 2.0 1e-06 
0.0 1.251 0 2.0 1e-06 
0.0 1.2511 0 2.0 1e-06 
0.0 1.2512 0 2.0 1e-06 
0.0 1.2513 0 2.0 1e-06 
0.0 1.2514 0 2.0 1e-06 
0.0 1.2515 0 2.0 1e-06 
0.0 1.2516 0 2.0 1e-06 
0.0 1.2517 0 2.0 1e-06 
0.0 1.2518 0 2.0 1e-06 
0.0 1.2519 0 2.0 1e-06 
0.0 1.252 0 2.0 1e-06 
0.0 1.2521 0 2.0 1e-06 
0.0 1.2522 0 2.0 1e-06 
0.0 1.2523 0 2.0 1e-06 
0.0 1.2524 0 2.0 1e-06 
0.0 1.2525 0 2.0 1e-06 
0.0 1.2526 0 2.0 1e-06 
0.0 1.2527 0 2.0 1e-06 
0.0 1.2528 0 2.0 1e-06 
0.0 1.2529 0 2.0 1e-06 
0.0 1.253 0 2.0 1e-06 
0.0 1.2531 0 2.0 1e-06 
0.0 1.2532 0 2.0 1e-06 
0.0 1.2533 0 2.0 1e-06 
0.0 1.2534 0 2.0 1e-06 
0.0 1.2535 0 2.0 1e-06 
0.0 1.2536 0 2.0 1e-06 
0.0 1.2537 0 2.0 1e-06 
0.0 1.2538 0 2.0 1e-06 
0.0 1.2539 0 2.0 1e-06 
0.0 1.254 0 2.0 1e-06 
0.0 1.2541 0 2.0 1e-06 
0.0 1.2542 0 2.0 1e-06 
0.0 1.2543 0 2.0 1e-06 
0.0 1.2544 0 2.0 1e-06 
0.0 1.2545 0 2.0 1e-06 
0.0 1.2546 0 2.0 1e-06 
0.0 1.2547 0 2.0 1e-06 
0.0 1.2548 0 2.0 1e-06 
0.0 1.2549 0 2.0 1e-06 
0.0 1.255 0 2.0 1e-06 
0.0 1.2551 0 2.0 1e-06 
0.0 1.2552 0 2.0 1e-06 
0.0 1.2553 0 2.0 1e-06 
0.0 1.2554 0 2.0 1e-06 
0.0 1.2555 0 2.0 1e-06 
0.0 1.2556 0 2.0 1e-06 
0.0 1.2557 0 2.0 1e-06 
0.0 1.2558 0 2.0 1e-06 
0.0 1.2559 0 2.0 1e-06 
0.0 1.256 0 2.0 1e-06 
0.0 1.2561 0 2.0 1e-06 
0.0 1.2562 0 2.0 1e-06 
0.0 1.2563 0 2.0 1e-06 
0.0 1.2564 0 2.0 1e-06 
0.0 1.2565 0 2.0 1e-06 
0.0 1.2566 0 2.0 1e-06 
0.0 1.2567 0 2.0 1e-06 
0.0 1.2568 0 2.0 1e-06 
0.0 1.2569 0 2.0 1e-06 
0.0 1.257 0 2.0 1e-06 
0.0 1.2571 0 2.0 1e-06 
0.0 1.2572 0 2.0 1e-06 
0.0 1.2573 0 2.0 1e-06 
0.0 1.2574 0 2.0 1e-06 
0.0 1.2575 0 2.0 1e-06 
0.0 1.2576 0 2.0 1e-06 
0.0 1.2577 0 2.0 1e-06 
0.0 1.2578 0 2.0 1e-06 
0.0 1.2579 0 2.0 1e-06 
0.0 1.258 0 2.0 1e-06 
0.0 1.2581 0 2.0 1e-06 
0.0 1.2582 0 2.0 1e-06 
0.0 1.2583 0 2.0 1e-06 
0.0 1.2584 0 2.0 1e-06 
0.0 1.2585 0 2.0 1e-06 
0.0 1.2586 0 2.0 1e-06 
0.0 1.2587 0 2.0 1e-06 
0.0 1.2588 0 2.0 1e-06 
0.0 1.2589 0 2.0 1e-06 
0.0 1.259 0 2.0 1e-06 
0.0 1.2591 0 2.0 1e-06 
0.0 1.2592 0 2.0 1e-06 
0.0 1.2593 0 2.0 1e-06 
0.0 1.2594 0 2.0 1e-06 
0.0 1.2595 0 2.0 1e-06 
0.0 1.2596 0 2.0 1e-06 
0.0 1.2597 0 2.0 1e-06 
0.0 1.2598 0 2.0 1e-06 
0.0 1.2599 0 2.0 1e-06 
0.0 1.26 0 2.0 1e-06 
0.0 1.2601 0 2.0 1e-06 
0.0 1.2602 0 2.0 1e-06 
0.0 1.2603 0 2.0 1e-06 
0.0 1.2604 0 2.0 1e-06 
0.0 1.2605 0 2.0 1e-06 
0.0 1.2606 0 2.0 1e-06 
0.0 1.2607 0 2.0 1e-06 
0.0 1.2608 0 2.0 1e-06 
0.0 1.2609 0 2.0 1e-06 
0.0 1.261 0 2.0 1e-06 
0.0 1.2611 0 2.0 1e-06 
0.0 1.2612 0 2.0 1e-06 
0.0 1.2613 0 2.0 1e-06 
0.0 1.2614 0 2.0 1e-06 
0.0 1.2615 0 2.0 1e-06 
0.0 1.2616 0 2.0 1e-06 
0.0 1.2617 0 2.0 1e-06 
0.0 1.2618 0 2.0 1e-06 
0.0 1.2619 0 2.0 1e-06 
0.0 1.262 0 2.0 1e-06 
0.0 1.2621 0 2.0 1e-06 
0.0 1.2622 0 2.0 1e-06 
0.0 1.2623 0 2.0 1e-06 
0.0 1.2624 0 2.0 1e-06 
0.0 1.2625 0 2.0 1e-06 
0.0 1.2626 0 2.0 1e-06 
0.0 1.2627 0 2.0 1e-06 
0.0 1.2628 0 2.0 1e-06 
0.0 1.2629 0 2.0 1e-06 
0.0 1.263 0 2.0 1e-06 
0.0 1.2631 0 2.0 1e-06 
0.0 1.2632 0 2.0 1e-06 
0.0 1.2633 0 2.0 1e-06 
0.0 1.2634 0 2.0 1e-06 
0.0 1.2635 0 2.0 1e-06 
0.0 1.2636 0 2.0 1e-06 
0.0 1.2637 0 2.0 1e-06 
0.0 1.2638 0 2.0 1e-06 
0.0 1.2639 0 2.0 1e-06 
0.0 1.264 0 2.0 1e-06 
0.0 1.2641 0 2.0 1e-06 
0.0 1.2642 0 2.0 1e-06 
0.0 1.2643 0 2.0 1e-06 
0.0 1.2644 0 2.0 1e-06 
0.0 1.2645 0 2.0 1e-06 
0.0 1.2646 0 2.0 1e-06 
0.0 1.2647 0 2.0 1e-06 
0.0 1.2648 0 2.0 1e-06 
0.0 1.2649 0 2.0 1e-06 
0.0 1.265 0 2.0 1e-06 
0.0 1.2651 0 2.0 1e-06 
0.0 1.2652 0 2.0 1e-06 
0.0 1.2653 0 2.0 1e-06 
0.0 1.2654 0 2.0 1e-06 
0.0 1.2655 0 2.0 1e-06 
0.0 1.2656 0 2.0 1e-06 
0.0 1.2657 0 2.0 1e-06 
0.0 1.2658 0 2.0 1e-06 
0.0 1.2659 0 2.0 1e-06 
0.0 1.266 0 2.0 1e-06 
0.0 1.2661 0 2.0 1e-06 
0.0 1.2662 0 2.0 1e-06 
0.0 1.2663 0 2.0 1e-06 
0.0 1.2664 0 2.0 1e-06 
0.0 1.2665 0 2.0 1e-06 
0.0 1.2666 0 2.0 1e-06 
0.0 1.2667 0 2.0 1e-06 
0.0 1.2668 0 2.0 1e-06 
0.0 1.2669 0 2.0 1e-06 
0.0 1.267 0 2.0 1e-06 
0.0 1.2671 0 2.0 1e-06 
0.0 1.2672 0 2.0 1e-06 
0.0 1.2673 0 2.0 1e-06 
0.0 1.2674 0 2.0 1e-06 
0.0 1.2675 0 2.0 1e-06 
0.0 1.2676 0 2.0 1e-06 
0.0 1.2677 0 2.0 1e-06 
0.0 1.2678 0 2.0 1e-06 
0.0 1.2679 0 2.0 1e-06 
0.0 1.268 0 2.0 1e-06 
0.0 1.2681 0 2.0 1e-06 
0.0 1.2682 0 2.0 1e-06 
0.0 1.2683 0 2.0 1e-06 
0.0 1.2684 0 2.0 1e-06 
0.0 1.2685 0 2.0 1e-06 
0.0 1.2686 0 2.0 1e-06 
0.0 1.2687 0 2.0 1e-06 
0.0 1.2688 0 2.0 1e-06 
0.0 1.2689 0 2.0 1e-06 
0.0 1.269 0 2.0 1e-06 
0.0 1.2691 0 2.0 1e-06 
0.0 1.2692 0 2.0 1e-06 
0.0 1.2693 0 2.0 1e-06 
0.0 1.2694 0 2.0 1e-06 
0.0 1.2695 0 2.0 1e-06 
0.0 1.2696 0 2.0 1e-06 
0.0 1.2697 0 2.0 1e-06 
0.0 1.2698 0 2.0 1e-06 
0.0 1.2699 0 2.0 1e-06 
0.0 1.27 0 2.0 1e-06 
0.0 1.2701 0 2.0 1e-06 
0.0 1.2702 0 2.0 1e-06 
0.0 1.2703 0 2.0 1e-06 
0.0 1.2704 0 2.0 1e-06 
0.0 1.2705 0 2.0 1e-06 
0.0 1.2706 0 2.0 1e-06 
0.0 1.2707 0 2.0 1e-06 
0.0 1.2708 0 2.0 1e-06 
0.0 1.2709 0 2.0 1e-06 
0.0 1.271 0 2.0 1e-06 
0.0 1.2711 0 2.0 1e-06 
0.0 1.2712 0 2.0 1e-06 
0.0 1.2713 0 2.0 1e-06 
0.0 1.2714 0 2.0 1e-06 
0.0 1.2715 0 2.0 1e-06 
0.0 1.2716 0 2.0 1e-06 
0.0 1.2717 0 2.0 1e-06 
0.0 1.2718 0 2.0 1e-06 
0.0 1.2719 0 2.0 1e-06 
0.0 1.272 0 2.0 1e-06 
0.0 1.2721 0 2.0 1e-06 
0.0 1.2722 0 2.0 1e-06 
0.0 1.2723 0 2.0 1e-06 
0.0 1.2724 0 2.0 1e-06 
0.0 1.2725 0 2.0 1e-06 
0.0 1.2726 0 2.0 1e-06 
0.0 1.2727 0 2.0 1e-06 
0.0 1.2728 0 2.0 1e-06 
0.0 1.2729 0 2.0 1e-06 
0.0 1.273 0 2.0 1e-06 
0.0 1.2731 0 2.0 1e-06 
0.0 1.2732 0 2.0 1e-06 
0.0 1.2733 0 2.0 1e-06 
0.0 1.2734 0 2.0 1e-06 
0.0 1.2735 0 2.0 1e-06 
0.0 1.2736 0 2.0 1e-06 
0.0 1.2737 0 2.0 1e-06 
0.0 1.2738 0 2.0 1e-06 
0.0 1.2739 0 2.0 1e-06 
0.0 1.274 0 2.0 1e-06 
0.0 1.2741 0 2.0 1e-06 
0.0 1.2742 0 2.0 1e-06 
0.0 1.2743 0 2.0 1e-06 
0.0 1.2744 0 2.0 1e-06 
0.0 1.2745 0 2.0 1e-06 
0.0 1.2746 0 2.0 1e-06 
0.0 1.2747 0 2.0 1e-06 
0.0 1.2748 0 2.0 1e-06 
0.0 1.2749 0 2.0 1e-06 
0.0 1.275 0 2.0 1e-06 
0.0 1.2751 0 2.0 1e-06 
0.0 1.2752 0 2.0 1e-06 
0.0 1.2753 0 2.0 1e-06 
0.0 1.2754 0 2.0 1e-06 
0.0 1.2755 0 2.0 1e-06 
0.0 1.2756 0 2.0 1e-06 
0.0 1.2757 0 2.0 1e-06 
0.0 1.2758 0 2.0 1e-06 
0.0 1.2759 0 2.0 1e-06 
0.0 1.276 0 2.0 1e-06 
0.0 1.2761 0 2.0 1e-06 
0.0 1.2762 0 2.0 1e-06 
0.0 1.2763 0 2.0 1e-06 
0.0 1.2764 0 2.0 1e-06 
0.0 1.2765 0 2.0 1e-06 
0.0 1.2766 0 2.0 1e-06 
0.0 1.2767 0 2.0 1e-06 
0.0 1.2768 0 2.0 1e-06 
0.0 1.2769 0 2.0 1e-06 
0.0 1.277 0 2.0 1e-06 
0.0 1.2771 0 2.0 1e-06 
0.0 1.2772 0 2.0 1e-06 
0.0 1.2773 0 2.0 1e-06 
0.0 1.2774 0 2.0 1e-06 
0.0 1.2775 0 2.0 1e-06 
0.0 1.2776 0 2.0 1e-06 
0.0 1.2777 0 2.0 1e-06 
0.0 1.2778 0 2.0 1e-06 
0.0 1.2779 0 2.0 1e-06 
0.0 1.278 0 2.0 1e-06 
0.0 1.2781 0 2.0 1e-06 
0.0 1.2782 0 2.0 1e-06 
0.0 1.2783 0 2.0 1e-06 
0.0 1.2784 0 2.0 1e-06 
0.0 1.2785 0 2.0 1e-06 
0.0 1.2786 0 2.0 1e-06 
0.0 1.2787 0 2.0 1e-06 
0.0 1.2788 0 2.0 1e-06 
0.0 1.2789 0 2.0 1e-06 
0.0 1.279 0 2.0 1e-06 
0.0 1.2791 0 2.0 1e-06 
0.0 1.2792 0 2.0 1e-06 
0.0 1.2793 0 2.0 1e-06 
0.0 1.2794 0 2.0 1e-06 
0.0 1.2795 0 2.0 1e-06 
0.0 1.2796 0 2.0 1e-06 
0.0 1.2797 0 2.0 1e-06 
0.0 1.2798 0 2.0 1e-06 
0.0 1.2799 0 2.0 1e-06 
0.0 1.28 0 2.0 1e-06 
0.0 1.2801 0 2.0 1e-06 
0.0 1.2802 0 2.0 1e-06 
0.0 1.2803 0 2.0 1e-06 
0.0 1.2804 0 2.0 1e-06 
0.0 1.2805 0 2.0 1e-06 
0.0 1.2806 0 2.0 1e-06 
0.0 1.2807 0 2.0 1e-06 
0.0 1.2808 0 2.0 1e-06 
0.0 1.2809 0 2.0 1e-06 
0.0 1.281 0 2.0 1e-06 
0.0 1.2811 0 2.0 1e-06 
0.0 1.2812 0 2.0 1e-06 
0.0 1.2813 0 2.0 1e-06 
0.0 1.2814 0 2.0 1e-06 
0.0 1.2815 0 2.0 1e-06 
0.0 1.2816 0 2.0 1e-06 
0.0 1.2817 0 2.0 1e-06 
0.0 1.2818 0 2.0 1e-06 
0.0 1.2819 0 2.0 1e-06 
0.0 1.282 0 2.0 1e-06 
0.0 1.2821 0 2.0 1e-06 
0.0 1.2822 0 2.0 1e-06 
0.0 1.2823 0 2.0 1e-06 
0.0 1.2824 0 2.0 1e-06 
0.0 1.2825 0 2.0 1e-06 
0.0 1.2826 0 2.0 1e-06 
0.0 1.2827 0 2.0 1e-06 
0.0 1.2828 0 2.0 1e-06 
0.0 1.2829 0 2.0 1e-06 
0.0 1.283 0 2.0 1e-06 
0.0 1.2831 0 2.0 1e-06 
0.0 1.2832 0 2.0 1e-06 
0.0 1.2833 0 2.0 1e-06 
0.0 1.2834 0 2.0 1e-06 
0.0 1.2835 0 2.0 1e-06 
0.0 1.2836 0 2.0 1e-06 
0.0 1.2837 0 2.0 1e-06 
0.0 1.2838 0 2.0 1e-06 
0.0 1.2839 0 2.0 1e-06 
0.0 1.284 0 2.0 1e-06 
0.0 1.2841 0 2.0 1e-06 
0.0 1.2842 0 2.0 1e-06 
0.0 1.2843 0 2.0 1e-06 
0.0 1.2844 0 2.0 1e-06 
0.0 1.2845 0 2.0 1e-06 
0.0 1.2846 0 2.0 1e-06 
0.0 1.2847 0 2.0 1e-06 
0.0 1.2848 0 2.0 1e-06 
0.0 1.2849 0 2.0 1e-06 
0.0 1.285 0 2.0 1e-06 
0.0 1.2851 0 2.0 1e-06 
0.0 1.2852 0 2.0 1e-06 
0.0 1.2853 0 2.0 1e-06 
0.0 1.2854 0 2.0 1e-06 
0.0 1.2855 0 2.0 1e-06 
0.0 1.2856 0 2.0 1e-06 
0.0 1.2857 0 2.0 1e-06 
0.0 1.2858 0 2.0 1e-06 
0.0 1.2859 0 2.0 1e-06 
0.0 1.286 0 2.0 1e-06 
0.0 1.2861 0 2.0 1e-06 
0.0 1.2862 0 2.0 1e-06 
0.0 1.2863 0 2.0 1e-06 
0.0 1.2864 0 2.0 1e-06 
0.0 1.2865 0 2.0 1e-06 
0.0 1.2866 0 2.0 1e-06 
0.0 1.2867 0 2.0 1e-06 
0.0 1.2868 0 2.0 1e-06 
0.0 1.2869 0 2.0 1e-06 
0.0 1.287 0 2.0 1e-06 
0.0 1.2871 0 2.0 1e-06 
0.0 1.2872 0 2.0 1e-06 
0.0 1.2873 0 2.0 1e-06 
0.0 1.2874 0 2.0 1e-06 
0.0 1.2875 0 2.0 1e-06 
0.0 1.2876 0 2.0 1e-06 
0.0 1.2877 0 2.0 1e-06 
0.0 1.2878 0 2.0 1e-06 
0.0 1.2879 0 2.0 1e-06 
0.0 1.288 0 2.0 1e-06 
0.0 1.2881 0 2.0 1e-06 
0.0 1.2882 0 2.0 1e-06 
0.0 1.2883 0 2.0 1e-06 
0.0 1.2884 0 2.0 1e-06 
0.0 1.2885 0 2.0 1e-06 
0.0 1.2886 0 2.0 1e-06 
0.0 1.2887 0 2.0 1e-06 
0.0 1.2888 0 2.0 1e-06 
0.0 1.2889 0 2.0 1e-06 
0.0 1.289 0 2.0 1e-06 
0.0 1.2891 0 2.0 1e-06 
0.0 1.2892 0 2.0 1e-06 
0.0 1.2893 0 2.0 1e-06 
0.0 1.2894 0 2.0 1e-06 
0.0 1.2895 0 2.0 1e-06 
0.0 1.2896 0 2.0 1e-06 
0.0 1.2897 0 2.0 1e-06 
0.0 1.2898 0 2.0 1e-06 
0.0 1.2899 0 2.0 1e-06 
0.0 1.29 0 2.0 1e-06 
0.0 1.2901 0 2.0 1e-06 
0.0 1.2902 0 2.0 1e-06 
0.0 1.2903 0 2.0 1e-06 
0.0 1.2904 0 2.0 1e-06 
0.0 1.2905 0 2.0 1e-06 
0.0 1.2906 0 2.0 1e-06 
0.0 1.2907 0 2.0 1e-06 
0.0 1.2908 0 2.0 1e-06 
0.0 1.2909 0 2.0 1e-06 
0.0 1.291 0 2.0 1e-06 
0.0 1.2911 0 2.0 1e-06 
0.0 1.2912 0 2.0 1e-06 
0.0 1.2913 0 2.0 1e-06 
0.0 1.2914 0 2.0 1e-06 
0.0 1.2915 0 2.0 1e-06 
0.0 1.2916 0 2.0 1e-06 
0.0 1.2917 0 2.0 1e-06 
0.0 1.2918 0 2.0 1e-06 
0.0 1.2919 0 2.0 1e-06 
0.0 1.292 0 2.0 1e-06 
0.0 1.2921 0 2.0 1e-06 
0.0 1.2922 0 2.0 1e-06 
0.0 1.2923 0 2.0 1e-06 
0.0 1.2924 0 2.0 1e-06 
0.0 1.2925 0 2.0 1e-06 
0.0 1.2926 0 2.0 1e-06 
0.0 1.2927 0 2.0 1e-06 
0.0 1.2928 0 2.0 1e-06 
0.0 1.2929 0 2.0 1e-06 
0.0 1.293 0 2.0 1e-06 
0.0 1.2931 0 2.0 1e-06 
0.0 1.2932 0 2.0 1e-06 
0.0 1.2933 0 2.0 1e-06 
0.0 1.2934 0 2.0 1e-06 
0.0 1.2935 0 2.0 1e-06 
0.0 1.2936 0 2.0 1e-06 
0.0 1.2937 0 2.0 1e-06 
0.0 1.2938 0 2.0 1e-06 
0.0 1.2939 0 2.0 1e-06 
0.0 1.294 0 2.0 1e-06 
0.0 1.2941 0 2.0 1e-06 
0.0 1.2942 0 2.0 1e-06 
0.0 1.2943 0 2.0 1e-06 
0.0 1.2944 0 2.0 1e-06 
0.0 1.2945 0 2.0 1e-06 
0.0 1.2946 0 2.0 1e-06 
0.0 1.2947 0 2.0 1e-06 
0.0 1.2948 0 2.0 1e-06 
0.0 1.2949 0 2.0 1e-06 
0.0 1.295 0 2.0 1e-06 
0.0 1.2951 0 2.0 1e-06 
0.0 1.2952 0 2.0 1e-06 
0.0 1.2953 0 2.0 1e-06 
0.0 1.2954 0 2.0 1e-06 
0.0 1.2955 0 2.0 1e-06 
0.0 1.2956 0 2.0 1e-06 
0.0 1.2957 0 2.0 1e-06 
0.0 1.2958 0 2.0 1e-06 
0.0 1.2959 0 2.0 1e-06 
0.0 1.296 0 2.0 1e-06 
0.0 1.2961 0 2.0 1e-06 
0.0 1.2962 0 2.0 1e-06 
0.0 1.2963 0 2.0 1e-06 
0.0 1.2964 0 2.0 1e-06 
0.0 1.2965 0 2.0 1e-06 
0.0 1.2966 0 2.0 1e-06 
0.0 1.2967 0 2.0 1e-06 
0.0 1.2968 0 2.0 1e-06 
0.0 1.2969 0 2.0 1e-06 
0.0 1.297 0 2.0 1e-06 
0.0 1.2971 0 2.0 1e-06 
0.0 1.2972 0 2.0 1e-06 
0.0 1.2973 0 2.0 1e-06 
0.0 1.2974 0 2.0 1e-06 
0.0 1.2975 0 2.0 1e-06 
0.0 1.2976 0 2.0 1e-06 
0.0 1.2977 0 2.0 1e-06 
0.0 1.2978 0 2.0 1e-06 
0.0 1.2979 0 2.0 1e-06 
0.0 1.298 0 2.0 1e-06 
0.0 1.2981 0 2.0 1e-06 
0.0 1.2982 0 2.0 1e-06 
0.0 1.2983 0 2.0 1e-06 
0.0 1.2984 0 2.0 1e-06 
0.0 1.2985 0 2.0 1e-06 
0.0 1.2986 0 2.0 1e-06 
0.0 1.2987 0 2.0 1e-06 
0.0 1.2988 0 2.0 1e-06 
0.0 1.2989 0 2.0 1e-06 
0.0 1.299 0 2.0 1e-06 
0.0 1.2991 0 2.0 1e-06 
0.0 1.2992 0 2.0 1e-06 
0.0 1.2993 0 2.0 1e-06 
0.0 1.2994 0 2.0 1e-06 
0.0 1.2995 0 2.0 1e-06 
0.0 1.2996 0 2.0 1e-06 
0.0 1.2997 0 2.0 1e-06 
0.0 1.2998 0 2.0 1e-06 
0.0 1.2999 0 2.0 1e-06 
0.0 1.3 0 2.0 1e-06 
0.0 1.3001 0 2.0 1e-06 
0.0 1.3002 0 2.0 1e-06 
0.0 1.3003 0 2.0 1e-06 
0.0 1.3004 0 2.0 1e-06 
0.0 1.3005 0 2.0 1e-06 
0.0 1.3006 0 2.0 1e-06 
0.0 1.3007 0 2.0 1e-06 
0.0 1.3008 0 2.0 1e-06 
0.0 1.3009 0 2.0 1e-06 
0.0 1.301 0 2.0 1e-06 
0.0 1.3011 0 2.0 1e-06 
0.0 1.3012 0 2.0 1e-06 
0.0 1.3013 0 2.0 1e-06 
0.0 1.3014 0 2.0 1e-06 
0.0 1.3015 0 2.0 1e-06 
0.0 1.3016 0 2.0 1e-06 
0.0 1.3017 0 2.0 1e-06 
0.0 1.3018 0 2.0 1e-06 
0.0 1.3019 0 2.0 1e-06 
0.0 1.302 0 2.0 1e-06 
0.0 1.3021 0 2.0 1e-06 
0.0 1.3022 0 2.0 1e-06 
0.0 1.3023 0 2.0 1e-06 
0.0 1.3024 0 2.0 1e-06 
0.0 1.3025 0 2.0 1e-06 
0.0 1.3026 0 2.0 1e-06 
0.0 1.3027 0 2.0 1e-06 
0.0 1.3028 0 2.0 1e-06 
0.0 1.3029 0 2.0 1e-06 
0.0 1.303 0 2.0 1e-06 
0.0 1.3031 0 2.0 1e-06 
0.0 1.3032 0 2.0 1e-06 
0.0 1.3033 0 2.0 1e-06 
0.0 1.3034 0 2.0 1e-06 
0.0 1.3035 0 2.0 1e-06 
0.0 1.3036 0 2.0 1e-06 
0.0 1.3037 0 2.0 1e-06 
0.0 1.3038 0 2.0 1e-06 
0.0 1.3039 0 2.0 1e-06 
0.0 1.304 0 2.0 1e-06 
0.0 1.3041 0 2.0 1e-06 
0.0 1.3042 0 2.0 1e-06 
0.0 1.3043 0 2.0 1e-06 
0.0 1.3044 0 2.0 1e-06 
0.0 1.3045 0 2.0 1e-06 
0.0 1.3046 0 2.0 1e-06 
0.0 1.3047 0 2.0 1e-06 
0.0 1.3048 0 2.0 1e-06 
0.0 1.3049 0 2.0 1e-06 
0.0 1.305 0 2.0 1e-06 
0.0 1.3051 0 2.0 1e-06 
0.0 1.3052 0 2.0 1e-06 
0.0 1.3053 0 2.0 1e-06 
0.0 1.3054 0 2.0 1e-06 
0.0 1.3055 0 2.0 1e-06 
0.0 1.3056 0 2.0 1e-06 
0.0 1.3057 0 2.0 1e-06 
0.0 1.3058 0 2.0 1e-06 
0.0 1.3059 0 2.0 1e-06 
0.0 1.306 0 2.0 1e-06 
0.0 1.3061 0 2.0 1e-06 
0.0 1.3062 0 2.0 1e-06 
0.0 1.3063 0 2.0 1e-06 
0.0 1.3064 0 2.0 1e-06 
0.0 1.3065 0 2.0 1e-06 
0.0 1.3066 0 2.0 1e-06 
0.0 1.3067 0 2.0 1e-06 
0.0 1.3068 0 2.0 1e-06 
0.0 1.3069 0 2.0 1e-06 
0.0 1.307 0 2.0 1e-06 
0.0 1.3071 0 2.0 1e-06 
0.0 1.3072 0 2.0 1e-06 
0.0 1.3073 0 2.0 1e-06 
0.0 1.3074 0 2.0 1e-06 
0.0 1.3075 0 2.0 1e-06 
0.0 1.3076 0 2.0 1e-06 
0.0 1.3077 0 2.0 1e-06 
0.0 1.3078 0 2.0 1e-06 
0.0 1.3079 0 2.0 1e-06 
0.0 1.308 0 2.0 1e-06 
0.0 1.3081 0 2.0 1e-06 
0.0 1.3082 0 2.0 1e-06 
0.0 1.3083 0 2.0 1e-06 
0.0 1.3084 0 2.0 1e-06 
0.0 1.3085 0 2.0 1e-06 
0.0 1.3086 0 2.0 1e-06 
0.0 1.3087 0 2.0 1e-06 
0.0 1.3088 0 2.0 1e-06 
0.0 1.3089 0 2.0 1e-06 
0.0 1.309 0 2.0 1e-06 
0.0 1.3091 0 2.0 1e-06 
0.0 1.3092 0 2.0 1e-06 
0.0 1.3093 0 2.0 1e-06 
0.0 1.3094 0 2.0 1e-06 
0.0 1.3095 0 2.0 1e-06 
0.0 1.3096 0 2.0 1e-06 
0.0 1.3097 0 2.0 1e-06 
0.0 1.3098 0 2.0 1e-06 
0.0 1.3099 0 2.0 1e-06 
0.0 1.31 0 2.0 1e-06 
0.0 1.3101 0 2.0 1e-06 
0.0 1.3102 0 2.0 1e-06 
0.0 1.3103 0 2.0 1e-06 
0.0 1.3104 0 2.0 1e-06 
0.0 1.3105 0 2.0 1e-06 
0.0 1.3106 0 2.0 1e-06 
0.0 1.3107 0 2.0 1e-06 
0.0 1.3108 0 2.0 1e-06 
0.0 1.3109 0 2.0 1e-06 
0.0 1.311 0 2.0 1e-06 
0.0 1.3111 0 2.0 1e-06 
0.0 1.3112 0 2.0 1e-06 
0.0 1.3113 0 2.0 1e-06 
0.0 1.3114 0 2.0 1e-06 
0.0 1.3115 0 2.0 1e-06 
0.0 1.3116 0 2.0 1e-06 
0.0 1.3117 0 2.0 1e-06 
0.0 1.3118 0 2.0 1e-06 
0.0 1.3119 0 2.0 1e-06 
0.0 1.312 0 2.0 1e-06 
0.0 1.3121 0 2.0 1e-06 
0.0 1.3122 0 2.0 1e-06 
0.0 1.3123 0 2.0 1e-06 
0.0 1.3124 0 2.0 1e-06 
0.0 1.3125 0 2.0 1e-06 
0.0 1.3126 0 2.0 1e-06 
0.0 1.3127 0 2.0 1e-06 
0.0 1.3128 0 2.0 1e-06 
0.0 1.3129 0 2.0 1e-06 
0.0 1.313 0 2.0 1e-06 
0.0 1.3131 0 2.0 1e-06 
0.0 1.3132 0 2.0 1e-06 
0.0 1.3133 0 2.0 1e-06 
0.0 1.3134 0 2.0 1e-06 
0.0 1.3135 0 2.0 1e-06 
0.0 1.3136 0 2.0 1e-06 
0.0 1.3137 0 2.0 1e-06 
0.0 1.3138 0 2.0 1e-06 
0.0 1.3139 0 2.0 1e-06 
0.0 1.314 0 2.0 1e-06 
0.0 1.3141 0 2.0 1e-06 
0.0 1.3142 0 2.0 1e-06 
0.0 1.3143 0 2.0 1e-06 
0.0 1.3144 0 2.0 1e-06 
0.0 1.3145 0 2.0 1e-06 
0.0 1.3146 0 2.0 1e-06 
0.0 1.3147 0 2.0 1e-06 
0.0 1.3148 0 2.0 1e-06 
0.0 1.3149 0 2.0 1e-06 
0.0 1.315 0 2.0 1e-06 
0.0 1.3151 0 2.0 1e-06 
0.0 1.3152 0 2.0 1e-06 
0.0 1.3153 0 2.0 1e-06 
0.0 1.3154 0 2.0 1e-06 
0.0 1.3155 0 2.0 1e-06 
0.0 1.3156 0 2.0 1e-06 
0.0 1.3157 0 2.0 1e-06 
0.0 1.3158 0 2.0 1e-06 
0.0 1.3159 0 2.0 1e-06 
0.0 1.316 0 2.0 1e-06 
0.0 1.3161 0 2.0 1e-06 
0.0 1.3162 0 2.0 1e-06 
0.0 1.3163 0 2.0 1e-06 
0.0 1.3164 0 2.0 1e-06 
0.0 1.3165 0 2.0 1e-06 
0.0 1.3166 0 2.0 1e-06 
0.0 1.3167 0 2.0 1e-06 
0.0 1.3168 0 2.0 1e-06 
0.0 1.3169 0 2.0 1e-06 
0.0 1.317 0 2.0 1e-06 
0.0 1.3171 0 2.0 1e-06 
0.0 1.3172 0 2.0 1e-06 
0.0 1.3173 0 2.0 1e-06 
0.0 1.3174 0 2.0 1e-06 
0.0 1.3175 0 2.0 1e-06 
0.0 1.3176 0 2.0 1e-06 
0.0 1.3177 0 2.0 1e-06 
0.0 1.3178 0 2.0 1e-06 
0.0 1.3179 0 2.0 1e-06 
0.0 1.318 0 2.0 1e-06 
0.0 1.3181 0 2.0 1e-06 
0.0 1.3182 0 2.0 1e-06 
0.0 1.3183 0 2.0 1e-06 
0.0 1.3184 0 2.0 1e-06 
0.0 1.3185 0 2.0 1e-06 
0.0 1.3186 0 2.0 1e-06 
0.0 1.3187 0 2.0 1e-06 
0.0 1.3188 0 2.0 1e-06 
0.0 1.3189 0 2.0 1e-06 
0.0 1.319 0 2.0 1e-06 
0.0 1.3191 0 2.0 1e-06 
0.0 1.3192 0 2.0 1e-06 
0.0 1.3193 0 2.0 1e-06 
0.0 1.3194 0 2.0 1e-06 
0.0 1.3195 0 2.0 1e-06 
0.0 1.3196 0 2.0 1e-06 
0.0 1.3197 0 2.0 1e-06 
0.0 1.3198 0 2.0 1e-06 
0.0 1.3199 0 2.0 1e-06 
0.0 1.32 0 2.0 1e-06 
0.0 1.3201 0 2.0 1e-06 
0.0 1.3202 0 2.0 1e-06 
0.0 1.3203 0 2.0 1e-06 
0.0 1.3204 0 2.0 1e-06 
0.0 1.3205 0 2.0 1e-06 
0.0 1.3206 0 2.0 1e-06 
0.0 1.3207 0 2.0 1e-06 
0.0 1.3208 0 2.0 1e-06 
0.0 1.3209 0 2.0 1e-06 
0.0 1.321 0 2.0 1e-06 
0.0 1.3211 0 2.0 1e-06 
0.0 1.3212 0 2.0 1e-06 
0.0 1.3213 0 2.0 1e-06 
0.0 1.3214 0 2.0 1e-06 
0.0 1.3215 0 2.0 1e-06 
0.0 1.3216 0 2.0 1e-06 
0.0 1.3217 0 2.0 1e-06 
0.0 1.3218 0 2.0 1e-06 
0.0 1.3219 0 2.0 1e-06 
0.0 1.322 0 2.0 1e-06 
0.0 1.3221 0 2.0 1e-06 
0.0 1.3222 0 2.0 1e-06 
0.0 1.3223 0 2.0 1e-06 
0.0 1.3224 0 2.0 1e-06 
0.0 1.3225 0 2.0 1e-06 
0.0 1.3226 0 2.0 1e-06 
0.0 1.3227 0 2.0 1e-06 
0.0 1.3228 0 2.0 1e-06 
0.0 1.3229 0 2.0 1e-06 
0.0 1.323 0 2.0 1e-06 
0.0 1.3231 0 2.0 1e-06 
0.0 1.3232 0 2.0 1e-06 
0.0 1.3233 0 2.0 1e-06 
0.0 1.3234 0 2.0 1e-06 
0.0 1.3235 0 2.0 1e-06 
0.0 1.3236 0 2.0 1e-06 
0.0 1.3237 0 2.0 1e-06 
0.0 1.3238 0 2.0 1e-06 
0.0 1.3239 0 2.0 1e-06 
0.0 1.324 0 2.0 1e-06 
0.0 1.3241 0 2.0 1e-06 
0.0 1.3242 0 2.0 1e-06 
0.0 1.3243 0 2.0 1e-06 
0.0 1.3244 0 2.0 1e-06 
0.0 1.3245 0 2.0 1e-06 
0.0 1.3246 0 2.0 1e-06 
0.0 1.3247 0 2.0 1e-06 
0.0 1.3248 0 2.0 1e-06 
0.0 1.3249 0 2.0 1e-06 
0.0 1.325 0 2.0 1e-06 
0.0 1.3251 0 2.0 1e-06 
0.0 1.3252 0 2.0 1e-06 
0.0 1.3253 0 2.0 1e-06 
0.0 1.3254 0 2.0 1e-06 
0.0 1.3255 0 2.0 1e-06 
0.0 1.3256 0 2.0 1e-06 
0.0 1.3257 0 2.0 1e-06 
0.0 1.3258 0 2.0 1e-06 
0.0 1.3259 0 2.0 1e-06 
0.0 1.326 0 2.0 1e-06 
0.0 1.3261 0 2.0 1e-06 
0.0 1.3262 0 2.0 1e-06 
0.0 1.3263 0 2.0 1e-06 
0.0 1.3264 0 2.0 1e-06 
0.0 1.3265 0 2.0 1e-06 
0.0 1.3266 0 2.0 1e-06 
0.0 1.3267 0 2.0 1e-06 
0.0 1.3268 0 2.0 1e-06 
0.0 1.3269 0 2.0 1e-06 
0.0 1.327 0 2.0 1e-06 
0.0 1.3271 0 2.0 1e-06 
0.0 1.3272 0 2.0 1e-06 
0.0 1.3273 0 2.0 1e-06 
0.0 1.3274 0 2.0 1e-06 
0.0 1.3275 0 2.0 1e-06 
0.0 1.3276 0 2.0 1e-06 
0.0 1.3277 0 2.0 1e-06 
0.0 1.3278 0 2.0 1e-06 
0.0 1.3279 0 2.0 1e-06 
0.0 1.328 0 2.0 1e-06 
0.0 1.3281 0 2.0 1e-06 
0.0 1.3282 0 2.0 1e-06 
0.0 1.3283 0 2.0 1e-06 
0.0 1.3284 0 2.0 1e-06 
0.0 1.3285 0 2.0 1e-06 
0.0 1.3286 0 2.0 1e-06 
0.0 1.3287 0 2.0 1e-06 
0.0 1.3288 0 2.0 1e-06 
0.0 1.3289 0 2.0 1e-06 
0.0 1.329 0 2.0 1e-06 
0.0 1.3291 0 2.0 1e-06 
0.0 1.3292 0 2.0 1e-06 
0.0 1.3293 0 2.0 1e-06 
0.0 1.3294 0 2.0 1e-06 
0.0 1.3295 0 2.0 1e-06 
0.0 1.3296 0 2.0 1e-06 
0.0 1.3297 0 2.0 1e-06 
0.0 1.3298 0 2.0 1e-06 
0.0 1.3299 0 2.0 1e-06 
0.0 1.33 0 2.0 1e-06 
0.0 1.3301 0 2.0 1e-06 
0.0 1.3302 0 2.0 1e-06 
0.0 1.3303 0 2.0 1e-06 
0.0 1.3304 0 2.0 1e-06 
0.0 1.3305 0 2.0 1e-06 
0.0 1.3306 0 2.0 1e-06 
0.0 1.3307 0 2.0 1e-06 
0.0 1.3308 0 2.0 1e-06 
0.0 1.3309 0 2.0 1e-06 
0.0 1.331 0 2.0 1e-06 
0.0 1.3311 0 2.0 1e-06 
0.0 1.3312 0 2.0 1e-06 
0.0 1.3313 0 2.0 1e-06 
0.0 1.3314 0 2.0 1e-06 
0.0 1.3315 0 2.0 1e-06 
0.0 1.3316 0 2.0 1e-06 
0.0 1.3317 0 2.0 1e-06 
0.0 1.3318 0 2.0 1e-06 
0.0 1.3319 0 2.0 1e-06 
0.0 1.332 0 2.0 1e-06 
0.0 1.3321 0 2.0 1e-06 
0.0 1.3322 0 2.0 1e-06 
0.0 1.3323 0 2.0 1e-06 
0.0 1.3324 0 2.0 1e-06 
0.0 1.3325 0 2.0 1e-06 
0.0 1.3326 0 2.0 1e-06 
0.0 1.3327 0 2.0 1e-06 
0.0 1.3328 0 2.0 1e-06 
0.0 1.3329 0 2.0 1e-06 
0.0 1.333 0 2.0 1e-06 
0.0 1.3331 0 2.0 1e-06 
0.0 1.3332 0 2.0 1e-06 
0.0 1.3333 0 2.0 1e-06 
0.0 1.3334 0 2.0 1e-06 
0.0 1.3335 0 2.0 1e-06 
0.0 1.3336 0 2.0 1e-06 
0.0 1.3337 0 2.0 1e-06 
0.0 1.3338 0 2.0 1e-06 
0.0 1.3339 0 2.0 1e-06 
0.0 1.334 0 2.0 1e-06 
0.0 1.3341 0 2.0 1e-06 
0.0 1.3342 0 2.0 1e-06 
0.0 1.3343 0 2.0 1e-06 
0.0 1.3344 0 2.0 1e-06 
0.0 1.3345 0 2.0 1e-06 
0.0 1.3346 0 2.0 1e-06 
0.0 1.3347 0 2.0 1e-06 
0.0 1.3348 0 2.0 1e-06 
0.0 1.3349 0 2.0 1e-06 
0.0 1.335 0 2.0 1e-06 
0.0 1.3351 0 2.0 1e-06 
0.0 1.3352 0 2.0 1e-06 
0.0 1.3353 0 2.0 1e-06 
0.0 1.3354 0 2.0 1e-06 
0.0 1.3355 0 2.0 1e-06 
0.0 1.3356 0 2.0 1e-06 
0.0 1.3357 0 2.0 1e-06 
0.0 1.3358 0 2.0 1e-06 
0.0 1.3359 0 2.0 1e-06 
0.0 1.336 0 2.0 1e-06 
0.0 1.3361 0 2.0 1e-06 
0.0 1.3362 0 2.0 1e-06 
0.0 1.3363 0 2.0 1e-06 
0.0 1.3364 0 2.0 1e-06 
0.0 1.3365 0 2.0 1e-06 
0.0 1.3366 0 2.0 1e-06 
0.0 1.3367 0 2.0 1e-06 
0.0 1.3368 0 2.0 1e-06 
0.0 1.3369 0 2.0 1e-06 
0.0 1.337 0 2.0 1e-06 
0.0 1.3371 0 2.0 1e-06 
0.0 1.3372 0 2.0 1e-06 
0.0 1.3373 0 2.0 1e-06 
0.0 1.3374 0 2.0 1e-06 
0.0 1.3375 0 2.0 1e-06 
0.0 1.3376 0 2.0 1e-06 
0.0 1.3377 0 2.0 1e-06 
0.0 1.3378 0 2.0 1e-06 
0.0 1.3379 0 2.0 1e-06 
0.0 1.338 0 2.0 1e-06 
0.0 1.3381 0 2.0 1e-06 
0.0 1.3382 0 2.0 1e-06 
0.0 1.3383 0 2.0 1e-06 
0.0 1.3384 0 2.0 1e-06 
0.0 1.3385 0 2.0 1e-06 
0.0 1.3386 0 2.0 1e-06 
0.0 1.3387 0 2.0 1e-06 
0.0 1.3388 0 2.0 1e-06 
0.0 1.3389 0 2.0 1e-06 
0.0 1.339 0 2.0 1e-06 
0.0 1.3391 0 2.0 1e-06 
0.0 1.3392 0 2.0 1e-06 
0.0 1.3393 0 2.0 1e-06 
0.0 1.3394 0 2.0 1e-06 
0.0 1.3395 0 2.0 1e-06 
0.0 1.3396 0 2.0 1e-06 
0.0 1.3397 0 2.0 1e-06 
0.0 1.3398 0 2.0 1e-06 
0.0 1.3399 0 2.0 1e-06 
0.0 1.34 0 2.0 1e-06 
0.0 1.3401 0 2.0 1e-06 
0.0 1.3402 0 2.0 1e-06 
0.0 1.3403 0 2.0 1e-06 
0.0 1.3404 0 2.0 1e-06 
0.0 1.3405 0 2.0 1e-06 
0.0 1.3406 0 2.0 1e-06 
0.0 1.3407 0 2.0 1e-06 
0.0 1.3408 0 2.0 1e-06 
0.0 1.3409 0 2.0 1e-06 
0.0 1.341 0 2.0 1e-06 
0.0 1.3411 0 2.0 1e-06 
0.0 1.3412 0 2.0 1e-06 
0.0 1.3413 0 2.0 1e-06 
0.0 1.3414 0 2.0 1e-06 
0.0 1.3415 0 2.0 1e-06 
0.0 1.3416 0 2.0 1e-06 
0.0 1.3417 0 2.0 1e-06 
0.0 1.3418 0 2.0 1e-06 
0.0 1.3419 0 2.0 1e-06 
0.0 1.342 0 2.0 1e-06 
0.0 1.3421 0 2.0 1e-06 
0.0 1.3422 0 2.0 1e-06 
0.0 1.3423 0 2.0 1e-06 
0.0 1.3424 0 2.0 1e-06 
0.0 1.3425 0 2.0 1e-06 
0.0 1.3426 0 2.0 1e-06 
0.0 1.3427 0 2.0 1e-06 
0.0 1.3428 0 2.0 1e-06 
0.0 1.3429 0 2.0 1e-06 
0.0 1.343 0 2.0 1e-06 
0.0 1.3431 0 2.0 1e-06 
0.0 1.3432 0 2.0 1e-06 
0.0 1.3433 0 2.0 1e-06 
0.0 1.3434 0 2.0 1e-06 
0.0 1.3435 0 2.0 1e-06 
0.0 1.3436 0 2.0 1e-06 
0.0 1.3437 0 2.0 1e-06 
0.0 1.3438 0 2.0 1e-06 
0.0 1.3439 0 2.0 1e-06 
0.0 1.344 0 2.0 1e-06 
0.0 1.3441 0 2.0 1e-06 
0.0 1.3442 0 2.0 1e-06 
0.0 1.3443 0 2.0 1e-06 
0.0 1.3444 0 2.0 1e-06 
0.0 1.3445 0 2.0 1e-06 
0.0 1.3446 0 2.0 1e-06 
0.0 1.3447 0 2.0 1e-06 
0.0 1.3448 0 2.0 1e-06 
0.0 1.3449 0 2.0 1e-06 
0.0 1.345 0 2.0 1e-06 
0.0 1.3451 0 2.0 1e-06 
0.0 1.3452 0 2.0 1e-06 
0.0 1.3453 0 2.0 1e-06 
0.0 1.3454 0 2.0 1e-06 
0.0 1.3455 0 2.0 1e-06 
0.0 1.3456 0 2.0 1e-06 
0.0 1.3457 0 2.0 1e-06 
0.0 1.3458 0 2.0 1e-06 
0.0 1.3459 0 2.0 1e-06 
0.0 1.346 0 2.0 1e-06 
0.0 1.3461 0 2.0 1e-06 
0.0 1.3462 0 2.0 1e-06 
0.0 1.3463 0 2.0 1e-06 
0.0 1.3464 0 2.0 1e-06 
0.0 1.3465 0 2.0 1e-06 
0.0 1.3466 0 2.0 1e-06 
0.0 1.3467 0 2.0 1e-06 
0.0 1.3468 0 2.0 1e-06 
0.0 1.3469 0 2.0 1e-06 
0.0 1.347 0 2.0 1e-06 
0.0 1.3471 0 2.0 1e-06 
0.0 1.3472 0 2.0 1e-06 
0.0 1.3473 0 2.0 1e-06 
0.0 1.3474 0 2.0 1e-06 
0.0 1.3475 0 2.0 1e-06 
0.0 1.3476 0 2.0 1e-06 
0.0 1.3477 0 2.0 1e-06 
0.0 1.3478 0 2.0 1e-06 
0.0 1.3479 0 2.0 1e-06 
0.0 1.348 0 2.0 1e-06 
0.0 1.3481 0 2.0 1e-06 
0.0 1.3482 0 2.0 1e-06 
0.0 1.3483 0 2.0 1e-06 
0.0 1.3484 0 2.0 1e-06 
0.0 1.3485 0 2.0 1e-06 
0.0 1.3486 0 2.0 1e-06 
0.0 1.3487 0 2.0 1e-06 
0.0 1.3488 0 2.0 1e-06 
0.0 1.3489 0 2.0 1e-06 
0.0 1.349 0 2.0 1e-06 
0.0 1.3491 0 2.0 1e-06 
0.0 1.3492 0 2.0 1e-06 
0.0 1.3493 0 2.0 1e-06 
0.0 1.3494 0 2.0 1e-06 
0.0 1.3495 0 2.0 1e-06 
0.0 1.3496 0 2.0 1e-06 
0.0 1.3497 0 2.0 1e-06 
0.0 1.3498 0 2.0 1e-06 
0.0 1.3499 0 2.0 1e-06 
0.0 1.35 0 2.0 1e-06 
0.0 1.3501 0 2.0 1e-06 
0.0 1.3502 0 2.0 1e-06 
0.0 1.3503 0 2.0 1e-06 
0.0 1.3504 0 2.0 1e-06 
0.0 1.3505 0 2.0 1e-06 
0.0 1.3506 0 2.0 1e-06 
0.0 1.3507 0 2.0 1e-06 
0.0 1.3508 0 2.0 1e-06 
0.0 1.3509 0 2.0 1e-06 
0.0 1.351 0 2.0 1e-06 
0.0 1.3511 0 2.0 1e-06 
0.0 1.3512 0 2.0 1e-06 
0.0 1.3513 0 2.0 1e-06 
0.0 1.3514 0 2.0 1e-06 
0.0 1.3515 0 2.0 1e-06 
0.0 1.3516 0 2.0 1e-06 
0.0 1.3517 0 2.0 1e-06 
0.0 1.3518 0 2.0 1e-06 
0.0 1.3519 0 2.0 1e-06 
0.0 1.352 0 2.0 1e-06 
0.0 1.3521 0 2.0 1e-06 
0.0 1.3522 0 2.0 1e-06 
0.0 1.3523 0 2.0 1e-06 
0.0 1.3524 0 2.0 1e-06 
0.0 1.3525 0 2.0 1e-06 
0.0 1.3526 0 2.0 1e-06 
0.0 1.3527 0 2.0 1e-06 
0.0 1.3528 0 2.0 1e-06 
0.0 1.3529 0 2.0 1e-06 
0.0 1.353 0 2.0 1e-06 
0.0 1.3531 0 2.0 1e-06 
0.0 1.3532 0 2.0 1e-06 
0.0 1.3533 0 2.0 1e-06 
0.0 1.3534 0 2.0 1e-06 
0.0 1.3535 0 2.0 1e-06 
0.0 1.3536 0 2.0 1e-06 
0.0 1.3537 0 2.0 1e-06 
0.0 1.3538 0 2.0 1e-06 
0.0 1.3539 0 2.0 1e-06 
0.0 1.354 0 2.0 1e-06 
0.0 1.3541 0 2.0 1e-06 
0.0 1.3542 0 2.0 1e-06 
0.0 1.3543 0 2.0 1e-06 
0.0 1.3544 0 2.0 1e-06 
0.0 1.3545 0 2.0 1e-06 
0.0 1.3546 0 2.0 1e-06 
0.0 1.3547 0 2.0 1e-06 
0.0 1.3548 0 2.0 1e-06 
0.0 1.3549 0 2.0 1e-06 
0.0 1.355 0 2.0 1e-06 
0.0 1.3551 0 2.0 1e-06 
0.0 1.3552 0 2.0 1e-06 
0.0 1.3553 0 2.0 1e-06 
0.0 1.3554 0 2.0 1e-06 
0.0 1.3555 0 2.0 1e-06 
0.0 1.3556 0 2.0 1e-06 
0.0 1.3557 0 2.0 1e-06 
0.0 1.3558 0 2.0 1e-06 
0.0 1.3559 0 2.0 1e-06 
0.0 1.356 0 2.0 1e-06 
0.0 1.3561 0 2.0 1e-06 
0.0 1.3562 0 2.0 1e-06 
0.0 1.3563 0 2.0 1e-06 
0.0 1.3564 0 2.0 1e-06 
0.0 1.3565 0 2.0 1e-06 
0.0 1.3566 0 2.0 1e-06 
0.0 1.3567 0 2.0 1e-06 
0.0 1.3568 0 2.0 1e-06 
0.0 1.3569 0 2.0 1e-06 
0.0 1.357 0 2.0 1e-06 
0.0 1.3571 0 2.0 1e-06 
0.0 1.3572 0 2.0 1e-06 
0.0 1.3573 0 2.0 1e-06 
0.0 1.3574 0 2.0 1e-06 
0.0 1.3575 0 2.0 1e-06 
0.0 1.3576 0 2.0 1e-06 
0.0 1.3577 0 2.0 1e-06 
0.0 1.3578 0 2.0 1e-06 
0.0 1.3579 0 2.0 1e-06 
0.0 1.358 0 2.0 1e-06 
0.0 1.3581 0 2.0 1e-06 
0.0 1.3582 0 2.0 1e-06 
0.0 1.3583 0 2.0 1e-06 
0.0 1.3584 0 2.0 1e-06 
0.0 1.3585 0 2.0 1e-06 
0.0 1.3586 0 2.0 1e-06 
0.0 1.3587 0 2.0 1e-06 
0.0 1.3588 0 2.0 1e-06 
0.0 1.3589 0 2.0 1e-06 
0.0 1.359 0 2.0 1e-06 
0.0 1.3591 0 2.0 1e-06 
0.0 1.3592 0 2.0 1e-06 
0.0 1.3593 0 2.0 1e-06 
0.0 1.3594 0 2.0 1e-06 
0.0 1.3595 0 2.0 1e-06 
0.0 1.3596 0 2.0 1e-06 
0.0 1.3597 0 2.0 1e-06 
0.0 1.3598 0 2.0 1e-06 
0.0 1.3599 0 2.0 1e-06 
0.0 1.36 0 2.0 1e-06 
0.0 1.3601 0 2.0 1e-06 
0.0 1.3602 0 2.0 1e-06 
0.0 1.3603 0 2.0 1e-06 
0.0 1.3604 0 2.0 1e-06 
0.0 1.3605 0 2.0 1e-06 
0.0 1.3606 0 2.0 1e-06 
0.0 1.3607 0 2.0 1e-06 
0.0 1.3608 0 2.0 1e-06 
0.0 1.3609 0 2.0 1e-06 
0.0 1.361 0 2.0 1e-06 
0.0 1.3611 0 2.0 1e-06 
0.0 1.3612 0 2.0 1e-06 
0.0 1.3613 0 2.0 1e-06 
0.0 1.3614 0 2.0 1e-06 
0.0 1.3615 0 2.0 1e-06 
0.0 1.3616 0 2.0 1e-06 
0.0 1.3617 0 2.0 1e-06 
0.0 1.3618 0 2.0 1e-06 
0.0 1.3619 0 2.0 1e-06 
0.0 1.362 0 2.0 1e-06 
0.0 1.3621 0 2.0 1e-06 
0.0 1.3622 0 2.0 1e-06 
0.0 1.3623 0 2.0 1e-06 
0.0 1.3624 0 2.0 1e-06 
0.0 1.3625 0 2.0 1e-06 
0.0 1.3626 0 2.0 1e-06 
0.0 1.3627 0 2.0 1e-06 
0.0 1.3628 0 2.0 1e-06 
0.0 1.3629 0 2.0 1e-06 
0.0 1.363 0 2.0 1e-06 
0.0 1.3631 0 2.0 1e-06 
0.0 1.3632 0 2.0 1e-06 
0.0 1.3633 0 2.0 1e-06 
0.0 1.3634 0 2.0 1e-06 
0.0 1.3635 0 2.0 1e-06 
0.0 1.3636 0 2.0 1e-06 
0.0 1.3637 0 2.0 1e-06 
0.0 1.3638 0 2.0 1e-06 
0.0 1.3639 0 2.0 1e-06 
0.0 1.364 0 2.0 1e-06 
0.0 1.3641 0 2.0 1e-06 
0.0 1.3642 0 2.0 1e-06 
0.0 1.3643 0 2.0 1e-06 
0.0 1.3644 0 2.0 1e-06 
0.0 1.3645 0 2.0 1e-06 
0.0 1.3646 0 2.0 1e-06 
0.0 1.3647 0 2.0 1e-06 
0.0 1.3648 0 2.0 1e-06 
0.0 1.3649 0 2.0 1e-06 
0.0 1.365 0 2.0 1e-06 
0.0 1.3651 0 2.0 1e-06 
0.0 1.3652 0 2.0 1e-06 
0.0 1.3653 0 2.0 1e-06 
0.0 1.3654 0 2.0 1e-06 
0.0 1.3655 0 2.0 1e-06 
0.0 1.3656 0 2.0 1e-06 
0.0 1.3657 0 2.0 1e-06 
0.0 1.3658 0 2.0 1e-06 
0.0 1.3659 0 2.0 1e-06 
0.0 1.366 0 2.0 1e-06 
0.0 1.3661 0 2.0 1e-06 
0.0 1.3662 0 2.0 1e-06 
0.0 1.3663 0 2.0 1e-06 
0.0 1.3664 0 2.0 1e-06 
0.0 1.3665 0 2.0 1e-06 
0.0 1.3666 0 2.0 1e-06 
0.0 1.3667 0 2.0 1e-06 
0.0 1.3668 0 2.0 1e-06 
0.0 1.3669 0 2.0 1e-06 
0.0 1.367 0 2.0 1e-06 
0.0 1.3671 0 2.0 1e-06 
0.0 1.3672 0 2.0 1e-06 
0.0 1.3673 0 2.0 1e-06 
0.0 1.3674 0 2.0 1e-06 
0.0 1.3675 0 2.0 1e-06 
0.0 1.3676 0 2.0 1e-06 
0.0 1.3677 0 2.0 1e-06 
0.0 1.3678 0 2.0 1e-06 
0.0 1.3679 0 2.0 1e-06 
0.0 1.368 0 2.0 1e-06 
0.0 1.3681 0 2.0 1e-06 
0.0 1.3682 0 2.0 1e-06 
0.0 1.3683 0 2.0 1e-06 
0.0 1.3684 0 2.0 1e-06 
0.0 1.3685 0 2.0 1e-06 
0.0 1.3686 0 2.0 1e-06 
0.0 1.3687 0 2.0 1e-06 
0.0 1.3688 0 2.0 1e-06 
0.0 1.3689 0 2.0 1e-06 
0.0 1.369 0 2.0 1e-06 
0.0 1.3691 0 2.0 1e-06 
0.0 1.3692 0 2.0 1e-06 
0.0 1.3693 0 2.0 1e-06 
0.0 1.3694 0 2.0 1e-06 
0.0 1.3695 0 2.0 1e-06 
0.0 1.3696 0 2.0 1e-06 
0.0 1.3697 0 2.0 1e-06 
0.0 1.3698 0 2.0 1e-06 
0.0 1.3699 0 2.0 1e-06 
0.0 1.37 0 2.0 1e-06 
0.0 1.3701 0 2.0 1e-06 
0.0 1.3702 0 2.0 1e-06 
0.0 1.3703 0 2.0 1e-06 
0.0 1.3704 0 2.0 1e-06 
0.0 1.3705 0 2.0 1e-06 
0.0 1.3706 0 2.0 1e-06 
0.0 1.3707 0 2.0 1e-06 
0.0 1.3708 0 2.0 1e-06 
0.0 1.3709 0 2.0 1e-06 
0.0 1.371 0 2.0 1e-06 
0.0 1.3711 0 2.0 1e-06 
0.0 1.3712 0 2.0 1e-06 
0.0 1.3713 0 2.0 1e-06 
0.0 1.3714 0 2.0 1e-06 
0.0 1.3715 0 2.0 1e-06 
0.0 1.3716 0 2.0 1e-06 
0.0 1.3717 0 2.0 1e-06 
0.0 1.3718 0 2.0 1e-06 
0.0 1.3719 0 2.0 1e-06 
0.0 1.372 0 2.0 1e-06 
0.0 1.3721 0 2.0 1e-06 
0.0 1.3722 0 2.0 1e-06 
0.0 1.3723 0 2.0 1e-06 
0.0 1.3724 0 2.0 1e-06 
0.0 1.3725 0 2.0 1e-06 
0.0 1.3726 0 2.0 1e-06 
0.0 1.3727 0 2.0 1e-06 
0.0 1.3728 0 2.0 1e-06 
0.0 1.3729 0 2.0 1e-06 
0.0 1.373 0 2.0 1e-06 
0.0 1.3731 0 2.0 1e-06 
0.0 1.3732 0 2.0 1e-06 
0.0 1.3733 0 2.0 1e-06 
0.0 1.3734 0 2.0 1e-06 
0.0 1.3735 0 2.0 1e-06 
0.0 1.3736 0 2.0 1e-06 
0.0 1.3737 0 2.0 1e-06 
0.0 1.3738 0 2.0 1e-06 
0.0 1.3739 0 2.0 1e-06 
0.0 1.374 0 2.0 1e-06 
0.0 1.3741 0 2.0 1e-06 
0.0 1.3742 0 2.0 1e-06 
0.0 1.3743 0 2.0 1e-06 
0.0 1.3744 0 2.0 1e-06 
0.0 1.3745 0 2.0 1e-06 
0.0 1.3746 0 2.0 1e-06 
0.0 1.3747 0 2.0 1e-06 
0.0 1.3748 0 2.0 1e-06 
0.0 1.3749 0 2.0 1e-06 
0.0 1.375 0 2.0 1e-06 
0.0 1.3751 0 2.0 1e-06 
0.0 1.3752 0 2.0 1e-06 
0.0 1.3753 0 2.0 1e-06 
0.0 1.3754 0 2.0 1e-06 
0.0 1.3755 0 2.0 1e-06 
0.0 1.3756 0 2.0 1e-06 
0.0 1.3757 0 2.0 1e-06 
0.0 1.3758 0 2.0 1e-06 
0.0 1.3759 0 2.0 1e-06 
0.0 1.376 0 2.0 1e-06 
0.0 1.3761 0 2.0 1e-06 
0.0 1.3762 0 2.0 1e-06 
0.0 1.3763 0 2.0 1e-06 
0.0 1.3764 0 2.0 1e-06 
0.0 1.3765 0 2.0 1e-06 
0.0 1.3766 0 2.0 1e-06 
0.0 1.3767 0 2.0 1e-06 
0.0 1.3768 0 2.0 1e-06 
0.0 1.3769 0 2.0 1e-06 
0.0 1.377 0 2.0 1e-06 
0.0 1.3771 0 2.0 1e-06 
0.0 1.3772 0 2.0 1e-06 
0.0 1.3773 0 2.0 1e-06 
0.0 1.3774 0 2.0 1e-06 
0.0 1.3775 0 2.0 1e-06 
0.0 1.3776 0 2.0 1e-06 
0.0 1.3777 0 2.0 1e-06 
0.0 1.3778 0 2.0 1e-06 
0.0 1.3779 0 2.0 1e-06 
0.0 1.378 0 2.0 1e-06 
0.0 1.3781 0 2.0 1e-06 
0.0 1.3782 0 2.0 1e-06 
0.0 1.3783 0 2.0 1e-06 
0.0 1.3784 0 2.0 1e-06 
0.0 1.3785 0 2.0 1e-06 
0.0 1.3786 0 2.0 1e-06 
0.0 1.3787 0 2.0 1e-06 
0.0 1.3788 0 2.0 1e-06 
0.0 1.3789 0 2.0 1e-06 
0.0 1.379 0 2.0 1e-06 
0.0 1.3791 0 2.0 1e-06 
0.0 1.3792 0 2.0 1e-06 
0.0 1.3793 0 2.0 1e-06 
0.0 1.3794 0 2.0 1e-06 
0.0 1.3795 0 2.0 1e-06 
0.0 1.3796 0 2.0 1e-06 
0.0 1.3797 0 2.0 1e-06 
0.0 1.3798 0 2.0 1e-06 
0.0 1.3799 0 2.0 1e-06 
0.0 1.38 0 2.0 1e-06 
0.0 1.3801 0 2.0 1e-06 
0.0 1.3802 0 2.0 1e-06 
0.0 1.3803 0 2.0 1e-06 
0.0 1.3804 0 2.0 1e-06 
0.0 1.3805 0 2.0 1e-06 
0.0 1.3806 0 2.0 1e-06 
0.0 1.3807 0 2.0 1e-06 
0.0 1.3808 0 2.0 1e-06 
0.0 1.3809 0 2.0 1e-06 
0.0 1.381 0 2.0 1e-06 
0.0 1.3811 0 2.0 1e-06 
0.0 1.3812 0 2.0 1e-06 
0.0 1.3813 0 2.0 1e-06 
0.0 1.3814 0 2.0 1e-06 
0.0 1.3815 0 2.0 1e-06 
0.0 1.3816 0 2.0 1e-06 
0.0 1.3817 0 2.0 1e-06 
0.0 1.3818 0 2.0 1e-06 
0.0 1.3819 0 2.0 1e-06 
0.0 1.382 0 2.0 1e-06 
0.0 1.3821 0 2.0 1e-06 
0.0 1.3822 0 2.0 1e-06 
0.0 1.3823 0 2.0 1e-06 
0.0 1.3824 0 2.0 1e-06 
0.0 1.3825 0 2.0 1e-06 
0.0 1.3826 0 2.0 1e-06 
0.0 1.3827 0 2.0 1e-06 
0.0 1.3828 0 2.0 1e-06 
0.0 1.3829 0 2.0 1e-06 
0.0 1.383 0 2.0 1e-06 
0.0 1.3831 0 2.0 1e-06 
0.0 1.3832 0 2.0 1e-06 
0.0 1.3833 0 2.0 1e-06 
0.0 1.3834 0 2.0 1e-06 
0.0 1.3835 0 2.0 1e-06 
0.0 1.3836 0 2.0 1e-06 
0.0 1.3837 0 2.0 1e-06 
0.0 1.3838 0 2.0 1e-06 
0.0 1.3839 0 2.0 1e-06 
0.0 1.384 0 2.0 1e-06 
0.0 1.3841 0 2.0 1e-06 
0.0 1.3842 0 2.0 1e-06 
0.0 1.3843 0 2.0 1e-06 
0.0 1.3844 0 2.0 1e-06 
0.0 1.3845 0 2.0 1e-06 
0.0 1.3846 0 2.0 1e-06 
0.0 1.3847 0 2.0 1e-06 
0.0 1.3848 0 2.0 1e-06 
0.0 1.3849 0 2.0 1e-06 
0.0 1.385 0 2.0 1e-06 
0.0 1.3851 0 2.0 1e-06 
0.0 1.3852 0 2.0 1e-06 
0.0 1.3853 0 2.0 1e-06 
0.0 1.3854 0 2.0 1e-06 
0.0 1.3855 0 2.0 1e-06 
0.0 1.3856 0 2.0 1e-06 
0.0 1.3857 0 2.0 1e-06 
0.0 1.3858 0 2.0 1e-06 
0.0 1.3859 0 2.0 1e-06 
0.0 1.386 0 2.0 1e-06 
0.0 1.3861 0 2.0 1e-06 
0.0 1.3862 0 2.0 1e-06 
0.0 1.3863 0 2.0 1e-06 
0.0 1.3864 0 2.0 1e-06 
0.0 1.3865 0 2.0 1e-06 
0.0 1.3866 0 2.0 1e-06 
0.0 1.3867 0 2.0 1e-06 
0.0 1.3868 0 2.0 1e-06 
0.0 1.3869 0 2.0 1e-06 
0.0 1.387 0 2.0 1e-06 
0.0 1.3871 0 2.0 1e-06 
0.0 1.3872 0 2.0 1e-06 
0.0 1.3873 0 2.0 1e-06 
0.0 1.3874 0 2.0 1e-06 
0.0 1.3875 0 2.0 1e-06 
0.0 1.3876 0 2.0 1e-06 
0.0 1.3877 0 2.0 1e-06 
0.0 1.3878 0 2.0 1e-06 
0.0 1.3879 0 2.0 1e-06 
0.0 1.388 0 2.0 1e-06 
0.0 1.3881 0 2.0 1e-06 
0.0 1.3882 0 2.0 1e-06 
0.0 1.3883 0 2.0 1e-06 
0.0 1.3884 0 2.0 1e-06 
0.0 1.3885 0 2.0 1e-06 
0.0 1.3886 0 2.0 1e-06 
0.0 1.3887 0 2.0 1e-06 
0.0 1.3888 0 2.0 1e-06 
0.0 1.3889 0 2.0 1e-06 
0.0 1.389 0 2.0 1e-06 
0.0 1.3891 0 2.0 1e-06 
0.0 1.3892 0 2.0 1e-06 
0.0 1.3893 0 2.0 1e-06 
0.0 1.3894 0 2.0 1e-06 
0.0 1.3895 0 2.0 1e-06 
0.0 1.3896 0 2.0 1e-06 
0.0 1.3897 0 2.0 1e-06 
0.0 1.3898 0 2.0 1e-06 
0.0 1.3899 0 2.0 1e-06 
0.0 1.39 0 2.0 1e-06 
0.0 1.3901 0 2.0 1e-06 
0.0 1.3902 0 2.0 1e-06 
0.0 1.3903 0 2.0 1e-06 
0.0 1.3904 0 2.0 1e-06 
0.0 1.3905 0 2.0 1e-06 
0.0 1.3906 0 2.0 1e-06 
0.0 1.3907 0 2.0 1e-06 
0.0 1.3908 0 2.0 1e-06 
0.0 1.3909 0 2.0 1e-06 
0.0 1.391 0 2.0 1e-06 
0.0 1.3911 0 2.0 1e-06 
0.0 1.3912 0 2.0 1e-06 
0.0 1.3913 0 2.0 1e-06 
0.0 1.3914 0 2.0 1e-06 
0.0 1.3915 0 2.0 1e-06 
0.0 1.3916 0 2.0 1e-06 
0.0 1.3917 0 2.0 1e-06 
0.0 1.3918 0 2.0 1e-06 
0.0 1.3919 0 2.0 1e-06 
0.0 1.392 0 2.0 1e-06 
0.0 1.3921 0 2.0 1e-06 
0.0 1.3922 0 2.0 1e-06 
0.0 1.3923 0 2.0 1e-06 
0.0 1.3924 0 2.0 1e-06 
0.0 1.3925 0 2.0 1e-06 
0.0 1.3926 0 2.0 1e-06 
0.0 1.3927 0 2.0 1e-06 
0.0 1.3928 0 2.0 1e-06 
0.0 1.3929 0 2.0 1e-06 
0.0 1.393 0 2.0 1e-06 
0.0 1.3931 0 2.0 1e-06 
0.0 1.3932 0 2.0 1e-06 
0.0 1.3933 0 2.0 1e-06 
0.0 1.3934 0 2.0 1e-06 
0.0 1.3935 0 2.0 1e-06 
0.0 1.3936 0 2.0 1e-06 
0.0 1.3937 0 2.0 1e-06 
0.0 1.3938 0 2.0 1e-06 
0.0 1.3939 0 2.0 1e-06 
0.0 1.394 0 2.0 1e-06 
0.0 1.3941 0 2.0 1e-06 
0.0 1.3942 0 2.0 1e-06 
0.0 1.3943 0 2.0 1e-06 
0.0 1.3944 0 2.0 1e-06 
0.0 1.3945 0 2.0 1e-06 
0.0 1.3946 0 2.0 1e-06 
0.0 1.3947 0 2.0 1e-06 
0.0 1.3948 0 2.0 1e-06 
0.0 1.3949 0 2.0 1e-06 
0.0 1.395 0 2.0 1e-06 
0.0 1.3951 0 2.0 1e-06 
0.0 1.3952 0 2.0 1e-06 
0.0 1.3953 0 2.0 1e-06 
0.0 1.3954 0 2.0 1e-06 
0.0 1.3955 0 2.0 1e-06 
0.0 1.3956 0 2.0 1e-06 
0.0 1.3957 0 2.0 1e-06 
0.0 1.3958 0 2.0 1e-06 
0.0 1.3959 0 2.0 1e-06 
0.0 1.396 0 2.0 1e-06 
0.0 1.3961 0 2.0 1e-06 
0.0 1.3962 0 2.0 1e-06 
0.0 1.3963 0 2.0 1e-06 
0.0 1.3964 0 2.0 1e-06 
0.0 1.3965 0 2.0 1e-06 
0.0 1.3966 0 2.0 1e-06 
0.0 1.3967 0 2.0 1e-06 
0.0 1.3968 0 2.0 1e-06 
0.0 1.3969 0 2.0 1e-06 
0.0 1.397 0 2.0 1e-06 
0.0 1.3971 0 2.0 1e-06 
0.0 1.3972 0 2.0 1e-06 
0.0 1.3973 0 2.0 1e-06 
0.0 1.3974 0 2.0 1e-06 
0.0 1.3975 0 2.0 1e-06 
0.0 1.3976 0 2.0 1e-06 
0.0 1.3977 0 2.0 1e-06 
0.0 1.3978 0 2.0 1e-06 
0.0 1.3979 0 2.0 1e-06 
0.0 1.398 0 2.0 1e-06 
0.0 1.3981 0 2.0 1e-06 
0.0 1.3982 0 2.0 1e-06 
0.0 1.3983 0 2.0 1e-06 
0.0 1.3984 0 2.0 1e-06 
0.0 1.3985 0 2.0 1e-06 
0.0 1.3986 0 2.0 1e-06 
0.0 1.3987 0 2.0 1e-06 
0.0 1.3988 0 2.0 1e-06 
0.0 1.3989 0 2.0 1e-06 
0.0 1.399 0 2.0 1e-06 
0.0 1.3991 0 2.0 1e-06 
0.0 1.3992 0 2.0 1e-06 
0.0 1.3993 0 2.0 1e-06 
0.0 1.3994 0 2.0 1e-06 
0.0 1.3995 0 2.0 1e-06 
0.0 1.3996 0 2.0 1e-06 
0.0 1.3997 0 2.0 1e-06 
0.0 1.3998 0 2.0 1e-06 
0.0 1.3999 0 2.0 1e-06 
0.0 1.4 0 2.0 1e-06 
0.0 1.4001 0 2.0 1e-06 
0.0 1.4002 0 2.0 1e-06 
0.0 1.4003 0 2.0 1e-06 
0.0 1.4004 0 2.0 1e-06 
0.0 1.4005 0 2.0 1e-06 
0.0 1.4006 0 2.0 1e-06 
0.0 1.4007 0 2.0 1e-06 
0.0 1.4008 0 2.0 1e-06 
0.0 1.4009 0 2.0 1e-06 
0.0 1.401 0 2.0 1e-06 
0.0 1.4011 0 2.0 1e-06 
0.0 1.4012 0 2.0 1e-06 
0.0 1.4013 0 2.0 1e-06 
0.0 1.4014 0 2.0 1e-06 
0.0 1.4015 0 2.0 1e-06 
0.0 1.4016 0 2.0 1e-06 
0.0 1.4017 0 2.0 1e-06 
0.0 1.4018 0 2.0 1e-06 
0.0 1.4019 0 2.0 1e-06 
0.0 1.402 0 2.0 1e-06 
0.0 1.4021 0 2.0 1e-06 
0.0 1.4022 0 2.0 1e-06 
0.0 1.4023 0 2.0 1e-06 
0.0 1.4024 0 2.0 1e-06 
0.0 1.4025 0 2.0 1e-06 
0.0 1.4026 0 2.0 1e-06 
0.0 1.4027 0 2.0 1e-06 
0.0 1.4028 0 2.0 1e-06 
0.0 1.4029 0 2.0 1e-06 
0.0 1.403 0 2.0 1e-06 
0.0 1.4031 0 2.0 1e-06 
0.0 1.4032 0 2.0 1e-06 
0.0 1.4033 0 2.0 1e-06 
0.0 1.4034 0 2.0 1e-06 
0.0 1.4035 0 2.0 1e-06 
0.0 1.4036 0 2.0 1e-06 
0.0 1.4037 0 2.0 1e-06 
0.0 1.4038 0 2.0 1e-06 
0.0 1.4039 0 2.0 1e-06 
0.0 1.404 0 2.0 1e-06 
0.0 1.4041 0 2.0 1e-06 
0.0 1.4042 0 2.0 1e-06 
0.0 1.4043 0 2.0 1e-06 
0.0 1.4044 0 2.0 1e-06 
0.0 1.4045 0 2.0 1e-06 
0.0 1.4046 0 2.0 1e-06 
0.0 1.4047 0 2.0 1e-06 
0.0 1.4048 0 2.0 1e-06 
0.0 1.4049 0 2.0 1e-06 
0.0 1.405 0 2.0 1e-06 
0.0 1.4051 0 2.0 1e-06 
0.0 1.4052 0 2.0 1e-06 
0.0 1.4053 0 2.0 1e-06 
0.0 1.4054 0 2.0 1e-06 
0.0 1.4055 0 2.0 1e-06 
0.0 1.4056 0 2.0 1e-06 
0.0 1.4057 0 2.0 1e-06 
0.0 1.4058 0 2.0 1e-06 
0.0 1.4059 0 2.0 1e-06 
0.0 1.406 0 2.0 1e-06 
0.0 1.4061 0 2.0 1e-06 
0.0 1.4062 0 2.0 1e-06 
0.0 1.4063 0 2.0 1e-06 
0.0 1.4064 0 2.0 1e-06 
0.0 1.4065 0 2.0 1e-06 
0.0 1.4066 0 2.0 1e-06 
0.0 1.4067 0 2.0 1e-06 
0.0 1.4068 0 2.0 1e-06 
0.0 1.4069 0 2.0 1e-06 
0.0 1.407 0 2.0 1e-06 
0.0 1.4071 0 2.0 1e-06 
0.0 1.4072 0 2.0 1e-06 
0.0 1.4073 0 2.0 1e-06 
0.0 1.4074 0 2.0 1e-06 
0.0 1.4075 0 2.0 1e-06 
0.0 1.4076 0 2.0 1e-06 
0.0 1.4077 0 2.0 1e-06 
0.0 1.4078 0 2.0 1e-06 
0.0 1.4079 0 2.0 1e-06 
0.0 1.408 0 2.0 1e-06 
0.0 1.4081 0 2.0 1e-06 
0.0 1.4082 0 2.0 1e-06 
0.0 1.4083 0 2.0 1e-06 
0.0 1.4084 0 2.0 1e-06 
0.0 1.4085 0 2.0 1e-06 
0.0 1.4086 0 2.0 1e-06 
0.0 1.4087 0 2.0 1e-06 
0.0 1.4088 0 2.0 1e-06 
0.0 1.4089 0 2.0 1e-06 
0.0 1.409 0 2.0 1e-06 
0.0 1.4091 0 2.0 1e-06 
0.0 1.4092 0 2.0 1e-06 
0.0 1.4093 0 2.0 1e-06 
0.0 1.4094 0 2.0 1e-06 
0.0 1.4095 0 2.0 1e-06 
0.0 1.4096 0 2.0 1e-06 
0.0 1.4097 0 2.0 1e-06 
0.0 1.4098 0 2.0 1e-06 
0.0 1.4099 0 2.0 1e-06 
0.0 1.41 0 2.0 1e-06 
0.0 1.4101 0 2.0 1e-06 
0.0 1.4102 0 2.0 1e-06 
0.0 1.4103 0 2.0 1e-06 
0.0 1.4104 0 2.0 1e-06 
0.0 1.4105 0 2.0 1e-06 
0.0 1.4106 0 2.0 1e-06 
0.0 1.4107 0 2.0 1e-06 
0.0 1.4108 0 2.0 1e-06 
0.0 1.4109 0 2.0 1e-06 
0.0 1.411 0 2.0 1e-06 
0.0 1.4111 0 2.0 1e-06 
0.0 1.4112 0 2.0 1e-06 
0.0 1.4113 0 2.0 1e-06 
0.0 1.4114 0 2.0 1e-06 
0.0 1.4115 0 2.0 1e-06 
0.0 1.4116 0 2.0 1e-06 
0.0 1.4117 0 2.0 1e-06 
0.0 1.4118 0 2.0 1e-06 
0.0 1.4119 0 2.0 1e-06 
0.0 1.412 0 2.0 1e-06 
0.0 1.4121 0 2.0 1e-06 
0.0 1.4122 0 2.0 1e-06 
0.0 1.4123 0 2.0 1e-06 
0.0 1.4124 0 2.0 1e-06 
0.0 1.4125 0 2.0 1e-06 
0.0 1.4126 0 2.0 1e-06 
0.0 1.4127 0 2.0 1e-06 
0.0 1.4128 0 2.0 1e-06 
0.0 1.4129 0 2.0 1e-06 
0.0 1.413 0 2.0 1e-06 
0.0 1.4131 0 2.0 1e-06 
0.0 1.4132 0 2.0 1e-06 
0.0 1.4133 0 2.0 1e-06 
0.0 1.4134 0 2.0 1e-06 
0.0 1.4135 0 2.0 1e-06 
0.0 1.4136 0 2.0 1e-06 
0.0 1.4137 0 2.0 1e-06 
0.0 1.4138 0 2.0 1e-06 
0.0 1.4139 0 2.0 1e-06 
0.0 1.414 0 2.0 1e-06 
0.0 1.4141 0 2.0 1e-06 
0.0 1.4142 0 2.0 1e-06 
0.0 1.4143 0 2.0 1e-06 
0.0 1.4144 0 2.0 1e-06 
0.0 1.4145 0 2.0 1e-06 
0.0 1.4146 0 2.0 1e-06 
0.0 1.4147 0 2.0 1e-06 
0.0 1.4148 0 2.0 1e-06 
0.0 1.4149 0 2.0 1e-06 
0.0 1.415 0 2.0 1e-06 
0.0 1.4151 0 2.0 1e-06 
0.0 1.4152 0 2.0 1e-06 
0.0 1.4153 0 2.0 1e-06 
0.0 1.4154 0 2.0 1e-06 
0.0 1.4155 0 2.0 1e-06 
0.0 1.4156 0 2.0 1e-06 
0.0 1.4157 0 2.0 1e-06 
0.0 1.4158 0 2.0 1e-06 
0.0 1.4159 0 2.0 1e-06 
0.0 1.416 0 2.0 1e-06 
0.0 1.4161 0 2.0 1e-06 
0.0 1.4162 0 2.0 1e-06 
0.0 1.4163 0 2.0 1e-06 
0.0 1.4164 0 2.0 1e-06 
0.0 1.4165 0 2.0 1e-06 
0.0 1.4166 0 2.0 1e-06 
0.0 1.4167 0 2.0 1e-06 
0.0 1.4168 0 2.0 1e-06 
0.0 1.4169 0 2.0 1e-06 
0.0 1.417 0 2.0 1e-06 
0.0 1.4171 0 2.0 1e-06 
0.0 1.4172 0 2.0 1e-06 
0.0 1.4173 0 2.0 1e-06 
0.0 1.4174 0 2.0 1e-06 
0.0 1.4175 0 2.0 1e-06 
0.0 1.4176 0 2.0 1e-06 
0.0 1.4177 0 2.0 1e-06 
0.0 1.4178 0 2.0 1e-06 
0.0 1.4179 0 2.0 1e-06 
0.0 1.418 0 2.0 1e-06 
0.0 1.4181 0 2.0 1e-06 
0.0 1.4182 0 2.0 1e-06 
0.0 1.4183 0 2.0 1e-06 
0.0 1.4184 0 2.0 1e-06 
0.0 1.4185 0 2.0 1e-06 
0.0 1.4186 0 2.0 1e-06 
0.0 1.4187 0 2.0 1e-06 
0.0 1.4188 0 2.0 1e-06 
0.0 1.4189 0 2.0 1e-06 
0.0 1.419 0 2.0 1e-06 
0.0 1.4191 0 2.0 1e-06 
0.0 1.4192 0 2.0 1e-06 
0.0 1.4193 0 2.0 1e-06 
0.0 1.4194 0 2.0 1e-06 
0.0 1.4195 0 2.0 1e-06 
0.0 1.4196 0 2.0 1e-06 
0.0 1.4197 0 2.0 1e-06 
0.0 1.4198 0 2.0 1e-06 
0.0 1.4199 0 2.0 1e-06 
0.0 1.42 0 2.0 1e-06 
0.0 1.4201 0 2.0 1e-06 
0.0 1.4202 0 2.0 1e-06 
0.0 1.4203 0 2.0 1e-06 
0.0 1.4204 0 2.0 1e-06 
0.0 1.4205 0 2.0 1e-06 
0.0 1.4206 0 2.0 1e-06 
0.0 1.4207 0 2.0 1e-06 
0.0 1.4208 0 2.0 1e-06 
0.0 1.4209 0 2.0 1e-06 
0.0 1.421 0 2.0 1e-06 
0.0 1.4211 0 2.0 1e-06 
0.0 1.4212 0 2.0 1e-06 
0.0 1.4213 0 2.0 1e-06 
0.0 1.4214 0 2.0 1e-06 
0.0 1.4215 0 2.0 1e-06 
0.0 1.4216 0 2.0 1e-06 
0.0 1.4217 0 2.0 1e-06 
0.0 1.4218 0 2.0 1e-06 
0.0 1.4219 0 2.0 1e-06 
0.0 1.422 0 2.0 1e-06 
0.0 1.4221 0 2.0 1e-06 
0.0 1.4222 0 2.0 1e-06 
0.0 1.4223 0 2.0 1e-06 
0.0 1.4224 0 2.0 1e-06 
0.0 1.4225 0 2.0 1e-06 
0.0 1.4226 0 2.0 1e-06 
0.0 1.4227 0 2.0 1e-06 
0.0 1.4228 0 2.0 1e-06 
0.0 1.4229 0 2.0 1e-06 
0.0 1.423 0 2.0 1e-06 
0.0 1.4231 0 2.0 1e-06 
0.0 1.4232 0 2.0 1e-06 
0.0 1.4233 0 2.0 1e-06 
0.0 1.4234 0 2.0 1e-06 
0.0 1.4235 0 2.0 1e-06 
0.0 1.4236 0 2.0 1e-06 
0.0 1.4237 0 2.0 1e-06 
0.0 1.4238 0 2.0 1e-06 
0.0 1.4239 0 2.0 1e-06 
0.0 1.424 0 2.0 1e-06 
0.0 1.4241 0 2.0 1e-06 
0.0 1.4242 0 2.0 1e-06 
0.0 1.4243 0 2.0 1e-06 
0.0 1.4244 0 2.0 1e-06 
0.0 1.4245 0 2.0 1e-06 
0.0 1.4246 0 2.0 1e-06 
0.0 1.4247 0 2.0 1e-06 
0.0 1.4248 0 2.0 1e-06 
0.0 1.4249 0 2.0 1e-06 
0.0 1.425 0 2.0 1e-06 
0.0 1.4251 0 2.0 1e-06 
0.0 1.4252 0 2.0 1e-06 
0.0 1.4253 0 2.0 1e-06 
0.0 1.4254 0 2.0 1e-06 
0.0 1.4255 0 2.0 1e-06 
0.0 1.4256 0 2.0 1e-06 
0.0 1.4257 0 2.0 1e-06 
0.0 1.4258 0 2.0 1e-06 
0.0 1.4259 0 2.0 1e-06 
0.0 1.426 0 2.0 1e-06 
0.0 1.4261 0 2.0 1e-06 
0.0 1.4262 0 2.0 1e-06 
0.0 1.4263 0 2.0 1e-06 
0.0 1.4264 0 2.0 1e-06 
0.0 1.4265 0 2.0 1e-06 
0.0 1.4266 0 2.0 1e-06 
0.0 1.4267 0 2.0 1e-06 
0.0 1.4268 0 2.0 1e-06 
0.0 1.4269 0 2.0 1e-06 
0.0 1.427 0 2.0 1e-06 
0.0 1.4271 0 2.0 1e-06 
0.0 1.4272 0 2.0 1e-06 
0.0 1.4273 0 2.0 1e-06 
0.0 1.4274 0 2.0 1e-06 
0.0 1.4275 0 2.0 1e-06 
0.0 1.4276 0 2.0 1e-06 
0.0 1.4277 0 2.0 1e-06 
0.0 1.4278 0 2.0 1e-06 
0.0 1.4279 0 2.0 1e-06 
0.0 1.428 0 2.0 1e-06 
0.0 1.4281 0 2.0 1e-06 
0.0 1.4282 0 2.0 1e-06 
0.0 1.4283 0 2.0 1e-06 
0.0 1.4284 0 2.0 1e-06 
0.0 1.4285 0 2.0 1e-06 
0.0 1.4286 0 2.0 1e-06 
0.0 1.4287 0 2.0 1e-06 
0.0 1.4288 0 2.0 1e-06 
0.0 1.4289 0 2.0 1e-06 
0.0 1.429 0 2.0 1e-06 
0.0 1.4291 0 2.0 1e-06 
0.0 1.4292 0 2.0 1e-06 
0.0 1.4293 0 2.0 1e-06 
0.0 1.4294 0 2.0 1e-06 
0.0 1.4295 0 2.0 1e-06 
0.0 1.4296 0 2.0 1e-06 
0.0 1.4297 0 2.0 1e-06 
0.0 1.4298 0 2.0 1e-06 
0.0 1.4299 0 2.0 1e-06 
0.0 1.43 0 2.0 1e-06 
0.0 1.4301 0 2.0 1e-06 
0.0 1.4302 0 2.0 1e-06 
0.0 1.4303 0 2.0 1e-06 
0.0 1.4304 0 2.0 1e-06 
0.0 1.4305 0 2.0 1e-06 
0.0 1.4306 0 2.0 1e-06 
0.0 1.4307 0 2.0 1e-06 
0.0 1.4308 0 2.0 1e-06 
0.0 1.4309 0 2.0 1e-06 
0.0 1.431 0 2.0 1e-06 
0.0 1.4311 0 2.0 1e-06 
0.0 1.4312 0 2.0 1e-06 
0.0 1.4313 0 2.0 1e-06 
0.0 1.4314 0 2.0 1e-06 
0.0 1.4315 0 2.0 1e-06 
0.0 1.4316 0 2.0 1e-06 
0.0 1.4317 0 2.0 1e-06 
0.0 1.4318 0 2.0 1e-06 
0.0 1.4319 0 2.0 1e-06 
0.0 1.432 0 2.0 1e-06 
0.0 1.4321 0 2.0 1e-06 
0.0 1.4322 0 2.0 1e-06 
0.0 1.4323 0 2.0 1e-06 
0.0 1.4324 0 2.0 1e-06 
0.0 1.4325 0 2.0 1e-06 
0.0 1.4326 0 2.0 1e-06 
0.0 1.4327 0 2.0 1e-06 
0.0 1.4328 0 2.0 1e-06 
0.0 1.4329 0 2.0 1e-06 
0.0 1.433 0 2.0 1e-06 
0.0 1.4331 0 2.0 1e-06 
0.0 1.4332 0 2.0 1e-06 
0.0 1.4333 0 2.0 1e-06 
0.0 1.4334 0 2.0 1e-06 
0.0 1.4335 0 2.0 1e-06 
0.0 1.4336 0 2.0 1e-06 
0.0 1.4337 0 2.0 1e-06 
0.0 1.4338 0 2.0 1e-06 
0.0 1.4339 0 2.0 1e-06 
0.0 1.434 0 2.0 1e-06 
0.0 1.4341 0 2.0 1e-06 
0.0 1.4342 0 2.0 1e-06 
0.0 1.4343 0 2.0 1e-06 
0.0 1.4344 0 2.0 1e-06 
0.0 1.4345 0 2.0 1e-06 
0.0 1.4346 0 2.0 1e-06 
0.0 1.4347 0 2.0 1e-06 
0.0 1.4348 0 2.0 1e-06 
0.0 1.4349 0 2.0 1e-06 
0.0 1.435 0 2.0 1e-06 
0.0 1.4351 0 2.0 1e-06 
0.0 1.4352 0 2.0 1e-06 
0.0 1.4353 0 2.0 1e-06 
0.0 1.4354 0 2.0 1e-06 
0.0 1.4355 0 2.0 1e-06 
0.0 1.4356 0 2.0 1e-06 
0.0 1.4357 0 2.0 1e-06 
0.0 1.4358 0 2.0 1e-06 
0.0 1.4359 0 2.0 1e-06 
0.0 1.436 0 2.0 1e-06 
0.0 1.4361 0 2.0 1e-06 
0.0 1.4362 0 2.0 1e-06 
0.0 1.4363 0 2.0 1e-06 
0.0 1.4364 0 2.0 1e-06 
0.0 1.4365 0 2.0 1e-06 
0.0 1.4366 0 2.0 1e-06 
0.0 1.4367 0 2.0 1e-06 
0.0 1.4368 0 2.0 1e-06 
0.0 1.4369 0 2.0 1e-06 
0.0 1.437 0 2.0 1e-06 
0.0 1.4371 0 2.0 1e-06 
0.0 1.4372 0 2.0 1e-06 
0.0 1.4373 0 2.0 1e-06 
0.0 1.4374 0 2.0 1e-06 
0.0 1.4375 0 2.0 1e-06 
0.0 1.4376 0 2.0 1e-06 
0.0 1.4377 0 2.0 1e-06 
0.0 1.4378 0 2.0 1e-06 
0.0 1.4379 0 2.0 1e-06 
0.0 1.438 0 2.0 1e-06 
0.0 1.4381 0 2.0 1e-06 
0.0 1.4382 0 2.0 1e-06 
0.0 1.4383 0 2.0 1e-06 
0.0 1.4384 0 2.0 1e-06 
0.0 1.4385 0 2.0 1e-06 
0.0 1.4386 0 2.0 1e-06 
0.0 1.4387 0 2.0 1e-06 
0.0 1.4388 0 2.0 1e-06 
0.0 1.4389 0 2.0 1e-06 
0.0 1.439 0 2.0 1e-06 
0.0 1.4391 0 2.0 1e-06 
0.0 1.4392 0 2.0 1e-06 
0.0 1.4393 0 2.0 1e-06 
0.0 1.4394 0 2.0 1e-06 
0.0 1.4395 0 2.0 1e-06 
0.0 1.4396 0 2.0 1e-06 
0.0 1.4397 0 2.0 1e-06 
0.0 1.4398 0 2.0 1e-06 
0.0 1.4399 0 2.0 1e-06 
0.0 1.44 0 2.0 1e-06 
0.0 1.4401 0 2.0 1e-06 
0.0 1.4402 0 2.0 1e-06 
0.0 1.4403 0 2.0 1e-06 
0.0 1.4404 0 2.0 1e-06 
0.0 1.4405 0 2.0 1e-06 
0.0 1.4406 0 2.0 1e-06 
0.0 1.4407 0 2.0 1e-06 
0.0 1.4408 0 2.0 1e-06 
0.0 1.4409 0 2.0 1e-06 
0.0 1.441 0 2.0 1e-06 
0.0 1.4411 0 2.0 1e-06 
0.0 1.4412 0 2.0 1e-06 
0.0 1.4413 0 2.0 1e-06 
0.0 1.4414 0 2.0 1e-06 
0.0 1.4415 0 2.0 1e-06 
0.0 1.4416 0 2.0 1e-06 
0.0 1.4417 0 2.0 1e-06 
0.0 1.4418 0 2.0 1e-06 
0.0 1.4419 0 2.0 1e-06 
0.0 1.442 0 2.0 1e-06 
0.0 1.4421 0 2.0 1e-06 
0.0 1.4422 0 2.0 1e-06 
0.0 1.4423 0 2.0 1e-06 
0.0 1.4424 0 2.0 1e-06 
0.0 1.4425 0 2.0 1e-06 
0.0 1.4426 0 2.0 1e-06 
0.0 1.4427 0 2.0 1e-06 
0.0 1.4428 0 2.0 1e-06 
0.0 1.4429 0 2.0 1e-06 
0.0 1.443 0 2.0 1e-06 
0.0 1.4431 0 2.0 1e-06 
0.0 1.4432 0 2.0 1e-06 
0.0 1.4433 0 2.0 1e-06 
0.0 1.4434 0 2.0 1e-06 
0.0 1.4435 0 2.0 1e-06 
0.0 1.4436 0 2.0 1e-06 
0.0 1.4437 0 2.0 1e-06 
0.0 1.4438 0 2.0 1e-06 
0.0 1.4439 0 2.0 1e-06 
0.0 1.444 0 2.0 1e-06 
0.0 1.4441 0 2.0 1e-06 
0.0 1.4442 0 2.0 1e-06 
0.0 1.4443 0 2.0 1e-06 
0.0 1.4444 0 2.0 1e-06 
0.0 1.4445 0 2.0 1e-06 
0.0 1.4446 0 2.0 1e-06 
0.0 1.4447 0 2.0 1e-06 
0.0 1.4448 0 2.0 1e-06 
0.0 1.4449 0 2.0 1e-06 
0.0 1.445 0 2.0 1e-06 
0.0 1.4451 0 2.0 1e-06 
0.0 1.4452 0 2.0 1e-06 
0.0 1.4453 0 2.0 1e-06 
0.0 1.4454 0 2.0 1e-06 
0.0 1.4455 0 2.0 1e-06 
0.0 1.4456 0 2.0 1e-06 
0.0 1.4457 0 2.0 1e-06 
0.0 1.4458 0 2.0 1e-06 
0.0 1.4459 0 2.0 1e-06 
0.0 1.446 0 2.0 1e-06 
0.0 1.4461 0 2.0 1e-06 
0.0 1.4462 0 2.0 1e-06 
0.0 1.4463 0 2.0 1e-06 
0.0 1.4464 0 2.0 1e-06 
0.0 1.4465 0 2.0 1e-06 
0.0 1.4466 0 2.0 1e-06 
0.0 1.4467 0 2.0 1e-06 
0.0 1.4468 0 2.0 1e-06 
0.0 1.4469 0 2.0 1e-06 
0.0 1.447 0 2.0 1e-06 
0.0 1.4471 0 2.0 1e-06 
0.0 1.4472 0 2.0 1e-06 
0.0 1.4473 0 2.0 1e-06 
0.0 1.4474 0 2.0 1e-06 
0.0 1.4475 0 2.0 1e-06 
0.0 1.4476 0 2.0 1e-06 
0.0 1.4477 0 2.0 1e-06 
0.0 1.4478 0 2.0 1e-06 
0.0 1.4479 0 2.0 1e-06 
0.0 1.448 0 2.0 1e-06 
0.0 1.4481 0 2.0 1e-06 
0.0 1.4482 0 2.0 1e-06 
0.0 1.4483 0 2.0 1e-06 
0.0 1.4484 0 2.0 1e-06 
0.0 1.4485 0 2.0 1e-06 
0.0 1.4486 0 2.0 1e-06 
0.0 1.4487 0 2.0 1e-06 
0.0 1.4488 0 2.0 1e-06 
0.0 1.4489 0 2.0 1e-06 
0.0 1.449 0 2.0 1e-06 
0.0 1.4491 0 2.0 1e-06 
0.0 1.4492 0 2.0 1e-06 
0.0 1.4493 0 2.0 1e-06 
0.0 1.4494 0 2.0 1e-06 
0.0 1.4495 0 2.0 1e-06 
0.0 1.4496 0 2.0 1e-06 
0.0 1.4497 0 2.0 1e-06 
0.0 1.4498 0 2.0 1e-06 
0.0 1.4499 0 2.0 1e-06 
0.0 1.45 0 2.0 1e-06 
0.0 1.4501 0 2.0 1e-06 
0.0 1.4502 0 2.0 1e-06 
0.0 1.4503 0 2.0 1e-06 
0.0 1.4504 0 2.0 1e-06 
0.0 1.4505 0 2.0 1e-06 
0.0 1.4506 0 2.0 1e-06 
0.0 1.4507 0 2.0 1e-06 
0.0 1.4508 0 2.0 1e-06 
0.0 1.4509 0 2.0 1e-06 
0.0 1.451 0 2.0 1e-06 
0.0 1.4511 0 2.0 1e-06 
0.0 1.4512 0 2.0 1e-06 
0.0 1.4513 0 2.0 1e-06 
0.0 1.4514 0 2.0 1e-06 
0.0 1.4515 0 2.0 1e-06 
0.0 1.4516 0 2.0 1e-06 
0.0 1.4517 0 2.0 1e-06 
0.0 1.4518 0 2.0 1e-06 
0.0 1.4519 0 2.0 1e-06 
0.0 1.452 0 2.0 1e-06 
0.0 1.4521 0 2.0 1e-06 
0.0 1.4522 0 2.0 1e-06 
0.0 1.4523 0 2.0 1e-06 
0.0 1.4524 0 2.0 1e-06 
0.0 1.4525 0 2.0 1e-06 
0.0 1.4526 0 2.0 1e-06 
0.0 1.4527 0 2.0 1e-06 
0.0 1.4528 0 2.0 1e-06 
0.0 1.4529 0 2.0 1e-06 
0.0 1.453 0 2.0 1e-06 
0.0 1.4531 0 2.0 1e-06 
0.0 1.4532 0 2.0 1e-06 
0.0 1.4533 0 2.0 1e-06 
0.0 1.4534 0 2.0 1e-06 
0.0 1.4535 0 2.0 1e-06 
0.0 1.4536 0 2.0 1e-06 
0.0 1.4537 0 2.0 1e-06 
0.0 1.4538 0 2.0 1e-06 
0.0 1.4539 0 2.0 1e-06 
0.0 1.454 0 2.0 1e-06 
0.0 1.4541 0 2.0 1e-06 
0.0 1.4542 0 2.0 1e-06 
0.0 1.4543 0 2.0 1e-06 
0.0 1.4544 0 2.0 1e-06 
0.0 1.4545 0 2.0 1e-06 
0.0 1.4546 0 2.0 1e-06 
0.0 1.4547 0 2.0 1e-06 
0.0 1.4548 0 2.0 1e-06 
0.0 1.4549 0 2.0 1e-06 
0.0 1.455 0 2.0 1e-06 
0.0 1.4551 0 2.0 1e-06 
0.0 1.4552 0 2.0 1e-06 
0.0 1.4553 0 2.0 1e-06 
0.0 1.4554 0 2.0 1e-06 
0.0 1.4555 0 2.0 1e-06 
0.0 1.4556 0 2.0 1e-06 
0.0 1.4557 0 2.0 1e-06 
0.0 1.4558 0 2.0 1e-06 
0.0 1.4559 0 2.0 1e-06 
0.0 1.456 0 2.0 1e-06 
0.0 1.4561 0 2.0 1e-06 
0.0 1.4562 0 2.0 1e-06 
0.0 1.4563 0 2.0 1e-06 
0.0 1.4564 0 2.0 1e-06 
0.0 1.4565 0 2.0 1e-06 
0.0 1.4566 0 2.0 1e-06 
0.0 1.4567 0 2.0 1e-06 
0.0 1.4568 0 2.0 1e-06 
0.0 1.4569 0 2.0 1e-06 
0.0 1.457 0 2.0 1e-06 
0.0 1.4571 0 2.0 1e-06 
0.0 1.4572 0 2.0 1e-06 
0.0 1.4573 0 2.0 1e-06 
0.0 1.4574 0 2.0 1e-06 
0.0 1.4575 0 2.0 1e-06 
0.0 1.4576 0 2.0 1e-06 
0.0 1.4577 0 2.0 1e-06 
0.0 1.4578 0 2.0 1e-06 
0.0 1.4579 0 2.0 1e-06 
0.0 1.458 0 2.0 1e-06 
0.0 1.4581 0 2.0 1e-06 
0.0 1.4582 0 2.0 1e-06 
0.0 1.4583 0 2.0 1e-06 
0.0 1.4584 0 2.0 1e-06 
0.0 1.4585 0 2.0 1e-06 
0.0 1.4586 0 2.0 1e-06 
0.0 1.4587 0 2.0 1e-06 
0.0 1.4588 0 2.0 1e-06 
0.0 1.4589 0 2.0 1e-06 
0.0 1.459 0 2.0 1e-06 
0.0 1.4591 0 2.0 1e-06 
0.0 1.4592 0 2.0 1e-06 
0.0 1.4593 0 2.0 1e-06 
0.0 1.4594 0 2.0 1e-06 
0.0 1.4595 0 2.0 1e-06 
0.0 1.4596 0 2.0 1e-06 
0.0 1.4597 0 2.0 1e-06 
0.0 1.4598 0 2.0 1e-06 
0.0 1.4599 0 2.0 1e-06 
0.0 1.46 0 2.0 1e-06 
0.0 1.4601 0 2.0 1e-06 
0.0 1.4602 0 2.0 1e-06 
0.0 1.4603 0 2.0 1e-06 
0.0 1.4604 0 2.0 1e-06 
0.0 1.4605 0 2.0 1e-06 
0.0 1.4606 0 2.0 1e-06 
0.0 1.4607 0 2.0 1e-06 
0.0 1.4608 0 2.0 1e-06 
0.0 1.4609 0 2.0 1e-06 
0.0 1.461 0 2.0 1e-06 
0.0 1.4611 0 2.0 1e-06 
0.0 1.4612 0 2.0 1e-06 
0.0 1.4613 0 2.0 1e-06 
0.0 1.4614 0 2.0 1e-06 
0.0 1.4615 0 2.0 1e-06 
0.0 1.4616 0 2.0 1e-06 
0.0 1.4617 0 2.0 1e-06 
0.0 1.4618 0 2.0 1e-06 
0.0 1.4619 0 2.0 1e-06 
0.0 1.462 0 2.0 1e-06 
0.0 1.4621 0 2.0 1e-06 
0.0 1.4622 0 2.0 1e-06 
0.0 1.4623 0 2.0 1e-06 
0.0 1.4624 0 2.0 1e-06 
0.0 1.4625 0 2.0 1e-06 
0.0 1.4626 0 2.0 1e-06 
0.0 1.4627 0 2.0 1e-06 
0.0 1.4628 0 2.0 1e-06 
0.0 1.4629 0 2.0 1e-06 
0.0 1.463 0 2.0 1e-06 
0.0 1.4631 0 2.0 1e-06 
0.0 1.4632 0 2.0 1e-06 
0.0 1.4633 0 2.0 1e-06 
0.0 1.4634 0 2.0 1e-06 
0.0 1.4635 0 2.0 1e-06 
0.0 1.4636 0 2.0 1e-06 
0.0 1.4637 0 2.0 1e-06 
0.0 1.4638 0 2.0 1e-06 
0.0 1.4639 0 2.0 1e-06 
0.0 1.464 0 2.0 1e-06 
0.0 1.4641 0 2.0 1e-06 
0.0 1.4642 0 2.0 1e-06 
0.0 1.4643 0 2.0 1e-06 
0.0 1.4644 0 2.0 1e-06 
0.0 1.4645 0 2.0 1e-06 
0.0 1.4646 0 2.0 1e-06 
0.0 1.4647 0 2.0 1e-06 
0.0 1.4648 0 2.0 1e-06 
0.0 1.4649 0 2.0 1e-06 
0.0 1.465 0 2.0 1e-06 
0.0 1.4651 0 2.0 1e-06 
0.0 1.4652 0 2.0 1e-06 
0.0 1.4653 0 2.0 1e-06 
0.0 1.4654 0 2.0 1e-06 
0.0 1.4655 0 2.0 1e-06 
0.0 1.4656 0 2.0 1e-06 
0.0 1.4657 0 2.0 1e-06 
0.0 1.4658 0 2.0 1e-06 
0.0 1.4659 0 2.0 1e-06 
0.0 1.466 0 2.0 1e-06 
0.0 1.4661 0 2.0 1e-06 
0.0 1.4662 0 2.0 1e-06 
0.0 1.4663 0 2.0 1e-06 
0.0 1.4664 0 2.0 1e-06 
0.0 1.4665 0 2.0 1e-06 
0.0 1.4666 0 2.0 1e-06 
0.0 1.4667 0 2.0 1e-06 
0.0 1.4668 0 2.0 1e-06 
0.0 1.4669 0 2.0 1e-06 
0.0 1.467 0 2.0 1e-06 
0.0 1.4671 0 2.0 1e-06 
0.0 1.4672 0 2.0 1e-06 
0.0 1.4673 0 2.0 1e-06 
0.0 1.4674 0 2.0 1e-06 
0.0 1.4675 0 2.0 1e-06 
0.0 1.4676 0 2.0 1e-06 
0.0 1.4677 0 2.0 1e-06 
0.0 1.4678 0 2.0 1e-06 
0.0 1.4679 0 2.0 1e-06 
0.0 1.468 0 2.0 1e-06 
0.0 1.4681 0 2.0 1e-06 
0.0 1.4682 0 2.0 1e-06 
0.0 1.4683 0 2.0 1e-06 
0.0 1.4684 0 2.0 1e-06 
0.0 1.4685 0 2.0 1e-06 
0.0 1.4686 0 2.0 1e-06 
0.0 1.4687 0 2.0 1e-06 
0.0 1.4688 0 2.0 1e-06 
0.0 1.4689 0 2.0 1e-06 
0.0 1.469 0 2.0 1e-06 
0.0 1.4691 0 2.0 1e-06 
0.0 1.4692 0 2.0 1e-06 
0.0 1.4693 0 2.0 1e-06 
0.0 1.4694 0 2.0 1e-06 
0.0 1.4695 0 2.0 1e-06 
0.0 1.4696 0 2.0 1e-06 
0.0 1.4697 0 2.0 1e-06 
0.0 1.4698 0 2.0 1e-06 
0.0 1.4699 0 2.0 1e-06 
0.0 1.47 0 2.0 1e-06 
0.0 1.4701 0 2.0 1e-06 
0.0 1.4702 0 2.0 1e-06 
0.0 1.4703 0 2.0 1e-06 
0.0 1.4704 0 2.0 1e-06 
0.0 1.4705 0 2.0 1e-06 
0.0 1.4706 0 2.0 1e-06 
0.0 1.4707 0 2.0 1e-06 
0.0 1.4708 0 2.0 1e-06 
0.0 1.4709 0 2.0 1e-06 
0.0 1.471 0 2.0 1e-06 
0.0 1.4711 0 2.0 1e-06 
0.0 1.4712 0 2.0 1e-06 
0.0 1.4713 0 2.0 1e-06 
0.0 1.4714 0 2.0 1e-06 
0.0 1.4715 0 2.0 1e-06 
0.0 1.4716 0 2.0 1e-06 
0.0 1.4717 0 2.0 1e-06 
0.0 1.4718 0 2.0 1e-06 
0.0 1.4719 0 2.0 1e-06 
0.0 1.472 0 2.0 1e-06 
0.0 1.4721 0 2.0 1e-06 
0.0 1.4722 0 2.0 1e-06 
0.0 1.4723 0 2.0 1e-06 
0.0 1.4724 0 2.0 1e-06 
0.0 1.4725 0 2.0 1e-06 
0.0 1.4726 0 2.0 1e-06 
0.0 1.4727 0 2.0 1e-06 
0.0 1.4728 0 2.0 1e-06 
0.0 1.4729 0 2.0 1e-06 
0.0 1.473 0 2.0 1e-06 
0.0 1.4731 0 2.0 1e-06 
0.0 1.4732 0 2.0 1e-06 
0.0 1.4733 0 2.0 1e-06 
0.0 1.4734 0 2.0 1e-06 
0.0 1.4735 0 2.0 1e-06 
0.0 1.4736 0 2.0 1e-06 
0.0 1.4737 0 2.0 1e-06 
0.0 1.4738 0 2.0 1e-06 
0.0 1.4739 0 2.0 1e-06 
0.0 1.474 0 2.0 1e-06 
0.0 1.4741 0 2.0 1e-06 
0.0 1.4742 0 2.0 1e-06 
0.0 1.4743 0 2.0 1e-06 
0.0 1.4744 0 2.0 1e-06 
0.0 1.4745 0 2.0 1e-06 
0.0 1.4746 0 2.0 1e-06 
0.0 1.4747 0 2.0 1e-06 
0.0 1.4748 0 2.0 1e-06 
0.0 1.4749 0 2.0 1e-06 
0.0 1.475 0 2.0 1e-06 
0.0 1.4751 0 2.0 1e-06 
0.0 1.4752 0 2.0 1e-06 
0.0 1.4753 0 2.0 1e-06 
0.0 1.4754 0 2.0 1e-06 
0.0 1.4755 0 2.0 1e-06 
0.0 1.4756 0 2.0 1e-06 
0.0 1.4757 0 2.0 1e-06 
0.0 1.4758 0 2.0 1e-06 
0.0 1.4759 0 2.0 1e-06 
0.0 1.476 0 2.0 1e-06 
0.0 1.4761 0 2.0 1e-06 
0.0 1.4762 0 2.0 1e-06 
0.0 1.4763 0 2.0 1e-06 
0.0 1.4764 0 2.0 1e-06 
0.0 1.4765 0 2.0 1e-06 
0.0 1.4766 0 2.0 1e-06 
0.0 1.4767 0 2.0 1e-06 
0.0 1.4768 0 2.0 1e-06 
0.0 1.4769 0 2.0 1e-06 
0.0 1.477 0 2.0 1e-06 
0.0 1.4771 0 2.0 1e-06 
0.0 1.4772 0 2.0 1e-06 
0.0 1.4773 0 2.0 1e-06 
0.0 1.4774 0 2.0 1e-06 
0.0 1.4775 0 2.0 1e-06 
0.0 1.4776 0 2.0 1e-06 
0.0 1.4777 0 2.0 1e-06 
0.0 1.4778 0 2.0 1e-06 
0.0 1.4779 0 2.0 1e-06 
0.0 1.478 0 2.0 1e-06 
0.0 1.4781 0 2.0 1e-06 
0.0 1.4782 0 2.0 1e-06 
0.0 1.4783 0 2.0 1e-06 
0.0 1.4784 0 2.0 1e-06 
0.0 1.4785 0 2.0 1e-06 
0.0 1.4786 0 2.0 1e-06 
0.0 1.4787 0 2.0 1e-06 
0.0 1.4788 0 2.0 1e-06 
0.0 1.4789 0 2.0 1e-06 
0.0 1.479 0 2.0 1e-06 
0.0 1.4791 0 2.0 1e-06 
0.0 1.4792 0 2.0 1e-06 
0.0 1.4793 0 2.0 1e-06 
0.0 1.4794 0 2.0 1e-06 
0.0 1.4795 0 2.0 1e-06 
0.0 1.4796 0 2.0 1e-06 
0.0 1.4797 0 2.0 1e-06 
0.0 1.4798 0 2.0 1e-06 
0.0 1.4799 0 2.0 1e-06 
0.0 1.48 0 2.0 1e-06 
0.0 1.4801 0 2.0 1e-06 
0.0 1.4802 0 2.0 1e-06 
0.0 1.4803 0 2.0 1e-06 
0.0 1.4804 0 2.0 1e-06 
0.0 1.4805 0 2.0 1e-06 
0.0 1.4806 0 2.0 1e-06 
0.0 1.4807 0 2.0 1e-06 
0.0 1.4808 0 2.0 1e-06 
0.0 1.4809 0 2.0 1e-06 
0.0 1.481 0 2.0 1e-06 
0.0 1.4811 0 2.0 1e-06 
0.0 1.4812 0 2.0 1e-06 
0.0 1.4813 0 2.0 1e-06 
0.0 1.4814 0 2.0 1e-06 
0.0 1.4815 0 2.0 1e-06 
0.0 1.4816 0 2.0 1e-06 
0.0 1.4817 0 2.0 1e-06 
0.0 1.4818 0 2.0 1e-06 
0.0 1.4819 0 2.0 1e-06 
0.0 1.482 0 2.0 1e-06 
0.0 1.4821 0 2.0 1e-06 
0.0 1.4822 0 2.0 1e-06 
0.0 1.4823 0 2.0 1e-06 
0.0 1.4824 0 2.0 1e-06 
0.0 1.4825 0 2.0 1e-06 
0.0 1.4826 0 2.0 1e-06 
0.0 1.4827 0 2.0 1e-06 
0.0 1.4828 0 2.0 1e-06 
0.0 1.4829 0 2.0 1e-06 
0.0 1.483 0 2.0 1e-06 
0.0 1.4831 0 2.0 1e-06 
0.0 1.4832 0 2.0 1e-06 
0.0 1.4833 0 2.0 1e-06 
0.0 1.4834 0 2.0 1e-06 
0.0 1.4835 0 2.0 1e-06 
0.0 1.4836 0 2.0 1e-06 
0.0 1.4837 0 2.0 1e-06 
0.0 1.4838 0 2.0 1e-06 
0.0 1.4839 0 2.0 1e-06 
0.0 1.484 0 2.0 1e-06 
0.0 1.4841 0 2.0 1e-06 
0.0 1.4842 0 2.0 1e-06 
0.0 1.4843 0 2.0 1e-06 
0.0 1.4844 0 2.0 1e-06 
0.0 1.4845 0 2.0 1e-06 
0.0 1.4846 0 2.0 1e-06 
0.0 1.4847 0 2.0 1e-06 
0.0 1.4848 0 2.0 1e-06 
0.0 1.4849 0 2.0 1e-06 
0.0 1.485 0 2.0 1e-06 
0.0 1.4851 0 2.0 1e-06 
0.0 1.4852 0 2.0 1e-06 
0.0 1.4853 0 2.0 1e-06 
0.0 1.4854 0 2.0 1e-06 
0.0 1.4855 0 2.0 1e-06 
0.0 1.4856 0 2.0 1e-06 
0.0 1.4857 0 2.0 1e-06 
0.0 1.4858 0 2.0 1e-06 
0.0 1.4859 0 2.0 1e-06 
0.0 1.486 0 2.0 1e-06 
0.0 1.4861 0 2.0 1e-06 
0.0 1.4862 0 2.0 1e-06 
0.0 1.4863 0 2.0 1e-06 
0.0 1.4864 0 2.0 1e-06 
0.0 1.4865 0 2.0 1e-06 
0.0 1.4866 0 2.0 1e-06 
0.0 1.4867 0 2.0 1e-06 
0.0 1.4868 0 2.0 1e-06 
0.0 1.4869 0 2.0 1e-06 
0.0 1.487 0 2.0 1e-06 
0.0 1.4871 0 2.0 1e-06 
0.0 1.4872 0 2.0 1e-06 
0.0 1.4873 0 2.0 1e-06 
0.0 1.4874 0 2.0 1e-06 
0.0 1.4875 0 2.0 1e-06 
0.0 1.4876 0 2.0 1e-06 
0.0 1.4877 0 2.0 1e-06 
0.0 1.4878 0 2.0 1e-06 
0.0 1.4879 0 2.0 1e-06 
0.0 1.488 0 2.0 1e-06 
0.0 1.4881 0 2.0 1e-06 
0.0 1.4882 0 2.0 1e-06 
0.0 1.4883 0 2.0 1e-06 
0.0 1.4884 0 2.0 1e-06 
0.0 1.4885 0 2.0 1e-06 
0.0 1.4886 0 2.0 1e-06 
0.0 1.4887 0 2.0 1e-06 
0.0 1.4888 0 2.0 1e-06 
0.0 1.4889 0 2.0 1e-06 
0.0 1.489 0 2.0 1e-06 
0.0 1.4891 0 2.0 1e-06 
0.0 1.4892 0 2.0 1e-06 
0.0 1.4893 0 2.0 1e-06 
0.0 1.4894 0 2.0 1e-06 
0.0 1.4895 0 2.0 1e-06 
0.0 1.4896 0 2.0 1e-06 
0.0 1.4897 0 2.0 1e-06 
0.0 1.4898 0 2.0 1e-06 
0.0 1.4899 0 2.0 1e-06 
0.0 1.49 0 2.0 1e-06 
0.0 1.4901 0 2.0 1e-06 
0.0 1.4902 0 2.0 1e-06 
0.0 1.4903 0 2.0 1e-06 
0.0 1.4904 0 2.0 1e-06 
0.0 1.4905 0 2.0 1e-06 
0.0 1.4906 0 2.0 1e-06 
0.0 1.4907 0 2.0 1e-06 
0.0 1.4908 0 2.0 1e-06 
0.0 1.4909 0 2.0 1e-06 
0.0 1.491 0 2.0 1e-06 
0.0 1.4911 0 2.0 1e-06 
0.0 1.4912 0 2.0 1e-06 
0.0 1.4913 0 2.0 1e-06 
0.0 1.4914 0 2.0 1e-06 
0.0 1.4915 0 2.0 1e-06 
0.0 1.4916 0 2.0 1e-06 
0.0 1.4917 0 2.0 1e-06 
0.0 1.4918 0 2.0 1e-06 
0.0 1.4919 0 2.0 1e-06 
0.0 1.492 0 2.0 1e-06 
0.0 1.4921 0 2.0 1e-06 
0.0 1.4922 0 2.0 1e-06 
0.0 1.4923 0 2.0 1e-06 
0.0 1.4924 0 2.0 1e-06 
0.0 1.4925 0 2.0 1e-06 
0.0 1.4926 0 2.0 1e-06 
0.0 1.4927 0 2.0 1e-06 
0.0 1.4928 0 2.0 1e-06 
0.0 1.4929 0 2.0 1e-06 
0.0 1.493 0 2.0 1e-06 
0.0 1.4931 0 2.0 1e-06 
0.0 1.4932 0 2.0 1e-06 
0.0 1.4933 0 2.0 1e-06 
0.0 1.4934 0 2.0 1e-06 
0.0 1.4935 0 2.0 1e-06 
0.0 1.4936 0 2.0 1e-06 
0.0 1.4937 0 2.0 1e-06 
0.0 1.4938 0 2.0 1e-06 
0.0 1.4939 0 2.0 1e-06 
0.0 1.494 0 2.0 1e-06 
0.0 1.4941 0 2.0 1e-06 
0.0 1.4942 0 2.0 1e-06 
0.0 1.4943 0 2.0 1e-06 
0.0 1.4944 0 2.0 1e-06 
0.0 1.4945 0 2.0 1e-06 
0.0 1.4946 0 2.0 1e-06 
0.0 1.4947 0 2.0 1e-06 
0.0 1.4948 0 2.0 1e-06 
0.0 1.4949 0 2.0 1e-06 
0.0 1.495 0 2.0 1e-06 
0.0 1.4951 0 2.0 1e-06 
0.0 1.4952 0 2.0 1e-06 
0.0 1.4953 0 2.0 1e-06 
0.0 1.4954 0 2.0 1e-06 
0.0 1.4955 0 2.0 1e-06 
0.0 1.4956 0 2.0 1e-06 
0.0 1.4957 0 2.0 1e-06 
0.0 1.4958 0 2.0 1e-06 
0.0 1.4959 0 2.0 1e-06 
0.0 1.496 0 2.0 1e-06 
0.0 1.4961 0 2.0 1e-06 
0.0 1.4962 0 2.0 1e-06 
0.0 1.4963 0 2.0 1e-06 
0.0 1.4964 0 2.0 1e-06 
0.0 1.4965 0 2.0 1e-06 
0.0 1.4966 0 2.0 1e-06 
0.0 1.4967 0 2.0 1e-06 
0.0 1.4968 0 2.0 1e-06 
0.0 1.4969 0 2.0 1e-06 
0.0 1.497 0 2.0 1e-06 
0.0 1.4971 0 2.0 1e-06 
0.0 1.4972 0 2.0 1e-06 
0.0 1.4973 0 2.0 1e-06 
0.0 1.4974 0 2.0 1e-06 
0.0 1.4975 0 2.0 1e-06 
0.0 1.4976 0 2.0 1e-06 
0.0 1.4977 0 2.0 1e-06 
0.0 1.4978 0 2.0 1e-06 
0.0 1.4979 0 2.0 1e-06 
0.0 1.498 0 2.0 1e-06 
0.0 1.4981 0 2.0 1e-06 
0.0 1.4982 0 2.0 1e-06 
0.0 1.4983 0 2.0 1e-06 
0.0 1.4984 0 2.0 1e-06 
0.0 1.4985 0 2.0 1e-06 
0.0 1.4986 0 2.0 1e-06 
0.0 1.4987 0 2.0 1e-06 
0.0 1.4988 0 2.0 1e-06 
0.0 1.4989 0 2.0 1e-06 
0.0 1.499 0 2.0 1e-06 
0.0 1.4991 0 2.0 1e-06 
0.0 1.4992 0 2.0 1e-06 
0.0 1.4993 0 2.0 1e-06 
0.0 1.4994 0 2.0 1e-06 
0.0 1.4995 0 2.0 1e-06 
0.0 1.4996 0 2.0 1e-06 
0.0 1.4997 0 2.0 1e-06 
0.0 1.4998 0 2.0 1e-06 
0.0 1.4999 0 2.0 1e-06 
.ENDDATA 
.dc sweep DATA = datadc 
.print dc X1:IDS X1:qicores X1:qicored X1:ids0 X1:qfronts X1:qbacks X1:CFGDI X1:CFGSI 
.end