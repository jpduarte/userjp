*script to generate hspice simulation using cmdp, Juan Duarte 
*Date: 10/13/2015, time: 23:13:04

.option abstol=1e-6 reltol=1e-6 post ingold 
.option measform=1 
.temp 27 

.hdl "/users/jpduarte/research/BSIMIMG/code/bsimimg.va" 
.include "/users/jpduarte/research/userjp/project4/modelcards/modelcardsimple.nmos" 

.PARAM Vd_value = 0 
.PARAM Vgf_value = 0 
.PARAM Vs_value = 0 
.PARAM Vgb_value = 0 
.PARAM L_value = 5.5e-08 

Vd Vd 0.0 dc = Vd_value 
Vgf Vgf 0.0 dc = Vgf_value 
Vs Vs 0.0 dc = Vs_value 
Vgb Vgb 0.0 dc = Vgb_value 

X1 Vd Vgf Vs Vgb nmos1 L = 'L_value'

.DATA datadc Vd_value Vgf_value Vs_value Vgb_value L_value 
1.0 -1.5 0 5.0 5.5e-08 
1.0 -1.48 0 5.0 5.5e-08 
1.0 -1.46 0 5.0 5.5e-08 
1.0 -1.44 0 5.0 5.5e-08 
1.0 -1.42 0 5.0 5.5e-08 
1.0 -1.4 0 5.0 5.5e-08 
1.0 -1.38 0 5.0 5.5e-08 
1.0 -1.36 0 5.0 5.5e-08 
1.0 -1.34 0 5.0 5.5e-08 
1.0 -1.32 0 5.0 5.5e-08 
1.0 -1.3 0 5.0 5.5e-08 
1.0 -1.28 0 5.0 5.5e-08 
1.0 -1.26 0 5.0 5.5e-08 
1.0 -1.24 0 5.0 5.5e-08 
1.0 -1.22 0 5.0 5.5e-08 
1.0 -1.2 0 5.0 5.5e-08 
1.0 -1.18 0 5.0 5.5e-08 
1.0 -1.16 0 5.0 5.5e-08 
1.0 -1.14 0 5.0 5.5e-08 
1.0 -1.12 0 5.0 5.5e-08 
1.0 -1.1 0 5.0 5.5e-08 
1.0 -1.08 0 5.0 5.5e-08 
1.0 -1.06 0 5.0 5.5e-08 
1.0 -1.04 0 5.0 5.5e-08 
1.0 -1.02 0 5.0 5.5e-08 
1.0 -1.0 0 5.0 5.5e-08 
1.0 -0.98 0 5.0 5.5e-08 
1.0 -0.96 0 5.0 5.5e-08 
1.0 -0.94 0 5.0 5.5e-08 
1.0 -0.92 0 5.0 5.5e-08 
1.0 -0.9 0 5.0 5.5e-08 
1.0 -0.88 0 5.0 5.5e-08 
1.0 -0.86 0 5.0 5.5e-08 
1.0 -0.84 0 5.0 5.5e-08 
1.0 -0.82 0 5.0 5.5e-08 
1.0 -0.8 0 5.0 5.5e-08 
1.0 -0.78 0 5.0 5.5e-08 
1.0 -0.76 0 5.0 5.5e-08 
1.0 -0.74 0 5.0 5.5e-08 
1.0 -0.72 0 5.0 5.5e-08 
1.0 -0.7 0 5.0 5.5e-08 
1.0 -0.68 0 5.0 5.5e-08 
1.0 -0.66 0 5.0 5.5e-08 
1.0 -0.64 0 5.0 5.5e-08 
1.0 -0.62 0 5.0 5.5e-08 
1.0 -0.6 0 5.0 5.5e-08 
1.0 -0.58 0 5.0 5.5e-08 
1.0 -0.56 0 5.0 5.5e-08 
1.0 -0.54 0 5.0 5.5e-08 
1.0 -0.52 0 5.0 5.5e-08 
1.0 -0.5 0 5.0 5.5e-08 
1.0 -0.48 0 5.0 5.5e-08 
1.0 -0.46 0 5.0 5.5e-08 
1.0 -0.44 0 5.0 5.5e-08 
1.0 -0.42 0 5.0 5.5e-08 
1.0 -0.4 0 5.0 5.5e-08 
1.0 -0.38 0 5.0 5.5e-08 
1.0 -0.36 0 5.0 5.5e-08 
1.0 -0.34 0 5.0 5.5e-08 
1.0 -0.32 0 5.0 5.5e-08 
1.0 -0.3 0 5.0 5.5e-08 
1.0 -0.28 0 5.0 5.5e-08 
1.0 -0.26 0 5.0 5.5e-08 
1.0 -0.24 0 5.0 5.5e-08 
1.0 -0.22 0 5.0 5.5e-08 
1.0 -0.2 0 5.0 5.5e-08 
1.0 -0.18 0 5.0 5.5e-08 
1.0 -0.16 0 5.0 5.5e-08 
1.0 -0.14 0 5.0 5.5e-08 
1.0 -0.12 0 5.0 5.5e-08 
1.0 -0.1 0 5.0 5.5e-08 
1.0 -0.08 0 5.0 5.5e-08 
1.0 -0.06 0 5.0 5.5e-08 
1.0 -0.04 0 5.0 5.5e-08 
1.0 -0.02 0 5.0 5.5e-08 
1.0 1.33226762955e-15 0 5.0 5.5e-08 
1.0 0.02 0 5.0 5.5e-08 
1.0 0.04 0 5.0 5.5e-08 
1.0 0.06 0 5.0 5.5e-08 
1.0 0.08 0 5.0 5.5e-08 
1.0 0.1 0 5.0 5.5e-08 
1.0 0.12 0 5.0 5.5e-08 
1.0 0.14 0 5.0 5.5e-08 
1.0 0.16 0 5.0 5.5e-08 
1.0 0.18 0 5.0 5.5e-08 
1.0 0.2 0 5.0 5.5e-08 
1.0 0.22 0 5.0 5.5e-08 
1.0 0.24 0 5.0 5.5e-08 
1.0 0.26 0 5.0 5.5e-08 
1.0 0.28 0 5.0 5.5e-08 
1.0 0.3 0 5.0 5.5e-08 
1.0 0.32 0 5.0 5.5e-08 
1.0 0.34 0 5.0 5.5e-08 
1.0 0.36 0 5.0 5.5e-08 
1.0 0.38 0 5.0 5.5e-08 
1.0 0.4 0 5.0 5.5e-08 
1.0 0.42 0 5.0 5.5e-08 
1.0 0.44 0 5.0 5.5e-08 
1.0 0.46 0 5.0 5.5e-08 
1.0 0.48 0 5.0 5.5e-08 
1.0 0.5 0 5.0 5.5e-08 
1.0 0.52 0 5.0 5.5e-08 
1.0 0.54 0 5.0 5.5e-08 
1.0 0.56 0 5.0 5.5e-08 
1.0 0.58 0 5.0 5.5e-08 
1.0 0.6 0 5.0 5.5e-08 
1.0 0.62 0 5.0 5.5e-08 
1.0 0.64 0 5.0 5.5e-08 
1.0 0.66 0 5.0 5.5e-08 
1.0 0.68 0 5.0 5.5e-08 
1.0 0.7 0 5.0 5.5e-08 
1.0 0.72 0 5.0 5.5e-08 
1.0 0.74 0 5.0 5.5e-08 
1.0 0.76 0 5.0 5.5e-08 
1.0 0.78 0 5.0 5.5e-08 
1.0 0.8 0 5.0 5.5e-08 
1.0 0.82 0 5.0 5.5e-08 
1.0 0.84 0 5.0 5.5e-08 
1.0 0.86 0 5.0 5.5e-08 
1.0 0.88 0 5.0 5.5e-08 
1.0 0.9 0 5.0 5.5e-08 
1.0 0.92 0 5.0 5.5e-08 
1.0 0.94 0 5.0 5.5e-08 
1.0 0.96 0 5.0 5.5e-08 
1.0 0.98 0 5.0 5.5e-08 
1.0 1.0 0 5.0 5.5e-08 
1.0 1.02 0 5.0 5.5e-08 
1.0 1.04 0 5.0 5.5e-08 
1.0 1.06 0 5.0 5.5e-08 
1.0 1.08 0 5.0 5.5e-08 
1.0 1.1 0 5.0 5.5e-08 
1.0 1.12 0 5.0 5.5e-08 
1.0 1.14 0 5.0 5.5e-08 
1.0 1.16 0 5.0 5.5e-08 
1.0 1.18 0 5.0 5.5e-08 
1.0 1.2 0 5.0 5.5e-08 
1.0 1.22 0 5.0 5.5e-08 
1.0 1.24 0 5.0 5.5e-08 
1.0 1.26 0 5.0 5.5e-08 
1.0 1.28 0 5.0 5.5e-08 
1.0 1.3 0 5.0 5.5e-08 
1.0 1.32 0 5.0 5.5e-08 
1.0 1.34 0 5.0 5.5e-08 
1.0 1.36 0 5.0 5.5e-08 
1.0 1.38 0 5.0 5.5e-08 
1.0 1.4 0 5.0 5.5e-08 
1.0 1.42 0 5.0 5.5e-08 
1.0 1.44 0 5.0 5.5e-08 
1.0 1.46 0 5.0 5.5e-08 
1.0 1.48 0 5.0 5.5e-08 
1.0 -1.5 0 4.5 5.5e-08 
1.0 -1.48 0 4.5 5.5e-08 
1.0 -1.46 0 4.5 5.5e-08 
1.0 -1.44 0 4.5 5.5e-08 
1.0 -1.42 0 4.5 5.5e-08 
1.0 -1.4 0 4.5 5.5e-08 
1.0 -1.38 0 4.5 5.5e-08 
1.0 -1.36 0 4.5 5.5e-08 
1.0 -1.34 0 4.5 5.5e-08 
1.0 -1.32 0 4.5 5.5e-08 
1.0 -1.3 0 4.5 5.5e-08 
1.0 -1.28 0 4.5 5.5e-08 
1.0 -1.26 0 4.5 5.5e-08 
1.0 -1.24 0 4.5 5.5e-08 
1.0 -1.22 0 4.5 5.5e-08 
1.0 -1.2 0 4.5 5.5e-08 
1.0 -1.18 0 4.5 5.5e-08 
1.0 -1.16 0 4.5 5.5e-08 
1.0 -1.14 0 4.5 5.5e-08 
1.0 -1.12 0 4.5 5.5e-08 
1.0 -1.1 0 4.5 5.5e-08 
1.0 -1.08 0 4.5 5.5e-08 
1.0 -1.06 0 4.5 5.5e-08 
1.0 -1.04 0 4.5 5.5e-08 
1.0 -1.02 0 4.5 5.5e-08 
1.0 -1.0 0 4.5 5.5e-08 
1.0 -0.98 0 4.5 5.5e-08 
1.0 -0.96 0 4.5 5.5e-08 
1.0 -0.94 0 4.5 5.5e-08 
1.0 -0.92 0 4.5 5.5e-08 
1.0 -0.9 0 4.5 5.5e-08 
1.0 -0.88 0 4.5 5.5e-08 
1.0 -0.86 0 4.5 5.5e-08 
1.0 -0.84 0 4.5 5.5e-08 
1.0 -0.82 0 4.5 5.5e-08 
1.0 -0.8 0 4.5 5.5e-08 
1.0 -0.78 0 4.5 5.5e-08 
1.0 -0.76 0 4.5 5.5e-08 
1.0 -0.74 0 4.5 5.5e-08 
1.0 -0.72 0 4.5 5.5e-08 
1.0 -0.7 0 4.5 5.5e-08 
1.0 -0.68 0 4.5 5.5e-08 
1.0 -0.66 0 4.5 5.5e-08 
1.0 -0.64 0 4.5 5.5e-08 
1.0 -0.62 0 4.5 5.5e-08 
1.0 -0.6 0 4.5 5.5e-08 
1.0 -0.58 0 4.5 5.5e-08 
1.0 -0.56 0 4.5 5.5e-08 
1.0 -0.54 0 4.5 5.5e-08 
1.0 -0.52 0 4.5 5.5e-08 
1.0 -0.5 0 4.5 5.5e-08 
1.0 -0.48 0 4.5 5.5e-08 
1.0 -0.46 0 4.5 5.5e-08 
1.0 -0.44 0 4.5 5.5e-08 
1.0 -0.42 0 4.5 5.5e-08 
1.0 -0.4 0 4.5 5.5e-08 
1.0 -0.38 0 4.5 5.5e-08 
1.0 -0.36 0 4.5 5.5e-08 
1.0 -0.34 0 4.5 5.5e-08 
1.0 -0.32 0 4.5 5.5e-08 
1.0 -0.3 0 4.5 5.5e-08 
1.0 -0.28 0 4.5 5.5e-08 
1.0 -0.26 0 4.5 5.5e-08 
1.0 -0.24 0 4.5 5.5e-08 
1.0 -0.22 0 4.5 5.5e-08 
1.0 -0.2 0 4.5 5.5e-08 
1.0 -0.18 0 4.5 5.5e-08 
1.0 -0.16 0 4.5 5.5e-08 
1.0 -0.14 0 4.5 5.5e-08 
1.0 -0.12 0 4.5 5.5e-08 
1.0 -0.1 0 4.5 5.5e-08 
1.0 -0.08 0 4.5 5.5e-08 
1.0 -0.06 0 4.5 5.5e-08 
1.0 -0.04 0 4.5 5.5e-08 
1.0 -0.02 0 4.5 5.5e-08 
1.0 1.33226762955e-15 0 4.5 5.5e-08 
1.0 0.02 0 4.5 5.5e-08 
1.0 0.04 0 4.5 5.5e-08 
1.0 0.06 0 4.5 5.5e-08 
1.0 0.08 0 4.5 5.5e-08 
1.0 0.1 0 4.5 5.5e-08 
1.0 0.12 0 4.5 5.5e-08 
1.0 0.14 0 4.5 5.5e-08 
1.0 0.16 0 4.5 5.5e-08 
1.0 0.18 0 4.5 5.5e-08 
1.0 0.2 0 4.5 5.5e-08 
1.0 0.22 0 4.5 5.5e-08 
1.0 0.24 0 4.5 5.5e-08 
1.0 0.26 0 4.5 5.5e-08 
1.0 0.28 0 4.5 5.5e-08 
1.0 0.3 0 4.5 5.5e-08 
1.0 0.32 0 4.5 5.5e-08 
1.0 0.34 0 4.5 5.5e-08 
1.0 0.36 0 4.5 5.5e-08 
1.0 0.38 0 4.5 5.5e-08 
1.0 0.4 0 4.5 5.5e-08 
1.0 0.42 0 4.5 5.5e-08 
1.0 0.44 0 4.5 5.5e-08 
1.0 0.46 0 4.5 5.5e-08 
1.0 0.48 0 4.5 5.5e-08 
1.0 0.5 0 4.5 5.5e-08 
1.0 0.52 0 4.5 5.5e-08 
1.0 0.54 0 4.5 5.5e-08 
1.0 0.56 0 4.5 5.5e-08 
1.0 0.58 0 4.5 5.5e-08 
1.0 0.6 0 4.5 5.5e-08 
1.0 0.62 0 4.5 5.5e-08 
1.0 0.64 0 4.5 5.5e-08 
1.0 0.66 0 4.5 5.5e-08 
1.0 0.68 0 4.5 5.5e-08 
1.0 0.7 0 4.5 5.5e-08 
1.0 0.72 0 4.5 5.5e-08 
1.0 0.74 0 4.5 5.5e-08 
1.0 0.76 0 4.5 5.5e-08 
1.0 0.78 0 4.5 5.5e-08 
1.0 0.8 0 4.5 5.5e-08 
1.0 0.82 0 4.5 5.5e-08 
1.0 0.84 0 4.5 5.5e-08 
1.0 0.86 0 4.5 5.5e-08 
1.0 0.88 0 4.5 5.5e-08 
1.0 0.9 0 4.5 5.5e-08 
1.0 0.92 0 4.5 5.5e-08 
1.0 0.94 0 4.5 5.5e-08 
1.0 0.96 0 4.5 5.5e-08 
1.0 0.98 0 4.5 5.5e-08 
1.0 1.0 0 4.5 5.5e-08 
1.0 1.02 0 4.5 5.5e-08 
1.0 1.04 0 4.5 5.5e-08 
1.0 1.06 0 4.5 5.5e-08 
1.0 1.08 0 4.5 5.5e-08 
1.0 1.1 0 4.5 5.5e-08 
1.0 1.12 0 4.5 5.5e-08 
1.0 1.14 0 4.5 5.5e-08 
1.0 1.16 0 4.5 5.5e-08 
1.0 1.18 0 4.5 5.5e-08 
1.0 1.2 0 4.5 5.5e-08 
1.0 1.22 0 4.5 5.5e-08 
1.0 1.24 0 4.5 5.5e-08 
1.0 1.26 0 4.5 5.5e-08 
1.0 1.28 0 4.5 5.5e-08 
1.0 1.3 0 4.5 5.5e-08 
1.0 1.32 0 4.5 5.5e-08 
1.0 1.34 0 4.5 5.5e-08 
1.0 1.36 0 4.5 5.5e-08 
1.0 1.38 0 4.5 5.5e-08 
1.0 1.4 0 4.5 5.5e-08 
1.0 1.42 0 4.5 5.5e-08 
1.0 1.44 0 4.5 5.5e-08 
1.0 1.46 0 4.5 5.5e-08 
1.0 1.48 0 4.5 5.5e-08 
1.0 -1.5 0 4.0 5.5e-08 
1.0 -1.48 0 4.0 5.5e-08 
1.0 -1.46 0 4.0 5.5e-08 
1.0 -1.44 0 4.0 5.5e-08 
1.0 -1.42 0 4.0 5.5e-08 
1.0 -1.4 0 4.0 5.5e-08 
1.0 -1.38 0 4.0 5.5e-08 
1.0 -1.36 0 4.0 5.5e-08 
1.0 -1.34 0 4.0 5.5e-08 
1.0 -1.32 0 4.0 5.5e-08 
1.0 -1.3 0 4.0 5.5e-08 
1.0 -1.28 0 4.0 5.5e-08 
1.0 -1.26 0 4.0 5.5e-08 
1.0 -1.24 0 4.0 5.5e-08 
1.0 -1.22 0 4.0 5.5e-08 
1.0 -1.2 0 4.0 5.5e-08 
1.0 -1.18 0 4.0 5.5e-08 
1.0 -1.16 0 4.0 5.5e-08 
1.0 -1.14 0 4.0 5.5e-08 
1.0 -1.12 0 4.0 5.5e-08 
1.0 -1.1 0 4.0 5.5e-08 
1.0 -1.08 0 4.0 5.5e-08 
1.0 -1.06 0 4.0 5.5e-08 
1.0 -1.04 0 4.0 5.5e-08 
1.0 -1.02 0 4.0 5.5e-08 
1.0 -1.0 0 4.0 5.5e-08 
1.0 -0.98 0 4.0 5.5e-08 
1.0 -0.96 0 4.0 5.5e-08 
1.0 -0.94 0 4.0 5.5e-08 
1.0 -0.92 0 4.0 5.5e-08 
1.0 -0.9 0 4.0 5.5e-08 
1.0 -0.88 0 4.0 5.5e-08 
1.0 -0.86 0 4.0 5.5e-08 
1.0 -0.84 0 4.0 5.5e-08 
1.0 -0.82 0 4.0 5.5e-08 
1.0 -0.8 0 4.0 5.5e-08 
1.0 -0.78 0 4.0 5.5e-08 
1.0 -0.76 0 4.0 5.5e-08 
1.0 -0.74 0 4.0 5.5e-08 
1.0 -0.72 0 4.0 5.5e-08 
1.0 -0.7 0 4.0 5.5e-08 
1.0 -0.68 0 4.0 5.5e-08 
1.0 -0.66 0 4.0 5.5e-08 
1.0 -0.64 0 4.0 5.5e-08 
1.0 -0.62 0 4.0 5.5e-08 
1.0 -0.6 0 4.0 5.5e-08 
1.0 -0.58 0 4.0 5.5e-08 
1.0 -0.56 0 4.0 5.5e-08 
1.0 -0.54 0 4.0 5.5e-08 
1.0 -0.52 0 4.0 5.5e-08 
1.0 -0.5 0 4.0 5.5e-08 
1.0 -0.48 0 4.0 5.5e-08 
1.0 -0.46 0 4.0 5.5e-08 
1.0 -0.44 0 4.0 5.5e-08 
1.0 -0.42 0 4.0 5.5e-08 
1.0 -0.4 0 4.0 5.5e-08 
1.0 -0.38 0 4.0 5.5e-08 
1.0 -0.36 0 4.0 5.5e-08 
1.0 -0.34 0 4.0 5.5e-08 
1.0 -0.32 0 4.0 5.5e-08 
1.0 -0.3 0 4.0 5.5e-08 
1.0 -0.28 0 4.0 5.5e-08 
1.0 -0.26 0 4.0 5.5e-08 
1.0 -0.24 0 4.0 5.5e-08 
1.0 -0.22 0 4.0 5.5e-08 
1.0 -0.2 0 4.0 5.5e-08 
1.0 -0.18 0 4.0 5.5e-08 
1.0 -0.16 0 4.0 5.5e-08 
1.0 -0.14 0 4.0 5.5e-08 
1.0 -0.12 0 4.0 5.5e-08 
1.0 -0.1 0 4.0 5.5e-08 
1.0 -0.08 0 4.0 5.5e-08 
1.0 -0.06 0 4.0 5.5e-08 
1.0 -0.04 0 4.0 5.5e-08 
1.0 -0.02 0 4.0 5.5e-08 
1.0 1.33226762955e-15 0 4.0 5.5e-08 
1.0 0.02 0 4.0 5.5e-08 
1.0 0.04 0 4.0 5.5e-08 
1.0 0.06 0 4.0 5.5e-08 
1.0 0.08 0 4.0 5.5e-08 
1.0 0.1 0 4.0 5.5e-08 
1.0 0.12 0 4.0 5.5e-08 
1.0 0.14 0 4.0 5.5e-08 
1.0 0.16 0 4.0 5.5e-08 
1.0 0.18 0 4.0 5.5e-08 
1.0 0.2 0 4.0 5.5e-08 
1.0 0.22 0 4.0 5.5e-08 
1.0 0.24 0 4.0 5.5e-08 
1.0 0.26 0 4.0 5.5e-08 
1.0 0.28 0 4.0 5.5e-08 
1.0 0.3 0 4.0 5.5e-08 
1.0 0.32 0 4.0 5.5e-08 
1.0 0.34 0 4.0 5.5e-08 
1.0 0.36 0 4.0 5.5e-08 
1.0 0.38 0 4.0 5.5e-08 
1.0 0.4 0 4.0 5.5e-08 
1.0 0.42 0 4.0 5.5e-08 
1.0 0.44 0 4.0 5.5e-08 
1.0 0.46 0 4.0 5.5e-08 
1.0 0.48 0 4.0 5.5e-08 
1.0 0.5 0 4.0 5.5e-08 
1.0 0.52 0 4.0 5.5e-08 
1.0 0.54 0 4.0 5.5e-08 
1.0 0.56 0 4.0 5.5e-08 
1.0 0.58 0 4.0 5.5e-08 
1.0 0.6 0 4.0 5.5e-08 
1.0 0.62 0 4.0 5.5e-08 
1.0 0.64 0 4.0 5.5e-08 
1.0 0.66 0 4.0 5.5e-08 
1.0 0.68 0 4.0 5.5e-08 
1.0 0.7 0 4.0 5.5e-08 
1.0 0.72 0 4.0 5.5e-08 
1.0 0.74 0 4.0 5.5e-08 
1.0 0.76 0 4.0 5.5e-08 
1.0 0.78 0 4.0 5.5e-08 
1.0 0.8 0 4.0 5.5e-08 
1.0 0.82 0 4.0 5.5e-08 
1.0 0.84 0 4.0 5.5e-08 
1.0 0.86 0 4.0 5.5e-08 
1.0 0.88 0 4.0 5.5e-08 
1.0 0.9 0 4.0 5.5e-08 
1.0 0.92 0 4.0 5.5e-08 
1.0 0.94 0 4.0 5.5e-08 
1.0 0.96 0 4.0 5.5e-08 
1.0 0.98 0 4.0 5.5e-08 
1.0 1.0 0 4.0 5.5e-08 
1.0 1.02 0 4.0 5.5e-08 
1.0 1.04 0 4.0 5.5e-08 
1.0 1.06 0 4.0 5.5e-08 
1.0 1.08 0 4.0 5.5e-08 
1.0 1.1 0 4.0 5.5e-08 
1.0 1.12 0 4.0 5.5e-08 
1.0 1.14 0 4.0 5.5e-08 
1.0 1.16 0 4.0 5.5e-08 
1.0 1.18 0 4.0 5.5e-08 
1.0 1.2 0 4.0 5.5e-08 
1.0 1.22 0 4.0 5.5e-08 
1.0 1.24 0 4.0 5.5e-08 
1.0 1.26 0 4.0 5.5e-08 
1.0 1.28 0 4.0 5.5e-08 
1.0 1.3 0 4.0 5.5e-08 
1.0 1.32 0 4.0 5.5e-08 
1.0 1.34 0 4.0 5.5e-08 
1.0 1.36 0 4.0 5.5e-08 
1.0 1.38 0 4.0 5.5e-08 
1.0 1.4 0 4.0 5.5e-08 
1.0 1.42 0 4.0 5.5e-08 
1.0 1.44 0 4.0 5.5e-08 
1.0 1.46 0 4.0 5.5e-08 
1.0 1.48 0 4.0 5.5e-08 
1.0 -1.5 0 3.5 5.5e-08 
1.0 -1.48 0 3.5 5.5e-08 
1.0 -1.46 0 3.5 5.5e-08 
1.0 -1.44 0 3.5 5.5e-08 
1.0 -1.42 0 3.5 5.5e-08 
1.0 -1.4 0 3.5 5.5e-08 
1.0 -1.38 0 3.5 5.5e-08 
1.0 -1.36 0 3.5 5.5e-08 
1.0 -1.34 0 3.5 5.5e-08 
1.0 -1.32 0 3.5 5.5e-08 
1.0 -1.3 0 3.5 5.5e-08 
1.0 -1.28 0 3.5 5.5e-08 
1.0 -1.26 0 3.5 5.5e-08 
1.0 -1.24 0 3.5 5.5e-08 
1.0 -1.22 0 3.5 5.5e-08 
1.0 -1.2 0 3.5 5.5e-08 
1.0 -1.18 0 3.5 5.5e-08 
1.0 -1.16 0 3.5 5.5e-08 
1.0 -1.14 0 3.5 5.5e-08 
1.0 -1.12 0 3.5 5.5e-08 
1.0 -1.1 0 3.5 5.5e-08 
1.0 -1.08 0 3.5 5.5e-08 
1.0 -1.06 0 3.5 5.5e-08 
1.0 -1.04 0 3.5 5.5e-08 
1.0 -1.02 0 3.5 5.5e-08 
1.0 -1.0 0 3.5 5.5e-08 
1.0 -0.98 0 3.5 5.5e-08 
1.0 -0.96 0 3.5 5.5e-08 
1.0 -0.94 0 3.5 5.5e-08 
1.0 -0.92 0 3.5 5.5e-08 
1.0 -0.9 0 3.5 5.5e-08 
1.0 -0.88 0 3.5 5.5e-08 
1.0 -0.86 0 3.5 5.5e-08 
1.0 -0.84 0 3.5 5.5e-08 
1.0 -0.82 0 3.5 5.5e-08 
1.0 -0.8 0 3.5 5.5e-08 
1.0 -0.78 0 3.5 5.5e-08 
1.0 -0.76 0 3.5 5.5e-08 
1.0 -0.74 0 3.5 5.5e-08 
1.0 -0.72 0 3.5 5.5e-08 
1.0 -0.7 0 3.5 5.5e-08 
1.0 -0.68 0 3.5 5.5e-08 
1.0 -0.66 0 3.5 5.5e-08 
1.0 -0.64 0 3.5 5.5e-08 
1.0 -0.62 0 3.5 5.5e-08 
1.0 -0.6 0 3.5 5.5e-08 
1.0 -0.58 0 3.5 5.5e-08 
1.0 -0.56 0 3.5 5.5e-08 
1.0 -0.54 0 3.5 5.5e-08 
1.0 -0.52 0 3.5 5.5e-08 
1.0 -0.5 0 3.5 5.5e-08 
1.0 -0.48 0 3.5 5.5e-08 
1.0 -0.46 0 3.5 5.5e-08 
1.0 -0.44 0 3.5 5.5e-08 
1.0 -0.42 0 3.5 5.5e-08 
1.0 -0.4 0 3.5 5.5e-08 
1.0 -0.38 0 3.5 5.5e-08 
1.0 -0.36 0 3.5 5.5e-08 
1.0 -0.34 0 3.5 5.5e-08 
1.0 -0.32 0 3.5 5.5e-08 
1.0 -0.3 0 3.5 5.5e-08 
1.0 -0.28 0 3.5 5.5e-08 
1.0 -0.26 0 3.5 5.5e-08 
1.0 -0.24 0 3.5 5.5e-08 
1.0 -0.22 0 3.5 5.5e-08 
1.0 -0.2 0 3.5 5.5e-08 
1.0 -0.18 0 3.5 5.5e-08 
1.0 -0.16 0 3.5 5.5e-08 
1.0 -0.14 0 3.5 5.5e-08 
1.0 -0.12 0 3.5 5.5e-08 
1.0 -0.1 0 3.5 5.5e-08 
1.0 -0.08 0 3.5 5.5e-08 
1.0 -0.06 0 3.5 5.5e-08 
1.0 -0.04 0 3.5 5.5e-08 
1.0 -0.02 0 3.5 5.5e-08 
1.0 1.33226762955e-15 0 3.5 5.5e-08 
1.0 0.02 0 3.5 5.5e-08 
1.0 0.04 0 3.5 5.5e-08 
1.0 0.06 0 3.5 5.5e-08 
1.0 0.08 0 3.5 5.5e-08 
1.0 0.1 0 3.5 5.5e-08 
1.0 0.12 0 3.5 5.5e-08 
1.0 0.14 0 3.5 5.5e-08 
1.0 0.16 0 3.5 5.5e-08 
1.0 0.18 0 3.5 5.5e-08 
1.0 0.2 0 3.5 5.5e-08 
1.0 0.22 0 3.5 5.5e-08 
1.0 0.24 0 3.5 5.5e-08 
1.0 0.26 0 3.5 5.5e-08 
1.0 0.28 0 3.5 5.5e-08 
1.0 0.3 0 3.5 5.5e-08 
1.0 0.32 0 3.5 5.5e-08 
1.0 0.34 0 3.5 5.5e-08 
1.0 0.36 0 3.5 5.5e-08 
1.0 0.38 0 3.5 5.5e-08 
1.0 0.4 0 3.5 5.5e-08 
1.0 0.42 0 3.5 5.5e-08 
1.0 0.44 0 3.5 5.5e-08 
1.0 0.46 0 3.5 5.5e-08 
1.0 0.48 0 3.5 5.5e-08 
1.0 0.5 0 3.5 5.5e-08 
1.0 0.52 0 3.5 5.5e-08 
1.0 0.54 0 3.5 5.5e-08 
1.0 0.56 0 3.5 5.5e-08 
1.0 0.58 0 3.5 5.5e-08 
1.0 0.6 0 3.5 5.5e-08 
1.0 0.62 0 3.5 5.5e-08 
1.0 0.64 0 3.5 5.5e-08 
1.0 0.66 0 3.5 5.5e-08 
1.0 0.68 0 3.5 5.5e-08 
1.0 0.7 0 3.5 5.5e-08 
1.0 0.72 0 3.5 5.5e-08 
1.0 0.74 0 3.5 5.5e-08 
1.0 0.76 0 3.5 5.5e-08 
1.0 0.78 0 3.5 5.5e-08 
1.0 0.8 0 3.5 5.5e-08 
1.0 0.82 0 3.5 5.5e-08 
1.0 0.84 0 3.5 5.5e-08 
1.0 0.86 0 3.5 5.5e-08 
1.0 0.88 0 3.5 5.5e-08 
1.0 0.9 0 3.5 5.5e-08 
1.0 0.92 0 3.5 5.5e-08 
1.0 0.94 0 3.5 5.5e-08 
1.0 0.96 0 3.5 5.5e-08 
1.0 0.98 0 3.5 5.5e-08 
1.0 1.0 0 3.5 5.5e-08 
1.0 1.02 0 3.5 5.5e-08 
1.0 1.04 0 3.5 5.5e-08 
1.0 1.06 0 3.5 5.5e-08 
1.0 1.08 0 3.5 5.5e-08 
1.0 1.1 0 3.5 5.5e-08 
1.0 1.12 0 3.5 5.5e-08 
1.0 1.14 0 3.5 5.5e-08 
1.0 1.16 0 3.5 5.5e-08 
1.0 1.18 0 3.5 5.5e-08 
1.0 1.2 0 3.5 5.5e-08 
1.0 1.22 0 3.5 5.5e-08 
1.0 1.24 0 3.5 5.5e-08 
1.0 1.26 0 3.5 5.5e-08 
1.0 1.28 0 3.5 5.5e-08 
1.0 1.3 0 3.5 5.5e-08 
1.0 1.32 0 3.5 5.5e-08 
1.0 1.34 0 3.5 5.5e-08 
1.0 1.36 0 3.5 5.5e-08 
1.0 1.38 0 3.5 5.5e-08 
1.0 1.4 0 3.5 5.5e-08 
1.0 1.42 0 3.5 5.5e-08 
1.0 1.44 0 3.5 5.5e-08 
1.0 1.46 0 3.5 5.5e-08 
1.0 1.48 0 3.5 5.5e-08 
1.0 -1.5 0 3.0 5.5e-08 
1.0 -1.48 0 3.0 5.5e-08 
1.0 -1.46 0 3.0 5.5e-08 
1.0 -1.44 0 3.0 5.5e-08 
1.0 -1.42 0 3.0 5.5e-08 
1.0 -1.4 0 3.0 5.5e-08 
1.0 -1.38 0 3.0 5.5e-08 
1.0 -1.36 0 3.0 5.5e-08 
1.0 -1.34 0 3.0 5.5e-08 
1.0 -1.32 0 3.0 5.5e-08 
1.0 -1.3 0 3.0 5.5e-08 
1.0 -1.28 0 3.0 5.5e-08 
1.0 -1.26 0 3.0 5.5e-08 
1.0 -1.24 0 3.0 5.5e-08 
1.0 -1.22 0 3.0 5.5e-08 
1.0 -1.2 0 3.0 5.5e-08 
1.0 -1.18 0 3.0 5.5e-08 
1.0 -1.16 0 3.0 5.5e-08 
1.0 -1.14 0 3.0 5.5e-08 
1.0 -1.12 0 3.0 5.5e-08 
1.0 -1.1 0 3.0 5.5e-08 
1.0 -1.08 0 3.0 5.5e-08 
1.0 -1.06 0 3.0 5.5e-08 
1.0 -1.04 0 3.0 5.5e-08 
1.0 -1.02 0 3.0 5.5e-08 
1.0 -1.0 0 3.0 5.5e-08 
1.0 -0.98 0 3.0 5.5e-08 
1.0 -0.96 0 3.0 5.5e-08 
1.0 -0.94 0 3.0 5.5e-08 
1.0 -0.92 0 3.0 5.5e-08 
1.0 -0.9 0 3.0 5.5e-08 
1.0 -0.88 0 3.0 5.5e-08 
1.0 -0.86 0 3.0 5.5e-08 
1.0 -0.84 0 3.0 5.5e-08 
1.0 -0.82 0 3.0 5.5e-08 
1.0 -0.8 0 3.0 5.5e-08 
1.0 -0.78 0 3.0 5.5e-08 
1.0 -0.76 0 3.0 5.5e-08 
1.0 -0.74 0 3.0 5.5e-08 
1.0 -0.72 0 3.0 5.5e-08 
1.0 -0.7 0 3.0 5.5e-08 
1.0 -0.68 0 3.0 5.5e-08 
1.0 -0.66 0 3.0 5.5e-08 
1.0 -0.64 0 3.0 5.5e-08 
1.0 -0.62 0 3.0 5.5e-08 
1.0 -0.6 0 3.0 5.5e-08 
1.0 -0.58 0 3.0 5.5e-08 
1.0 -0.56 0 3.0 5.5e-08 
1.0 -0.54 0 3.0 5.5e-08 
1.0 -0.52 0 3.0 5.5e-08 
1.0 -0.5 0 3.0 5.5e-08 
1.0 -0.48 0 3.0 5.5e-08 
1.0 -0.46 0 3.0 5.5e-08 
1.0 -0.44 0 3.0 5.5e-08 
1.0 -0.42 0 3.0 5.5e-08 
1.0 -0.4 0 3.0 5.5e-08 
1.0 -0.38 0 3.0 5.5e-08 
1.0 -0.36 0 3.0 5.5e-08 
1.0 -0.34 0 3.0 5.5e-08 
1.0 -0.32 0 3.0 5.5e-08 
1.0 -0.3 0 3.0 5.5e-08 
1.0 -0.28 0 3.0 5.5e-08 
1.0 -0.26 0 3.0 5.5e-08 
1.0 -0.24 0 3.0 5.5e-08 
1.0 -0.22 0 3.0 5.5e-08 
1.0 -0.2 0 3.0 5.5e-08 
1.0 -0.18 0 3.0 5.5e-08 
1.0 -0.16 0 3.0 5.5e-08 
1.0 -0.14 0 3.0 5.5e-08 
1.0 -0.12 0 3.0 5.5e-08 
1.0 -0.1 0 3.0 5.5e-08 
1.0 -0.08 0 3.0 5.5e-08 
1.0 -0.06 0 3.0 5.5e-08 
1.0 -0.04 0 3.0 5.5e-08 
1.0 -0.02 0 3.0 5.5e-08 
1.0 1.33226762955e-15 0 3.0 5.5e-08 
1.0 0.02 0 3.0 5.5e-08 
1.0 0.04 0 3.0 5.5e-08 
1.0 0.06 0 3.0 5.5e-08 
1.0 0.08 0 3.0 5.5e-08 
1.0 0.1 0 3.0 5.5e-08 
1.0 0.12 0 3.0 5.5e-08 
1.0 0.14 0 3.0 5.5e-08 
1.0 0.16 0 3.0 5.5e-08 
1.0 0.18 0 3.0 5.5e-08 
1.0 0.2 0 3.0 5.5e-08 
1.0 0.22 0 3.0 5.5e-08 
1.0 0.24 0 3.0 5.5e-08 
1.0 0.26 0 3.0 5.5e-08 
1.0 0.28 0 3.0 5.5e-08 
1.0 0.3 0 3.0 5.5e-08 
1.0 0.32 0 3.0 5.5e-08 
1.0 0.34 0 3.0 5.5e-08 
1.0 0.36 0 3.0 5.5e-08 
1.0 0.38 0 3.0 5.5e-08 
1.0 0.4 0 3.0 5.5e-08 
1.0 0.42 0 3.0 5.5e-08 
1.0 0.44 0 3.0 5.5e-08 
1.0 0.46 0 3.0 5.5e-08 
1.0 0.48 0 3.0 5.5e-08 
1.0 0.5 0 3.0 5.5e-08 
1.0 0.52 0 3.0 5.5e-08 
1.0 0.54 0 3.0 5.5e-08 
1.0 0.56 0 3.0 5.5e-08 
1.0 0.58 0 3.0 5.5e-08 
1.0 0.6 0 3.0 5.5e-08 
1.0 0.62 0 3.0 5.5e-08 
1.0 0.64 0 3.0 5.5e-08 
1.0 0.66 0 3.0 5.5e-08 
1.0 0.68 0 3.0 5.5e-08 
1.0 0.7 0 3.0 5.5e-08 
1.0 0.72 0 3.0 5.5e-08 
1.0 0.74 0 3.0 5.5e-08 
1.0 0.76 0 3.0 5.5e-08 
1.0 0.78 0 3.0 5.5e-08 
1.0 0.8 0 3.0 5.5e-08 
1.0 0.82 0 3.0 5.5e-08 
1.0 0.84 0 3.0 5.5e-08 
1.0 0.86 0 3.0 5.5e-08 
1.0 0.88 0 3.0 5.5e-08 
1.0 0.9 0 3.0 5.5e-08 
1.0 0.92 0 3.0 5.5e-08 
1.0 0.94 0 3.0 5.5e-08 
1.0 0.96 0 3.0 5.5e-08 
1.0 0.98 0 3.0 5.5e-08 
1.0 1.0 0 3.0 5.5e-08 
1.0 1.02 0 3.0 5.5e-08 
1.0 1.04 0 3.0 5.5e-08 
1.0 1.06 0 3.0 5.5e-08 
1.0 1.08 0 3.0 5.5e-08 
1.0 1.1 0 3.0 5.5e-08 
1.0 1.12 0 3.0 5.5e-08 
1.0 1.14 0 3.0 5.5e-08 
1.0 1.16 0 3.0 5.5e-08 
1.0 1.18 0 3.0 5.5e-08 
1.0 1.2 0 3.0 5.5e-08 
1.0 1.22 0 3.0 5.5e-08 
1.0 1.24 0 3.0 5.5e-08 
1.0 1.26 0 3.0 5.5e-08 
1.0 1.28 0 3.0 5.5e-08 
1.0 1.3 0 3.0 5.5e-08 
1.0 1.32 0 3.0 5.5e-08 
1.0 1.34 0 3.0 5.5e-08 
1.0 1.36 0 3.0 5.5e-08 
1.0 1.38 0 3.0 5.5e-08 
1.0 1.4 0 3.0 5.5e-08 
1.0 1.42 0 3.0 5.5e-08 
1.0 1.44 0 3.0 5.5e-08 
1.0 1.46 0 3.0 5.5e-08 
1.0 1.48 0 3.0 5.5e-08 
1.0 -1.5 0 2.5 5.5e-08 
1.0 -1.48 0 2.5 5.5e-08 
1.0 -1.46 0 2.5 5.5e-08 
1.0 -1.44 0 2.5 5.5e-08 
1.0 -1.42 0 2.5 5.5e-08 
1.0 -1.4 0 2.5 5.5e-08 
1.0 -1.38 0 2.5 5.5e-08 
1.0 -1.36 0 2.5 5.5e-08 
1.0 -1.34 0 2.5 5.5e-08 
1.0 -1.32 0 2.5 5.5e-08 
1.0 -1.3 0 2.5 5.5e-08 
1.0 -1.28 0 2.5 5.5e-08 
1.0 -1.26 0 2.5 5.5e-08 
1.0 -1.24 0 2.5 5.5e-08 
1.0 -1.22 0 2.5 5.5e-08 
1.0 -1.2 0 2.5 5.5e-08 
1.0 -1.18 0 2.5 5.5e-08 
1.0 -1.16 0 2.5 5.5e-08 
1.0 -1.14 0 2.5 5.5e-08 
1.0 -1.12 0 2.5 5.5e-08 
1.0 -1.1 0 2.5 5.5e-08 
1.0 -1.08 0 2.5 5.5e-08 
1.0 -1.06 0 2.5 5.5e-08 
1.0 -1.04 0 2.5 5.5e-08 
1.0 -1.02 0 2.5 5.5e-08 
1.0 -1.0 0 2.5 5.5e-08 
1.0 -0.98 0 2.5 5.5e-08 
1.0 -0.96 0 2.5 5.5e-08 
1.0 -0.94 0 2.5 5.5e-08 
1.0 -0.92 0 2.5 5.5e-08 
1.0 -0.9 0 2.5 5.5e-08 
1.0 -0.88 0 2.5 5.5e-08 
1.0 -0.86 0 2.5 5.5e-08 
1.0 -0.84 0 2.5 5.5e-08 
1.0 -0.82 0 2.5 5.5e-08 
1.0 -0.8 0 2.5 5.5e-08 
1.0 -0.78 0 2.5 5.5e-08 
1.0 -0.76 0 2.5 5.5e-08 
1.0 -0.74 0 2.5 5.5e-08 
1.0 -0.72 0 2.5 5.5e-08 
1.0 -0.7 0 2.5 5.5e-08 
1.0 -0.68 0 2.5 5.5e-08 
1.0 -0.66 0 2.5 5.5e-08 
1.0 -0.64 0 2.5 5.5e-08 
1.0 -0.62 0 2.5 5.5e-08 
1.0 -0.6 0 2.5 5.5e-08 
1.0 -0.58 0 2.5 5.5e-08 
1.0 -0.56 0 2.5 5.5e-08 
1.0 -0.54 0 2.5 5.5e-08 
1.0 -0.52 0 2.5 5.5e-08 
1.0 -0.5 0 2.5 5.5e-08 
1.0 -0.48 0 2.5 5.5e-08 
1.0 -0.46 0 2.5 5.5e-08 
1.0 -0.44 0 2.5 5.5e-08 
1.0 -0.42 0 2.5 5.5e-08 
1.0 -0.4 0 2.5 5.5e-08 
1.0 -0.38 0 2.5 5.5e-08 
1.0 -0.36 0 2.5 5.5e-08 
1.0 -0.34 0 2.5 5.5e-08 
1.0 -0.32 0 2.5 5.5e-08 
1.0 -0.3 0 2.5 5.5e-08 
1.0 -0.28 0 2.5 5.5e-08 
1.0 -0.26 0 2.5 5.5e-08 
1.0 -0.24 0 2.5 5.5e-08 
1.0 -0.22 0 2.5 5.5e-08 
1.0 -0.2 0 2.5 5.5e-08 
1.0 -0.18 0 2.5 5.5e-08 
1.0 -0.16 0 2.5 5.5e-08 
1.0 -0.14 0 2.5 5.5e-08 
1.0 -0.12 0 2.5 5.5e-08 
1.0 -0.1 0 2.5 5.5e-08 
1.0 -0.08 0 2.5 5.5e-08 
1.0 -0.06 0 2.5 5.5e-08 
1.0 -0.04 0 2.5 5.5e-08 
1.0 -0.02 0 2.5 5.5e-08 
1.0 1.33226762955e-15 0 2.5 5.5e-08 
1.0 0.02 0 2.5 5.5e-08 
1.0 0.04 0 2.5 5.5e-08 
1.0 0.06 0 2.5 5.5e-08 
1.0 0.08 0 2.5 5.5e-08 
1.0 0.1 0 2.5 5.5e-08 
1.0 0.12 0 2.5 5.5e-08 
1.0 0.14 0 2.5 5.5e-08 
1.0 0.16 0 2.5 5.5e-08 
1.0 0.18 0 2.5 5.5e-08 
1.0 0.2 0 2.5 5.5e-08 
1.0 0.22 0 2.5 5.5e-08 
1.0 0.24 0 2.5 5.5e-08 
1.0 0.26 0 2.5 5.5e-08 
1.0 0.28 0 2.5 5.5e-08 
1.0 0.3 0 2.5 5.5e-08 
1.0 0.32 0 2.5 5.5e-08 
1.0 0.34 0 2.5 5.5e-08 
1.0 0.36 0 2.5 5.5e-08 
1.0 0.38 0 2.5 5.5e-08 
1.0 0.4 0 2.5 5.5e-08 
1.0 0.42 0 2.5 5.5e-08 
1.0 0.44 0 2.5 5.5e-08 
1.0 0.46 0 2.5 5.5e-08 
1.0 0.48 0 2.5 5.5e-08 
1.0 0.5 0 2.5 5.5e-08 
1.0 0.52 0 2.5 5.5e-08 
1.0 0.54 0 2.5 5.5e-08 
1.0 0.56 0 2.5 5.5e-08 
1.0 0.58 0 2.5 5.5e-08 
1.0 0.6 0 2.5 5.5e-08 
1.0 0.62 0 2.5 5.5e-08 
1.0 0.64 0 2.5 5.5e-08 
1.0 0.66 0 2.5 5.5e-08 
1.0 0.68 0 2.5 5.5e-08 
1.0 0.7 0 2.5 5.5e-08 
1.0 0.72 0 2.5 5.5e-08 
1.0 0.74 0 2.5 5.5e-08 
1.0 0.76 0 2.5 5.5e-08 
1.0 0.78 0 2.5 5.5e-08 
1.0 0.8 0 2.5 5.5e-08 
1.0 0.82 0 2.5 5.5e-08 
1.0 0.84 0 2.5 5.5e-08 
1.0 0.86 0 2.5 5.5e-08 
1.0 0.88 0 2.5 5.5e-08 
1.0 0.9 0 2.5 5.5e-08 
1.0 0.92 0 2.5 5.5e-08 
1.0 0.94 0 2.5 5.5e-08 
1.0 0.96 0 2.5 5.5e-08 
1.0 0.98 0 2.5 5.5e-08 
1.0 1.0 0 2.5 5.5e-08 
1.0 1.02 0 2.5 5.5e-08 
1.0 1.04 0 2.5 5.5e-08 
1.0 1.06 0 2.5 5.5e-08 
1.0 1.08 0 2.5 5.5e-08 
1.0 1.1 0 2.5 5.5e-08 
1.0 1.12 0 2.5 5.5e-08 
1.0 1.14 0 2.5 5.5e-08 
1.0 1.16 0 2.5 5.5e-08 
1.0 1.18 0 2.5 5.5e-08 
1.0 1.2 0 2.5 5.5e-08 
1.0 1.22 0 2.5 5.5e-08 
1.0 1.24 0 2.5 5.5e-08 
1.0 1.26 0 2.5 5.5e-08 
1.0 1.28 0 2.5 5.5e-08 
1.0 1.3 0 2.5 5.5e-08 
1.0 1.32 0 2.5 5.5e-08 
1.0 1.34 0 2.5 5.5e-08 
1.0 1.36 0 2.5 5.5e-08 
1.0 1.38 0 2.5 5.5e-08 
1.0 1.4 0 2.5 5.5e-08 
1.0 1.42 0 2.5 5.5e-08 
1.0 1.44 0 2.5 5.5e-08 
1.0 1.46 0 2.5 5.5e-08 
1.0 1.48 0 2.5 5.5e-08 
1.0 -1.5 0 2.0 5.5e-08 
1.0 -1.48 0 2.0 5.5e-08 
1.0 -1.46 0 2.0 5.5e-08 
1.0 -1.44 0 2.0 5.5e-08 
1.0 -1.42 0 2.0 5.5e-08 
1.0 -1.4 0 2.0 5.5e-08 
1.0 -1.38 0 2.0 5.5e-08 
1.0 -1.36 0 2.0 5.5e-08 
1.0 -1.34 0 2.0 5.5e-08 
1.0 -1.32 0 2.0 5.5e-08 
1.0 -1.3 0 2.0 5.5e-08 
1.0 -1.28 0 2.0 5.5e-08 
1.0 -1.26 0 2.0 5.5e-08 
1.0 -1.24 0 2.0 5.5e-08 
1.0 -1.22 0 2.0 5.5e-08 
1.0 -1.2 0 2.0 5.5e-08 
1.0 -1.18 0 2.0 5.5e-08 
1.0 -1.16 0 2.0 5.5e-08 
1.0 -1.14 0 2.0 5.5e-08 
1.0 -1.12 0 2.0 5.5e-08 
1.0 -1.1 0 2.0 5.5e-08 
1.0 -1.08 0 2.0 5.5e-08 
1.0 -1.06 0 2.0 5.5e-08 
1.0 -1.04 0 2.0 5.5e-08 
1.0 -1.02 0 2.0 5.5e-08 
1.0 -1.0 0 2.0 5.5e-08 
1.0 -0.98 0 2.0 5.5e-08 
1.0 -0.96 0 2.0 5.5e-08 
1.0 -0.94 0 2.0 5.5e-08 
1.0 -0.92 0 2.0 5.5e-08 
1.0 -0.9 0 2.0 5.5e-08 
1.0 -0.88 0 2.0 5.5e-08 
1.0 -0.86 0 2.0 5.5e-08 
1.0 -0.84 0 2.0 5.5e-08 
1.0 -0.82 0 2.0 5.5e-08 
1.0 -0.8 0 2.0 5.5e-08 
1.0 -0.78 0 2.0 5.5e-08 
1.0 -0.76 0 2.0 5.5e-08 
1.0 -0.74 0 2.0 5.5e-08 
1.0 -0.72 0 2.0 5.5e-08 
1.0 -0.7 0 2.0 5.5e-08 
1.0 -0.68 0 2.0 5.5e-08 
1.0 -0.66 0 2.0 5.5e-08 
1.0 -0.64 0 2.0 5.5e-08 
1.0 -0.62 0 2.0 5.5e-08 
1.0 -0.6 0 2.0 5.5e-08 
1.0 -0.58 0 2.0 5.5e-08 
1.0 -0.56 0 2.0 5.5e-08 
1.0 -0.54 0 2.0 5.5e-08 
1.0 -0.52 0 2.0 5.5e-08 
1.0 -0.5 0 2.0 5.5e-08 
1.0 -0.48 0 2.0 5.5e-08 
1.0 -0.46 0 2.0 5.5e-08 
1.0 -0.44 0 2.0 5.5e-08 
1.0 -0.42 0 2.0 5.5e-08 
1.0 -0.4 0 2.0 5.5e-08 
1.0 -0.38 0 2.0 5.5e-08 
1.0 -0.36 0 2.0 5.5e-08 
1.0 -0.34 0 2.0 5.5e-08 
1.0 -0.32 0 2.0 5.5e-08 
1.0 -0.3 0 2.0 5.5e-08 
1.0 -0.28 0 2.0 5.5e-08 
1.0 -0.26 0 2.0 5.5e-08 
1.0 -0.24 0 2.0 5.5e-08 
1.0 -0.22 0 2.0 5.5e-08 
1.0 -0.2 0 2.0 5.5e-08 
1.0 -0.18 0 2.0 5.5e-08 
1.0 -0.16 0 2.0 5.5e-08 
1.0 -0.14 0 2.0 5.5e-08 
1.0 -0.12 0 2.0 5.5e-08 
1.0 -0.1 0 2.0 5.5e-08 
1.0 -0.08 0 2.0 5.5e-08 
1.0 -0.06 0 2.0 5.5e-08 
1.0 -0.04 0 2.0 5.5e-08 
1.0 -0.02 0 2.0 5.5e-08 
1.0 1.33226762955e-15 0 2.0 5.5e-08 
1.0 0.02 0 2.0 5.5e-08 
1.0 0.04 0 2.0 5.5e-08 
1.0 0.06 0 2.0 5.5e-08 
1.0 0.08 0 2.0 5.5e-08 
1.0 0.1 0 2.0 5.5e-08 
1.0 0.12 0 2.0 5.5e-08 
1.0 0.14 0 2.0 5.5e-08 
1.0 0.16 0 2.0 5.5e-08 
1.0 0.18 0 2.0 5.5e-08 
1.0 0.2 0 2.0 5.5e-08 
1.0 0.22 0 2.0 5.5e-08 
1.0 0.24 0 2.0 5.5e-08 
1.0 0.26 0 2.0 5.5e-08 
1.0 0.28 0 2.0 5.5e-08 
1.0 0.3 0 2.0 5.5e-08 
1.0 0.32 0 2.0 5.5e-08 
1.0 0.34 0 2.0 5.5e-08 
1.0 0.36 0 2.0 5.5e-08 
1.0 0.38 0 2.0 5.5e-08 
1.0 0.4 0 2.0 5.5e-08 
1.0 0.42 0 2.0 5.5e-08 
1.0 0.44 0 2.0 5.5e-08 
1.0 0.46 0 2.0 5.5e-08 
1.0 0.48 0 2.0 5.5e-08 
1.0 0.5 0 2.0 5.5e-08 
1.0 0.52 0 2.0 5.5e-08 
1.0 0.54 0 2.0 5.5e-08 
1.0 0.56 0 2.0 5.5e-08 
1.0 0.58 0 2.0 5.5e-08 
1.0 0.6 0 2.0 5.5e-08 
1.0 0.62 0 2.0 5.5e-08 
1.0 0.64 0 2.0 5.5e-08 
1.0 0.66 0 2.0 5.5e-08 
1.0 0.68 0 2.0 5.5e-08 
1.0 0.7 0 2.0 5.5e-08 
1.0 0.72 0 2.0 5.5e-08 
1.0 0.74 0 2.0 5.5e-08 
1.0 0.76 0 2.0 5.5e-08 
1.0 0.78 0 2.0 5.5e-08 
1.0 0.8 0 2.0 5.5e-08 
1.0 0.82 0 2.0 5.5e-08 
1.0 0.84 0 2.0 5.5e-08 
1.0 0.86 0 2.0 5.5e-08 
1.0 0.88 0 2.0 5.5e-08 
1.0 0.9 0 2.0 5.5e-08 
1.0 0.92 0 2.0 5.5e-08 
1.0 0.94 0 2.0 5.5e-08 
1.0 0.96 0 2.0 5.5e-08 
1.0 0.98 0 2.0 5.5e-08 
1.0 1.0 0 2.0 5.5e-08 
1.0 1.02 0 2.0 5.5e-08 
1.0 1.04 0 2.0 5.5e-08 
1.0 1.06 0 2.0 5.5e-08 
1.0 1.08 0 2.0 5.5e-08 
1.0 1.1 0 2.0 5.5e-08 
1.0 1.12 0 2.0 5.5e-08 
1.0 1.14 0 2.0 5.5e-08 
1.0 1.16 0 2.0 5.5e-08 
1.0 1.18 0 2.0 5.5e-08 
1.0 1.2 0 2.0 5.5e-08 
1.0 1.22 0 2.0 5.5e-08 
1.0 1.24 0 2.0 5.5e-08 
1.0 1.26 0 2.0 5.5e-08 
1.0 1.28 0 2.0 5.5e-08 
1.0 1.3 0 2.0 5.5e-08 
1.0 1.32 0 2.0 5.5e-08 
1.0 1.34 0 2.0 5.5e-08 
1.0 1.36 0 2.0 5.5e-08 
1.0 1.38 0 2.0 5.5e-08 
1.0 1.4 0 2.0 5.5e-08 
1.0 1.42 0 2.0 5.5e-08 
1.0 1.44 0 2.0 5.5e-08 
1.0 1.46 0 2.0 5.5e-08 
1.0 1.48 0 2.0 5.5e-08 
1.0 -1.5 0 1.5 5.5e-08 
1.0 -1.48 0 1.5 5.5e-08 
1.0 -1.46 0 1.5 5.5e-08 
1.0 -1.44 0 1.5 5.5e-08 
1.0 -1.42 0 1.5 5.5e-08 
1.0 -1.4 0 1.5 5.5e-08 
1.0 -1.38 0 1.5 5.5e-08 
1.0 -1.36 0 1.5 5.5e-08 
1.0 -1.34 0 1.5 5.5e-08 
1.0 -1.32 0 1.5 5.5e-08 
1.0 -1.3 0 1.5 5.5e-08 
1.0 -1.28 0 1.5 5.5e-08 
1.0 -1.26 0 1.5 5.5e-08 
1.0 -1.24 0 1.5 5.5e-08 
1.0 -1.22 0 1.5 5.5e-08 
1.0 -1.2 0 1.5 5.5e-08 
1.0 -1.18 0 1.5 5.5e-08 
1.0 -1.16 0 1.5 5.5e-08 
1.0 -1.14 0 1.5 5.5e-08 
1.0 -1.12 0 1.5 5.5e-08 
1.0 -1.1 0 1.5 5.5e-08 
1.0 -1.08 0 1.5 5.5e-08 
1.0 -1.06 0 1.5 5.5e-08 
1.0 -1.04 0 1.5 5.5e-08 
1.0 -1.02 0 1.5 5.5e-08 
1.0 -1.0 0 1.5 5.5e-08 
1.0 -0.98 0 1.5 5.5e-08 
1.0 -0.96 0 1.5 5.5e-08 
1.0 -0.94 0 1.5 5.5e-08 
1.0 -0.92 0 1.5 5.5e-08 
1.0 -0.9 0 1.5 5.5e-08 
1.0 -0.88 0 1.5 5.5e-08 
1.0 -0.86 0 1.5 5.5e-08 
1.0 -0.84 0 1.5 5.5e-08 
1.0 -0.82 0 1.5 5.5e-08 
1.0 -0.8 0 1.5 5.5e-08 
1.0 -0.78 0 1.5 5.5e-08 
1.0 -0.76 0 1.5 5.5e-08 
1.0 -0.74 0 1.5 5.5e-08 
1.0 -0.72 0 1.5 5.5e-08 
1.0 -0.7 0 1.5 5.5e-08 
1.0 -0.68 0 1.5 5.5e-08 
1.0 -0.66 0 1.5 5.5e-08 
1.0 -0.64 0 1.5 5.5e-08 
1.0 -0.62 0 1.5 5.5e-08 
1.0 -0.6 0 1.5 5.5e-08 
1.0 -0.58 0 1.5 5.5e-08 
1.0 -0.56 0 1.5 5.5e-08 
1.0 -0.54 0 1.5 5.5e-08 
1.0 -0.52 0 1.5 5.5e-08 
1.0 -0.5 0 1.5 5.5e-08 
1.0 -0.48 0 1.5 5.5e-08 
1.0 -0.46 0 1.5 5.5e-08 
1.0 -0.44 0 1.5 5.5e-08 
1.0 -0.42 0 1.5 5.5e-08 
1.0 -0.4 0 1.5 5.5e-08 
1.0 -0.38 0 1.5 5.5e-08 
1.0 -0.36 0 1.5 5.5e-08 
1.0 -0.34 0 1.5 5.5e-08 
1.0 -0.32 0 1.5 5.5e-08 
1.0 -0.3 0 1.5 5.5e-08 
1.0 -0.28 0 1.5 5.5e-08 
1.0 -0.26 0 1.5 5.5e-08 
1.0 -0.24 0 1.5 5.5e-08 
1.0 -0.22 0 1.5 5.5e-08 
1.0 -0.2 0 1.5 5.5e-08 
1.0 -0.18 0 1.5 5.5e-08 
1.0 -0.16 0 1.5 5.5e-08 
1.0 -0.14 0 1.5 5.5e-08 
1.0 -0.12 0 1.5 5.5e-08 
1.0 -0.1 0 1.5 5.5e-08 
1.0 -0.08 0 1.5 5.5e-08 
1.0 -0.06 0 1.5 5.5e-08 
1.0 -0.04 0 1.5 5.5e-08 
1.0 -0.02 0 1.5 5.5e-08 
1.0 1.33226762955e-15 0 1.5 5.5e-08 
1.0 0.02 0 1.5 5.5e-08 
1.0 0.04 0 1.5 5.5e-08 
1.0 0.06 0 1.5 5.5e-08 
1.0 0.08 0 1.5 5.5e-08 
1.0 0.1 0 1.5 5.5e-08 
1.0 0.12 0 1.5 5.5e-08 
1.0 0.14 0 1.5 5.5e-08 
1.0 0.16 0 1.5 5.5e-08 
1.0 0.18 0 1.5 5.5e-08 
1.0 0.2 0 1.5 5.5e-08 
1.0 0.22 0 1.5 5.5e-08 
1.0 0.24 0 1.5 5.5e-08 
1.0 0.26 0 1.5 5.5e-08 
1.0 0.28 0 1.5 5.5e-08 
1.0 0.3 0 1.5 5.5e-08 
1.0 0.32 0 1.5 5.5e-08 
1.0 0.34 0 1.5 5.5e-08 
1.0 0.36 0 1.5 5.5e-08 
1.0 0.38 0 1.5 5.5e-08 
1.0 0.4 0 1.5 5.5e-08 
1.0 0.42 0 1.5 5.5e-08 
1.0 0.44 0 1.5 5.5e-08 
1.0 0.46 0 1.5 5.5e-08 
1.0 0.48 0 1.5 5.5e-08 
1.0 0.5 0 1.5 5.5e-08 
1.0 0.52 0 1.5 5.5e-08 
1.0 0.54 0 1.5 5.5e-08 
1.0 0.56 0 1.5 5.5e-08 
1.0 0.58 0 1.5 5.5e-08 
1.0 0.6 0 1.5 5.5e-08 
1.0 0.62 0 1.5 5.5e-08 
1.0 0.64 0 1.5 5.5e-08 
1.0 0.66 0 1.5 5.5e-08 
1.0 0.68 0 1.5 5.5e-08 
1.0 0.7 0 1.5 5.5e-08 
1.0 0.72 0 1.5 5.5e-08 
1.0 0.74 0 1.5 5.5e-08 
1.0 0.76 0 1.5 5.5e-08 
1.0 0.78 0 1.5 5.5e-08 
1.0 0.8 0 1.5 5.5e-08 
1.0 0.82 0 1.5 5.5e-08 
1.0 0.84 0 1.5 5.5e-08 
1.0 0.86 0 1.5 5.5e-08 
1.0 0.88 0 1.5 5.5e-08 
1.0 0.9 0 1.5 5.5e-08 
1.0 0.92 0 1.5 5.5e-08 
1.0 0.94 0 1.5 5.5e-08 
1.0 0.96 0 1.5 5.5e-08 
1.0 0.98 0 1.5 5.5e-08 
1.0 1.0 0 1.5 5.5e-08 
1.0 1.02 0 1.5 5.5e-08 
1.0 1.04 0 1.5 5.5e-08 
1.0 1.06 0 1.5 5.5e-08 
1.0 1.08 0 1.5 5.5e-08 
1.0 1.1 0 1.5 5.5e-08 
1.0 1.12 0 1.5 5.5e-08 
1.0 1.14 0 1.5 5.5e-08 
1.0 1.16 0 1.5 5.5e-08 
1.0 1.18 0 1.5 5.5e-08 
1.0 1.2 0 1.5 5.5e-08 
1.0 1.22 0 1.5 5.5e-08 
1.0 1.24 0 1.5 5.5e-08 
1.0 1.26 0 1.5 5.5e-08 
1.0 1.28 0 1.5 5.5e-08 
1.0 1.3 0 1.5 5.5e-08 
1.0 1.32 0 1.5 5.5e-08 
1.0 1.34 0 1.5 5.5e-08 
1.0 1.36 0 1.5 5.5e-08 
1.0 1.38 0 1.5 5.5e-08 
1.0 1.4 0 1.5 5.5e-08 
1.0 1.42 0 1.5 5.5e-08 
1.0 1.44 0 1.5 5.5e-08 
1.0 1.46 0 1.5 5.5e-08 
1.0 1.48 0 1.5 5.5e-08 
1.0 -1.5 0 1.0 5.5e-08 
1.0 -1.48 0 1.0 5.5e-08 
1.0 -1.46 0 1.0 5.5e-08 
1.0 -1.44 0 1.0 5.5e-08 
1.0 -1.42 0 1.0 5.5e-08 
1.0 -1.4 0 1.0 5.5e-08 
1.0 -1.38 0 1.0 5.5e-08 
1.0 -1.36 0 1.0 5.5e-08 
1.0 -1.34 0 1.0 5.5e-08 
1.0 -1.32 0 1.0 5.5e-08 
1.0 -1.3 0 1.0 5.5e-08 
1.0 -1.28 0 1.0 5.5e-08 
1.0 -1.26 0 1.0 5.5e-08 
1.0 -1.24 0 1.0 5.5e-08 
1.0 -1.22 0 1.0 5.5e-08 
1.0 -1.2 0 1.0 5.5e-08 
1.0 -1.18 0 1.0 5.5e-08 
1.0 -1.16 0 1.0 5.5e-08 
1.0 -1.14 0 1.0 5.5e-08 
1.0 -1.12 0 1.0 5.5e-08 
1.0 -1.1 0 1.0 5.5e-08 
1.0 -1.08 0 1.0 5.5e-08 
1.0 -1.06 0 1.0 5.5e-08 
1.0 -1.04 0 1.0 5.5e-08 
1.0 -1.02 0 1.0 5.5e-08 
1.0 -1.0 0 1.0 5.5e-08 
1.0 -0.98 0 1.0 5.5e-08 
1.0 -0.96 0 1.0 5.5e-08 
1.0 -0.94 0 1.0 5.5e-08 
1.0 -0.92 0 1.0 5.5e-08 
1.0 -0.9 0 1.0 5.5e-08 
1.0 -0.88 0 1.0 5.5e-08 
1.0 -0.86 0 1.0 5.5e-08 
1.0 -0.84 0 1.0 5.5e-08 
1.0 -0.82 0 1.0 5.5e-08 
1.0 -0.8 0 1.0 5.5e-08 
1.0 -0.78 0 1.0 5.5e-08 
1.0 -0.76 0 1.0 5.5e-08 
1.0 -0.74 0 1.0 5.5e-08 
1.0 -0.72 0 1.0 5.5e-08 
1.0 -0.7 0 1.0 5.5e-08 
1.0 -0.68 0 1.0 5.5e-08 
1.0 -0.66 0 1.0 5.5e-08 
1.0 -0.64 0 1.0 5.5e-08 
1.0 -0.62 0 1.0 5.5e-08 
1.0 -0.6 0 1.0 5.5e-08 
1.0 -0.58 0 1.0 5.5e-08 
1.0 -0.56 0 1.0 5.5e-08 
1.0 -0.54 0 1.0 5.5e-08 
1.0 -0.52 0 1.0 5.5e-08 
1.0 -0.5 0 1.0 5.5e-08 
1.0 -0.48 0 1.0 5.5e-08 
1.0 -0.46 0 1.0 5.5e-08 
1.0 -0.44 0 1.0 5.5e-08 
1.0 -0.42 0 1.0 5.5e-08 
1.0 -0.4 0 1.0 5.5e-08 
1.0 -0.38 0 1.0 5.5e-08 
1.0 -0.36 0 1.0 5.5e-08 
1.0 -0.34 0 1.0 5.5e-08 
1.0 -0.32 0 1.0 5.5e-08 
1.0 -0.3 0 1.0 5.5e-08 
1.0 -0.28 0 1.0 5.5e-08 
1.0 -0.26 0 1.0 5.5e-08 
1.0 -0.24 0 1.0 5.5e-08 
1.0 -0.22 0 1.0 5.5e-08 
1.0 -0.2 0 1.0 5.5e-08 
1.0 -0.18 0 1.0 5.5e-08 
1.0 -0.16 0 1.0 5.5e-08 
1.0 -0.14 0 1.0 5.5e-08 
1.0 -0.12 0 1.0 5.5e-08 
1.0 -0.1 0 1.0 5.5e-08 
1.0 -0.08 0 1.0 5.5e-08 
1.0 -0.06 0 1.0 5.5e-08 
1.0 -0.04 0 1.0 5.5e-08 
1.0 -0.02 0 1.0 5.5e-08 
1.0 1.33226762955e-15 0 1.0 5.5e-08 
1.0 0.02 0 1.0 5.5e-08 
1.0 0.04 0 1.0 5.5e-08 
1.0 0.06 0 1.0 5.5e-08 
1.0 0.08 0 1.0 5.5e-08 
1.0 0.1 0 1.0 5.5e-08 
1.0 0.12 0 1.0 5.5e-08 
1.0 0.14 0 1.0 5.5e-08 
1.0 0.16 0 1.0 5.5e-08 
1.0 0.18 0 1.0 5.5e-08 
1.0 0.2 0 1.0 5.5e-08 
1.0 0.22 0 1.0 5.5e-08 
1.0 0.24 0 1.0 5.5e-08 
1.0 0.26 0 1.0 5.5e-08 
1.0 0.28 0 1.0 5.5e-08 
1.0 0.3 0 1.0 5.5e-08 
1.0 0.32 0 1.0 5.5e-08 
1.0 0.34 0 1.0 5.5e-08 
1.0 0.36 0 1.0 5.5e-08 
1.0 0.38 0 1.0 5.5e-08 
1.0 0.4 0 1.0 5.5e-08 
1.0 0.42 0 1.0 5.5e-08 
1.0 0.44 0 1.0 5.5e-08 
1.0 0.46 0 1.0 5.5e-08 
1.0 0.48 0 1.0 5.5e-08 
1.0 0.5 0 1.0 5.5e-08 
1.0 0.52 0 1.0 5.5e-08 
1.0 0.54 0 1.0 5.5e-08 
1.0 0.56 0 1.0 5.5e-08 
1.0 0.58 0 1.0 5.5e-08 
1.0 0.6 0 1.0 5.5e-08 
1.0 0.62 0 1.0 5.5e-08 
1.0 0.64 0 1.0 5.5e-08 
1.0 0.66 0 1.0 5.5e-08 
1.0 0.68 0 1.0 5.5e-08 
1.0 0.7 0 1.0 5.5e-08 
1.0 0.72 0 1.0 5.5e-08 
1.0 0.74 0 1.0 5.5e-08 
1.0 0.76 0 1.0 5.5e-08 
1.0 0.78 0 1.0 5.5e-08 
1.0 0.8 0 1.0 5.5e-08 
1.0 0.82 0 1.0 5.5e-08 
1.0 0.84 0 1.0 5.5e-08 
1.0 0.86 0 1.0 5.5e-08 
1.0 0.88 0 1.0 5.5e-08 
1.0 0.9 0 1.0 5.5e-08 
1.0 0.92 0 1.0 5.5e-08 
1.0 0.94 0 1.0 5.5e-08 
1.0 0.96 0 1.0 5.5e-08 
1.0 0.98 0 1.0 5.5e-08 
1.0 1.0 0 1.0 5.5e-08 
1.0 1.02 0 1.0 5.5e-08 
1.0 1.04 0 1.0 5.5e-08 
1.0 1.06 0 1.0 5.5e-08 
1.0 1.08 0 1.0 5.5e-08 
1.0 1.1 0 1.0 5.5e-08 
1.0 1.12 0 1.0 5.5e-08 
1.0 1.14 0 1.0 5.5e-08 
1.0 1.16 0 1.0 5.5e-08 
1.0 1.18 0 1.0 5.5e-08 
1.0 1.2 0 1.0 5.5e-08 
1.0 1.22 0 1.0 5.5e-08 
1.0 1.24 0 1.0 5.5e-08 
1.0 1.26 0 1.0 5.5e-08 
1.0 1.28 0 1.0 5.5e-08 
1.0 1.3 0 1.0 5.5e-08 
1.0 1.32 0 1.0 5.5e-08 
1.0 1.34 0 1.0 5.5e-08 
1.0 1.36 0 1.0 5.5e-08 
1.0 1.38 0 1.0 5.5e-08 
1.0 1.4 0 1.0 5.5e-08 
1.0 1.42 0 1.0 5.5e-08 
1.0 1.44 0 1.0 5.5e-08 
1.0 1.46 0 1.0 5.5e-08 
1.0 1.48 0 1.0 5.5e-08 
1.0 -1.5 0 0.5 5.5e-08 
1.0 -1.48 0 0.5 5.5e-08 
1.0 -1.46 0 0.5 5.5e-08 
1.0 -1.44 0 0.5 5.5e-08 
1.0 -1.42 0 0.5 5.5e-08 
1.0 -1.4 0 0.5 5.5e-08 
1.0 -1.38 0 0.5 5.5e-08 
1.0 -1.36 0 0.5 5.5e-08 
1.0 -1.34 0 0.5 5.5e-08 
1.0 -1.32 0 0.5 5.5e-08 
1.0 -1.3 0 0.5 5.5e-08 
1.0 -1.28 0 0.5 5.5e-08 
1.0 -1.26 0 0.5 5.5e-08 
1.0 -1.24 0 0.5 5.5e-08 
1.0 -1.22 0 0.5 5.5e-08 
1.0 -1.2 0 0.5 5.5e-08 
1.0 -1.18 0 0.5 5.5e-08 
1.0 -1.16 0 0.5 5.5e-08 
1.0 -1.14 0 0.5 5.5e-08 
1.0 -1.12 0 0.5 5.5e-08 
1.0 -1.1 0 0.5 5.5e-08 
1.0 -1.08 0 0.5 5.5e-08 
1.0 -1.06 0 0.5 5.5e-08 
1.0 -1.04 0 0.5 5.5e-08 
1.0 -1.02 0 0.5 5.5e-08 
1.0 -1.0 0 0.5 5.5e-08 
1.0 -0.98 0 0.5 5.5e-08 
1.0 -0.96 0 0.5 5.5e-08 
1.0 -0.94 0 0.5 5.5e-08 
1.0 -0.92 0 0.5 5.5e-08 
1.0 -0.9 0 0.5 5.5e-08 
1.0 -0.88 0 0.5 5.5e-08 
1.0 -0.86 0 0.5 5.5e-08 
1.0 -0.84 0 0.5 5.5e-08 
1.0 -0.82 0 0.5 5.5e-08 
1.0 -0.8 0 0.5 5.5e-08 
1.0 -0.78 0 0.5 5.5e-08 
1.0 -0.76 0 0.5 5.5e-08 
1.0 -0.74 0 0.5 5.5e-08 
1.0 -0.72 0 0.5 5.5e-08 
1.0 -0.7 0 0.5 5.5e-08 
1.0 -0.68 0 0.5 5.5e-08 
1.0 -0.66 0 0.5 5.5e-08 
1.0 -0.64 0 0.5 5.5e-08 
1.0 -0.62 0 0.5 5.5e-08 
1.0 -0.6 0 0.5 5.5e-08 
1.0 -0.58 0 0.5 5.5e-08 
1.0 -0.56 0 0.5 5.5e-08 
1.0 -0.54 0 0.5 5.5e-08 
1.0 -0.52 0 0.5 5.5e-08 
1.0 -0.5 0 0.5 5.5e-08 
1.0 -0.48 0 0.5 5.5e-08 
1.0 -0.46 0 0.5 5.5e-08 
1.0 -0.44 0 0.5 5.5e-08 
1.0 -0.42 0 0.5 5.5e-08 
1.0 -0.4 0 0.5 5.5e-08 
1.0 -0.38 0 0.5 5.5e-08 
1.0 -0.36 0 0.5 5.5e-08 
1.0 -0.34 0 0.5 5.5e-08 
1.0 -0.32 0 0.5 5.5e-08 
1.0 -0.3 0 0.5 5.5e-08 
1.0 -0.28 0 0.5 5.5e-08 
1.0 -0.26 0 0.5 5.5e-08 
1.0 -0.24 0 0.5 5.5e-08 
1.0 -0.22 0 0.5 5.5e-08 
1.0 -0.2 0 0.5 5.5e-08 
1.0 -0.18 0 0.5 5.5e-08 
1.0 -0.16 0 0.5 5.5e-08 
1.0 -0.14 0 0.5 5.5e-08 
1.0 -0.12 0 0.5 5.5e-08 
1.0 -0.1 0 0.5 5.5e-08 
1.0 -0.08 0 0.5 5.5e-08 
1.0 -0.06 0 0.5 5.5e-08 
1.0 -0.04 0 0.5 5.5e-08 
1.0 -0.02 0 0.5 5.5e-08 
1.0 1.33226762955e-15 0 0.5 5.5e-08 
1.0 0.02 0 0.5 5.5e-08 
1.0 0.04 0 0.5 5.5e-08 
1.0 0.06 0 0.5 5.5e-08 
1.0 0.08 0 0.5 5.5e-08 
1.0 0.1 0 0.5 5.5e-08 
1.0 0.12 0 0.5 5.5e-08 
1.0 0.14 0 0.5 5.5e-08 
1.0 0.16 0 0.5 5.5e-08 
1.0 0.18 0 0.5 5.5e-08 
1.0 0.2 0 0.5 5.5e-08 
1.0 0.22 0 0.5 5.5e-08 
1.0 0.24 0 0.5 5.5e-08 
1.0 0.26 0 0.5 5.5e-08 
1.0 0.28 0 0.5 5.5e-08 
1.0 0.3 0 0.5 5.5e-08 
1.0 0.32 0 0.5 5.5e-08 
1.0 0.34 0 0.5 5.5e-08 
1.0 0.36 0 0.5 5.5e-08 
1.0 0.38 0 0.5 5.5e-08 
1.0 0.4 0 0.5 5.5e-08 
1.0 0.42 0 0.5 5.5e-08 
1.0 0.44 0 0.5 5.5e-08 
1.0 0.46 0 0.5 5.5e-08 
1.0 0.48 0 0.5 5.5e-08 
1.0 0.5 0 0.5 5.5e-08 
1.0 0.52 0 0.5 5.5e-08 
1.0 0.54 0 0.5 5.5e-08 
1.0 0.56 0 0.5 5.5e-08 
1.0 0.58 0 0.5 5.5e-08 
1.0 0.6 0 0.5 5.5e-08 
1.0 0.62 0 0.5 5.5e-08 
1.0 0.64 0 0.5 5.5e-08 
1.0 0.66 0 0.5 5.5e-08 
1.0 0.68 0 0.5 5.5e-08 
1.0 0.7 0 0.5 5.5e-08 
1.0 0.72 0 0.5 5.5e-08 
1.0 0.74 0 0.5 5.5e-08 
1.0 0.76 0 0.5 5.5e-08 
1.0 0.78 0 0.5 5.5e-08 
1.0 0.8 0 0.5 5.5e-08 
1.0 0.82 0 0.5 5.5e-08 
1.0 0.84 0 0.5 5.5e-08 
1.0 0.86 0 0.5 5.5e-08 
1.0 0.88 0 0.5 5.5e-08 
1.0 0.9 0 0.5 5.5e-08 
1.0 0.92 0 0.5 5.5e-08 
1.0 0.94 0 0.5 5.5e-08 
1.0 0.96 0 0.5 5.5e-08 
1.0 0.98 0 0.5 5.5e-08 
1.0 1.0 0 0.5 5.5e-08 
1.0 1.02 0 0.5 5.5e-08 
1.0 1.04 0 0.5 5.5e-08 
1.0 1.06 0 0.5 5.5e-08 
1.0 1.08 0 0.5 5.5e-08 
1.0 1.1 0 0.5 5.5e-08 
1.0 1.12 0 0.5 5.5e-08 
1.0 1.14 0 0.5 5.5e-08 
1.0 1.16 0 0.5 5.5e-08 
1.0 1.18 0 0.5 5.5e-08 
1.0 1.2 0 0.5 5.5e-08 
1.0 1.22 0 0.5 5.5e-08 
1.0 1.24 0 0.5 5.5e-08 
1.0 1.26 0 0.5 5.5e-08 
1.0 1.28 0 0.5 5.5e-08 
1.0 1.3 0 0.5 5.5e-08 
1.0 1.32 0 0.5 5.5e-08 
1.0 1.34 0 0.5 5.5e-08 
1.0 1.36 0 0.5 5.5e-08 
1.0 1.38 0 0.5 5.5e-08 
1.0 1.4 0 0.5 5.5e-08 
1.0 1.42 0 0.5 5.5e-08 
1.0 1.44 0 0.5 5.5e-08 
1.0 1.46 0 0.5 5.5e-08 
1.0 1.48 0 0.5 5.5e-08 
1.0 -1.5 0 0.0 5.5e-08 
1.0 -1.48 0 0.0 5.5e-08 
1.0 -1.46 0 0.0 5.5e-08 
1.0 -1.44 0 0.0 5.5e-08 
1.0 -1.42 0 0.0 5.5e-08 
1.0 -1.4 0 0.0 5.5e-08 
1.0 -1.38 0 0.0 5.5e-08 
1.0 -1.36 0 0.0 5.5e-08 
1.0 -1.34 0 0.0 5.5e-08 
1.0 -1.32 0 0.0 5.5e-08 
1.0 -1.3 0 0.0 5.5e-08 
1.0 -1.28 0 0.0 5.5e-08 
1.0 -1.26 0 0.0 5.5e-08 
1.0 -1.24 0 0.0 5.5e-08 
1.0 -1.22 0 0.0 5.5e-08 
1.0 -1.2 0 0.0 5.5e-08 
1.0 -1.18 0 0.0 5.5e-08 
1.0 -1.16 0 0.0 5.5e-08 
1.0 -1.14 0 0.0 5.5e-08 
1.0 -1.12 0 0.0 5.5e-08 
1.0 -1.1 0 0.0 5.5e-08 
1.0 -1.08 0 0.0 5.5e-08 
1.0 -1.06 0 0.0 5.5e-08 
1.0 -1.04 0 0.0 5.5e-08 
1.0 -1.02 0 0.0 5.5e-08 
1.0 -1.0 0 0.0 5.5e-08 
1.0 -0.98 0 0.0 5.5e-08 
1.0 -0.96 0 0.0 5.5e-08 
1.0 -0.94 0 0.0 5.5e-08 
1.0 -0.92 0 0.0 5.5e-08 
1.0 -0.9 0 0.0 5.5e-08 
1.0 -0.88 0 0.0 5.5e-08 
1.0 -0.86 0 0.0 5.5e-08 
1.0 -0.84 0 0.0 5.5e-08 
1.0 -0.82 0 0.0 5.5e-08 
1.0 -0.8 0 0.0 5.5e-08 
1.0 -0.78 0 0.0 5.5e-08 
1.0 -0.76 0 0.0 5.5e-08 
1.0 -0.74 0 0.0 5.5e-08 
1.0 -0.72 0 0.0 5.5e-08 
1.0 -0.7 0 0.0 5.5e-08 
1.0 -0.68 0 0.0 5.5e-08 
1.0 -0.66 0 0.0 5.5e-08 
1.0 -0.64 0 0.0 5.5e-08 
1.0 -0.62 0 0.0 5.5e-08 
1.0 -0.6 0 0.0 5.5e-08 
1.0 -0.58 0 0.0 5.5e-08 
1.0 -0.56 0 0.0 5.5e-08 
1.0 -0.54 0 0.0 5.5e-08 
1.0 -0.52 0 0.0 5.5e-08 
1.0 -0.5 0 0.0 5.5e-08 
1.0 -0.48 0 0.0 5.5e-08 
1.0 -0.46 0 0.0 5.5e-08 
1.0 -0.44 0 0.0 5.5e-08 
1.0 -0.42 0 0.0 5.5e-08 
1.0 -0.4 0 0.0 5.5e-08 
1.0 -0.38 0 0.0 5.5e-08 
1.0 -0.36 0 0.0 5.5e-08 
1.0 -0.34 0 0.0 5.5e-08 
1.0 -0.32 0 0.0 5.5e-08 
1.0 -0.3 0 0.0 5.5e-08 
1.0 -0.28 0 0.0 5.5e-08 
1.0 -0.26 0 0.0 5.5e-08 
1.0 -0.24 0 0.0 5.5e-08 
1.0 -0.22 0 0.0 5.5e-08 
1.0 -0.2 0 0.0 5.5e-08 
1.0 -0.18 0 0.0 5.5e-08 
1.0 -0.16 0 0.0 5.5e-08 
1.0 -0.14 0 0.0 5.5e-08 
1.0 -0.12 0 0.0 5.5e-08 
1.0 -0.1 0 0.0 5.5e-08 
1.0 -0.08 0 0.0 5.5e-08 
1.0 -0.06 0 0.0 5.5e-08 
1.0 -0.04 0 0.0 5.5e-08 
1.0 -0.02 0 0.0 5.5e-08 
1.0 1.33226762955e-15 0 0.0 5.5e-08 
1.0 0.02 0 0.0 5.5e-08 
1.0 0.04 0 0.0 5.5e-08 
1.0 0.06 0 0.0 5.5e-08 
1.0 0.08 0 0.0 5.5e-08 
1.0 0.1 0 0.0 5.5e-08 
1.0 0.12 0 0.0 5.5e-08 
1.0 0.14 0 0.0 5.5e-08 
1.0 0.16 0 0.0 5.5e-08 
1.0 0.18 0 0.0 5.5e-08 
1.0 0.2 0 0.0 5.5e-08 
1.0 0.22 0 0.0 5.5e-08 
1.0 0.24 0 0.0 5.5e-08 
1.0 0.26 0 0.0 5.5e-08 
1.0 0.28 0 0.0 5.5e-08 
1.0 0.3 0 0.0 5.5e-08 
1.0 0.32 0 0.0 5.5e-08 
1.0 0.34 0 0.0 5.5e-08 
1.0 0.36 0 0.0 5.5e-08 
1.0 0.38 0 0.0 5.5e-08 
1.0 0.4 0 0.0 5.5e-08 
1.0 0.42 0 0.0 5.5e-08 
1.0 0.44 0 0.0 5.5e-08 
1.0 0.46 0 0.0 5.5e-08 
1.0 0.48 0 0.0 5.5e-08 
1.0 0.5 0 0.0 5.5e-08 
1.0 0.52 0 0.0 5.5e-08 
1.0 0.54 0 0.0 5.5e-08 
1.0 0.56 0 0.0 5.5e-08 
1.0 0.58 0 0.0 5.5e-08 
1.0 0.6 0 0.0 5.5e-08 
1.0 0.62 0 0.0 5.5e-08 
1.0 0.64 0 0.0 5.5e-08 
1.0 0.66 0 0.0 5.5e-08 
1.0 0.68 0 0.0 5.5e-08 
1.0 0.7 0 0.0 5.5e-08 
1.0 0.72 0 0.0 5.5e-08 
1.0 0.74 0 0.0 5.5e-08 
1.0 0.76 0 0.0 5.5e-08 
1.0 0.78 0 0.0 5.5e-08 
1.0 0.8 0 0.0 5.5e-08 
1.0 0.82 0 0.0 5.5e-08 
1.0 0.84 0 0.0 5.5e-08 
1.0 0.86 0 0.0 5.5e-08 
1.0 0.88 0 0.0 5.5e-08 
1.0 0.9 0 0.0 5.5e-08 
1.0 0.92 0 0.0 5.5e-08 
1.0 0.94 0 0.0 5.5e-08 
1.0 0.96 0 0.0 5.5e-08 
1.0 0.98 0 0.0 5.5e-08 
1.0 1.0 0 0.0 5.5e-08 
1.0 1.02 0 0.0 5.5e-08 
1.0 1.04 0 0.0 5.5e-08 
1.0 1.06 0 0.0 5.5e-08 
1.0 1.08 0 0.0 5.5e-08 
1.0 1.1 0 0.0 5.5e-08 
1.0 1.12 0 0.0 5.5e-08 
1.0 1.14 0 0.0 5.5e-08 
1.0 1.16 0 0.0 5.5e-08 
1.0 1.18 0 0.0 5.5e-08 
1.0 1.2 0 0.0 5.5e-08 
1.0 1.22 0 0.0 5.5e-08 
1.0 1.24 0 0.0 5.5e-08 
1.0 1.26 0 0.0 5.5e-08 
1.0 1.28 0 0.0 5.5e-08 
1.0 1.3 0 0.0 5.5e-08 
1.0 1.32 0 0.0 5.5e-08 
1.0 1.34 0 0.0 5.5e-08 
1.0 1.36 0 0.0 5.5e-08 
1.0 1.38 0 0.0 5.5e-08 
1.0 1.4 0 0.0 5.5e-08 
1.0 1.42 0 0.0 5.5e-08 
1.0 1.44 0 0.0 5.5e-08 
1.0 1.46 0 0.0 5.5e-08 
1.0 1.48 0 0.0 5.5e-08 
1.0 -1.5 0 -0.5 5.5e-08 
1.0 -1.48 0 -0.5 5.5e-08 
1.0 -1.46 0 -0.5 5.5e-08 
1.0 -1.44 0 -0.5 5.5e-08 
1.0 -1.42 0 -0.5 5.5e-08 
1.0 -1.4 0 -0.5 5.5e-08 
1.0 -1.38 0 -0.5 5.5e-08 
1.0 -1.36 0 -0.5 5.5e-08 
1.0 -1.34 0 -0.5 5.5e-08 
1.0 -1.32 0 -0.5 5.5e-08 
1.0 -1.3 0 -0.5 5.5e-08 
1.0 -1.28 0 -0.5 5.5e-08 
1.0 -1.26 0 -0.5 5.5e-08 
1.0 -1.24 0 -0.5 5.5e-08 
1.0 -1.22 0 -0.5 5.5e-08 
1.0 -1.2 0 -0.5 5.5e-08 
1.0 -1.18 0 -0.5 5.5e-08 
1.0 -1.16 0 -0.5 5.5e-08 
1.0 -1.14 0 -0.5 5.5e-08 
1.0 -1.12 0 -0.5 5.5e-08 
1.0 -1.1 0 -0.5 5.5e-08 
1.0 -1.08 0 -0.5 5.5e-08 
1.0 -1.06 0 -0.5 5.5e-08 
1.0 -1.04 0 -0.5 5.5e-08 
1.0 -1.02 0 -0.5 5.5e-08 
1.0 -1.0 0 -0.5 5.5e-08 
1.0 -0.98 0 -0.5 5.5e-08 
1.0 -0.96 0 -0.5 5.5e-08 
1.0 -0.94 0 -0.5 5.5e-08 
1.0 -0.92 0 -0.5 5.5e-08 
1.0 -0.9 0 -0.5 5.5e-08 
1.0 -0.88 0 -0.5 5.5e-08 
1.0 -0.86 0 -0.5 5.5e-08 
1.0 -0.84 0 -0.5 5.5e-08 
1.0 -0.82 0 -0.5 5.5e-08 
1.0 -0.8 0 -0.5 5.5e-08 
1.0 -0.78 0 -0.5 5.5e-08 
1.0 -0.76 0 -0.5 5.5e-08 
1.0 -0.74 0 -0.5 5.5e-08 
1.0 -0.72 0 -0.5 5.5e-08 
1.0 -0.7 0 -0.5 5.5e-08 
1.0 -0.68 0 -0.5 5.5e-08 
1.0 -0.66 0 -0.5 5.5e-08 
1.0 -0.64 0 -0.5 5.5e-08 
1.0 -0.62 0 -0.5 5.5e-08 
1.0 -0.6 0 -0.5 5.5e-08 
1.0 -0.58 0 -0.5 5.5e-08 
1.0 -0.56 0 -0.5 5.5e-08 
1.0 -0.54 0 -0.5 5.5e-08 
1.0 -0.52 0 -0.5 5.5e-08 
1.0 -0.5 0 -0.5 5.5e-08 
1.0 -0.48 0 -0.5 5.5e-08 
1.0 -0.46 0 -0.5 5.5e-08 
1.0 -0.44 0 -0.5 5.5e-08 
1.0 -0.42 0 -0.5 5.5e-08 
1.0 -0.4 0 -0.5 5.5e-08 
1.0 -0.38 0 -0.5 5.5e-08 
1.0 -0.36 0 -0.5 5.5e-08 
1.0 -0.34 0 -0.5 5.5e-08 
1.0 -0.32 0 -0.5 5.5e-08 
1.0 -0.3 0 -0.5 5.5e-08 
1.0 -0.28 0 -0.5 5.5e-08 
1.0 -0.26 0 -0.5 5.5e-08 
1.0 -0.24 0 -0.5 5.5e-08 
1.0 -0.22 0 -0.5 5.5e-08 
1.0 -0.2 0 -0.5 5.5e-08 
1.0 -0.18 0 -0.5 5.5e-08 
1.0 -0.16 0 -0.5 5.5e-08 
1.0 -0.14 0 -0.5 5.5e-08 
1.0 -0.12 0 -0.5 5.5e-08 
1.0 -0.1 0 -0.5 5.5e-08 
1.0 -0.08 0 -0.5 5.5e-08 
1.0 -0.06 0 -0.5 5.5e-08 
1.0 -0.04 0 -0.5 5.5e-08 
1.0 -0.02 0 -0.5 5.5e-08 
1.0 1.33226762955e-15 0 -0.5 5.5e-08 
1.0 0.02 0 -0.5 5.5e-08 
1.0 0.04 0 -0.5 5.5e-08 
1.0 0.06 0 -0.5 5.5e-08 
1.0 0.08 0 -0.5 5.5e-08 
1.0 0.1 0 -0.5 5.5e-08 
1.0 0.12 0 -0.5 5.5e-08 
1.0 0.14 0 -0.5 5.5e-08 
1.0 0.16 0 -0.5 5.5e-08 
1.0 0.18 0 -0.5 5.5e-08 
1.0 0.2 0 -0.5 5.5e-08 
1.0 0.22 0 -0.5 5.5e-08 
1.0 0.24 0 -0.5 5.5e-08 
1.0 0.26 0 -0.5 5.5e-08 
1.0 0.28 0 -0.5 5.5e-08 
1.0 0.3 0 -0.5 5.5e-08 
1.0 0.32 0 -0.5 5.5e-08 
1.0 0.34 0 -0.5 5.5e-08 
1.0 0.36 0 -0.5 5.5e-08 
1.0 0.38 0 -0.5 5.5e-08 
1.0 0.4 0 -0.5 5.5e-08 
1.0 0.42 0 -0.5 5.5e-08 
1.0 0.44 0 -0.5 5.5e-08 
1.0 0.46 0 -0.5 5.5e-08 
1.0 0.48 0 -0.5 5.5e-08 
1.0 0.5 0 -0.5 5.5e-08 
1.0 0.52 0 -0.5 5.5e-08 
1.0 0.54 0 -0.5 5.5e-08 
1.0 0.56 0 -0.5 5.5e-08 
1.0 0.58 0 -0.5 5.5e-08 
1.0 0.6 0 -0.5 5.5e-08 
1.0 0.62 0 -0.5 5.5e-08 
1.0 0.64 0 -0.5 5.5e-08 
1.0 0.66 0 -0.5 5.5e-08 
1.0 0.68 0 -0.5 5.5e-08 
1.0 0.7 0 -0.5 5.5e-08 
1.0 0.72 0 -0.5 5.5e-08 
1.0 0.74 0 -0.5 5.5e-08 
1.0 0.76 0 -0.5 5.5e-08 
1.0 0.78 0 -0.5 5.5e-08 
1.0 0.8 0 -0.5 5.5e-08 
1.0 0.82 0 -0.5 5.5e-08 
1.0 0.84 0 -0.5 5.5e-08 
1.0 0.86 0 -0.5 5.5e-08 
1.0 0.88 0 -0.5 5.5e-08 
1.0 0.9 0 -0.5 5.5e-08 
1.0 0.92 0 -0.5 5.5e-08 
1.0 0.94 0 -0.5 5.5e-08 
1.0 0.96 0 -0.5 5.5e-08 
1.0 0.98 0 -0.5 5.5e-08 
1.0 1.0 0 -0.5 5.5e-08 
1.0 1.02 0 -0.5 5.5e-08 
1.0 1.04 0 -0.5 5.5e-08 
1.0 1.06 0 -0.5 5.5e-08 
1.0 1.08 0 -0.5 5.5e-08 
1.0 1.1 0 -0.5 5.5e-08 
1.0 1.12 0 -0.5 5.5e-08 
1.0 1.14 0 -0.5 5.5e-08 
1.0 1.16 0 -0.5 5.5e-08 
1.0 1.18 0 -0.5 5.5e-08 
1.0 1.2 0 -0.5 5.5e-08 
1.0 1.22 0 -0.5 5.5e-08 
1.0 1.24 0 -0.5 5.5e-08 
1.0 1.26 0 -0.5 5.5e-08 
1.0 1.28 0 -0.5 5.5e-08 
1.0 1.3 0 -0.5 5.5e-08 
1.0 1.32 0 -0.5 5.5e-08 
1.0 1.34 0 -0.5 5.5e-08 
1.0 1.36 0 -0.5 5.5e-08 
1.0 1.38 0 -0.5 5.5e-08 
1.0 1.4 0 -0.5 5.5e-08 
1.0 1.42 0 -0.5 5.5e-08 
1.0 1.44 0 -0.5 5.5e-08 
1.0 1.46 0 -0.5 5.5e-08 
1.0 1.48 0 -0.5 5.5e-08 
1.0 -1.5 0 -1.0 5.5e-08 
1.0 -1.48 0 -1.0 5.5e-08 
1.0 -1.46 0 -1.0 5.5e-08 
1.0 -1.44 0 -1.0 5.5e-08 
1.0 -1.42 0 -1.0 5.5e-08 
1.0 -1.4 0 -1.0 5.5e-08 
1.0 -1.38 0 -1.0 5.5e-08 
1.0 -1.36 0 -1.0 5.5e-08 
1.0 -1.34 0 -1.0 5.5e-08 
1.0 -1.32 0 -1.0 5.5e-08 
1.0 -1.3 0 -1.0 5.5e-08 
1.0 -1.28 0 -1.0 5.5e-08 
1.0 -1.26 0 -1.0 5.5e-08 
1.0 -1.24 0 -1.0 5.5e-08 
1.0 -1.22 0 -1.0 5.5e-08 
1.0 -1.2 0 -1.0 5.5e-08 
1.0 -1.18 0 -1.0 5.5e-08 
1.0 -1.16 0 -1.0 5.5e-08 
1.0 -1.14 0 -1.0 5.5e-08 
1.0 -1.12 0 -1.0 5.5e-08 
1.0 -1.1 0 -1.0 5.5e-08 
1.0 -1.08 0 -1.0 5.5e-08 
1.0 -1.06 0 -1.0 5.5e-08 
1.0 -1.04 0 -1.0 5.5e-08 
1.0 -1.02 0 -1.0 5.5e-08 
1.0 -1.0 0 -1.0 5.5e-08 
1.0 -0.98 0 -1.0 5.5e-08 
1.0 -0.96 0 -1.0 5.5e-08 
1.0 -0.94 0 -1.0 5.5e-08 
1.0 -0.92 0 -1.0 5.5e-08 
1.0 -0.9 0 -1.0 5.5e-08 
1.0 -0.88 0 -1.0 5.5e-08 
1.0 -0.86 0 -1.0 5.5e-08 
1.0 -0.84 0 -1.0 5.5e-08 
1.0 -0.82 0 -1.0 5.5e-08 
1.0 -0.8 0 -1.0 5.5e-08 
1.0 -0.78 0 -1.0 5.5e-08 
1.0 -0.76 0 -1.0 5.5e-08 
1.0 -0.74 0 -1.0 5.5e-08 
1.0 -0.72 0 -1.0 5.5e-08 
1.0 -0.7 0 -1.0 5.5e-08 
1.0 -0.68 0 -1.0 5.5e-08 
1.0 -0.66 0 -1.0 5.5e-08 
1.0 -0.64 0 -1.0 5.5e-08 
1.0 -0.62 0 -1.0 5.5e-08 
1.0 -0.6 0 -1.0 5.5e-08 
1.0 -0.58 0 -1.0 5.5e-08 
1.0 -0.56 0 -1.0 5.5e-08 
1.0 -0.54 0 -1.0 5.5e-08 
1.0 -0.52 0 -1.0 5.5e-08 
1.0 -0.5 0 -1.0 5.5e-08 
1.0 -0.48 0 -1.0 5.5e-08 
1.0 -0.46 0 -1.0 5.5e-08 
1.0 -0.44 0 -1.0 5.5e-08 
1.0 -0.42 0 -1.0 5.5e-08 
1.0 -0.4 0 -1.0 5.5e-08 
1.0 -0.38 0 -1.0 5.5e-08 
1.0 -0.36 0 -1.0 5.5e-08 
1.0 -0.34 0 -1.0 5.5e-08 
1.0 -0.32 0 -1.0 5.5e-08 
1.0 -0.3 0 -1.0 5.5e-08 
1.0 -0.28 0 -1.0 5.5e-08 
1.0 -0.26 0 -1.0 5.5e-08 
1.0 -0.24 0 -1.0 5.5e-08 
1.0 -0.22 0 -1.0 5.5e-08 
1.0 -0.2 0 -1.0 5.5e-08 
1.0 -0.18 0 -1.0 5.5e-08 
1.0 -0.16 0 -1.0 5.5e-08 
1.0 -0.14 0 -1.0 5.5e-08 
1.0 -0.12 0 -1.0 5.5e-08 
1.0 -0.1 0 -1.0 5.5e-08 
1.0 -0.08 0 -1.0 5.5e-08 
1.0 -0.06 0 -1.0 5.5e-08 
1.0 -0.04 0 -1.0 5.5e-08 
1.0 -0.02 0 -1.0 5.5e-08 
1.0 1.33226762955e-15 0 -1.0 5.5e-08 
1.0 0.02 0 -1.0 5.5e-08 
1.0 0.04 0 -1.0 5.5e-08 
1.0 0.06 0 -1.0 5.5e-08 
1.0 0.08 0 -1.0 5.5e-08 
1.0 0.1 0 -1.0 5.5e-08 
1.0 0.12 0 -1.0 5.5e-08 
1.0 0.14 0 -1.0 5.5e-08 
1.0 0.16 0 -1.0 5.5e-08 
1.0 0.18 0 -1.0 5.5e-08 
1.0 0.2 0 -1.0 5.5e-08 
1.0 0.22 0 -1.0 5.5e-08 
1.0 0.24 0 -1.0 5.5e-08 
1.0 0.26 0 -1.0 5.5e-08 
1.0 0.28 0 -1.0 5.5e-08 
1.0 0.3 0 -1.0 5.5e-08 
1.0 0.32 0 -1.0 5.5e-08 
1.0 0.34 0 -1.0 5.5e-08 
1.0 0.36 0 -1.0 5.5e-08 
1.0 0.38 0 -1.0 5.5e-08 
1.0 0.4 0 -1.0 5.5e-08 
1.0 0.42 0 -1.0 5.5e-08 
1.0 0.44 0 -1.0 5.5e-08 
1.0 0.46 0 -1.0 5.5e-08 
1.0 0.48 0 -1.0 5.5e-08 
1.0 0.5 0 -1.0 5.5e-08 
1.0 0.52 0 -1.0 5.5e-08 
1.0 0.54 0 -1.0 5.5e-08 
1.0 0.56 0 -1.0 5.5e-08 
1.0 0.58 0 -1.0 5.5e-08 
1.0 0.6 0 -1.0 5.5e-08 
1.0 0.62 0 -1.0 5.5e-08 
1.0 0.64 0 -1.0 5.5e-08 
1.0 0.66 0 -1.0 5.5e-08 
1.0 0.68 0 -1.0 5.5e-08 
1.0 0.7 0 -1.0 5.5e-08 
1.0 0.72 0 -1.0 5.5e-08 
1.0 0.74 0 -1.0 5.5e-08 
1.0 0.76 0 -1.0 5.5e-08 
1.0 0.78 0 -1.0 5.5e-08 
1.0 0.8 0 -1.0 5.5e-08 
1.0 0.82 0 -1.0 5.5e-08 
1.0 0.84 0 -1.0 5.5e-08 
1.0 0.86 0 -1.0 5.5e-08 
1.0 0.88 0 -1.0 5.5e-08 
1.0 0.9 0 -1.0 5.5e-08 
1.0 0.92 0 -1.0 5.5e-08 
1.0 0.94 0 -1.0 5.5e-08 
1.0 0.96 0 -1.0 5.5e-08 
1.0 0.98 0 -1.0 5.5e-08 
1.0 1.0 0 -1.0 5.5e-08 
1.0 1.02 0 -1.0 5.5e-08 
1.0 1.04 0 -1.0 5.5e-08 
1.0 1.06 0 -1.0 5.5e-08 
1.0 1.08 0 -1.0 5.5e-08 
1.0 1.1 0 -1.0 5.5e-08 
1.0 1.12 0 -1.0 5.5e-08 
1.0 1.14 0 -1.0 5.5e-08 
1.0 1.16 0 -1.0 5.5e-08 
1.0 1.18 0 -1.0 5.5e-08 
1.0 1.2 0 -1.0 5.5e-08 
1.0 1.22 0 -1.0 5.5e-08 
1.0 1.24 0 -1.0 5.5e-08 
1.0 1.26 0 -1.0 5.5e-08 
1.0 1.28 0 -1.0 5.5e-08 
1.0 1.3 0 -1.0 5.5e-08 
1.0 1.32 0 -1.0 5.5e-08 
1.0 1.34 0 -1.0 5.5e-08 
1.0 1.36 0 -1.0 5.5e-08 
1.0 1.38 0 -1.0 5.5e-08 
1.0 1.4 0 -1.0 5.5e-08 
1.0 1.42 0 -1.0 5.5e-08 
1.0 1.44 0 -1.0 5.5e-08 
1.0 1.46 0 -1.0 5.5e-08 
1.0 1.48 0 -1.0 5.5e-08 
1.0 -1.5 0 -1.5 5.5e-08 
1.0 -1.48 0 -1.5 5.5e-08 
1.0 -1.46 0 -1.5 5.5e-08 
1.0 -1.44 0 -1.5 5.5e-08 
1.0 -1.42 0 -1.5 5.5e-08 
1.0 -1.4 0 -1.5 5.5e-08 
1.0 -1.38 0 -1.5 5.5e-08 
1.0 -1.36 0 -1.5 5.5e-08 
1.0 -1.34 0 -1.5 5.5e-08 
1.0 -1.32 0 -1.5 5.5e-08 
1.0 -1.3 0 -1.5 5.5e-08 
1.0 -1.28 0 -1.5 5.5e-08 
1.0 -1.26 0 -1.5 5.5e-08 
1.0 -1.24 0 -1.5 5.5e-08 
1.0 -1.22 0 -1.5 5.5e-08 
1.0 -1.2 0 -1.5 5.5e-08 
1.0 -1.18 0 -1.5 5.5e-08 
1.0 -1.16 0 -1.5 5.5e-08 
1.0 -1.14 0 -1.5 5.5e-08 
1.0 -1.12 0 -1.5 5.5e-08 
1.0 -1.1 0 -1.5 5.5e-08 
1.0 -1.08 0 -1.5 5.5e-08 
1.0 -1.06 0 -1.5 5.5e-08 
1.0 -1.04 0 -1.5 5.5e-08 
1.0 -1.02 0 -1.5 5.5e-08 
1.0 -1.0 0 -1.5 5.5e-08 
1.0 -0.98 0 -1.5 5.5e-08 
1.0 -0.96 0 -1.5 5.5e-08 
1.0 -0.94 0 -1.5 5.5e-08 
1.0 -0.92 0 -1.5 5.5e-08 
1.0 -0.9 0 -1.5 5.5e-08 
1.0 -0.88 0 -1.5 5.5e-08 
1.0 -0.86 0 -1.5 5.5e-08 
1.0 -0.84 0 -1.5 5.5e-08 
1.0 -0.82 0 -1.5 5.5e-08 
1.0 -0.8 0 -1.5 5.5e-08 
1.0 -0.78 0 -1.5 5.5e-08 
1.0 -0.76 0 -1.5 5.5e-08 
1.0 -0.74 0 -1.5 5.5e-08 
1.0 -0.72 0 -1.5 5.5e-08 
1.0 -0.7 0 -1.5 5.5e-08 
1.0 -0.68 0 -1.5 5.5e-08 
1.0 -0.66 0 -1.5 5.5e-08 
1.0 -0.64 0 -1.5 5.5e-08 
1.0 -0.62 0 -1.5 5.5e-08 
1.0 -0.6 0 -1.5 5.5e-08 
1.0 -0.58 0 -1.5 5.5e-08 
1.0 -0.56 0 -1.5 5.5e-08 
1.0 -0.54 0 -1.5 5.5e-08 
1.0 -0.52 0 -1.5 5.5e-08 
1.0 -0.5 0 -1.5 5.5e-08 
1.0 -0.48 0 -1.5 5.5e-08 
1.0 -0.46 0 -1.5 5.5e-08 
1.0 -0.44 0 -1.5 5.5e-08 
1.0 -0.42 0 -1.5 5.5e-08 
1.0 -0.4 0 -1.5 5.5e-08 
1.0 -0.38 0 -1.5 5.5e-08 
1.0 -0.36 0 -1.5 5.5e-08 
1.0 -0.34 0 -1.5 5.5e-08 
1.0 -0.32 0 -1.5 5.5e-08 
1.0 -0.3 0 -1.5 5.5e-08 
1.0 -0.28 0 -1.5 5.5e-08 
1.0 -0.26 0 -1.5 5.5e-08 
1.0 -0.24 0 -1.5 5.5e-08 
1.0 -0.22 0 -1.5 5.5e-08 
1.0 -0.2 0 -1.5 5.5e-08 
1.0 -0.18 0 -1.5 5.5e-08 
1.0 -0.16 0 -1.5 5.5e-08 
1.0 -0.14 0 -1.5 5.5e-08 
1.0 -0.12 0 -1.5 5.5e-08 
1.0 -0.1 0 -1.5 5.5e-08 
1.0 -0.08 0 -1.5 5.5e-08 
1.0 -0.06 0 -1.5 5.5e-08 
1.0 -0.04 0 -1.5 5.5e-08 
1.0 -0.02 0 -1.5 5.5e-08 
1.0 1.33226762955e-15 0 -1.5 5.5e-08 
1.0 0.02 0 -1.5 5.5e-08 
1.0 0.04 0 -1.5 5.5e-08 
1.0 0.06 0 -1.5 5.5e-08 
1.0 0.08 0 -1.5 5.5e-08 
1.0 0.1 0 -1.5 5.5e-08 
1.0 0.12 0 -1.5 5.5e-08 
1.0 0.14 0 -1.5 5.5e-08 
1.0 0.16 0 -1.5 5.5e-08 
1.0 0.18 0 -1.5 5.5e-08 
1.0 0.2 0 -1.5 5.5e-08 
1.0 0.22 0 -1.5 5.5e-08 
1.0 0.24 0 -1.5 5.5e-08 
1.0 0.26 0 -1.5 5.5e-08 
1.0 0.28 0 -1.5 5.5e-08 
1.0 0.3 0 -1.5 5.5e-08 
1.0 0.32 0 -1.5 5.5e-08 
1.0 0.34 0 -1.5 5.5e-08 
1.0 0.36 0 -1.5 5.5e-08 
1.0 0.38 0 -1.5 5.5e-08 
1.0 0.4 0 -1.5 5.5e-08 
1.0 0.42 0 -1.5 5.5e-08 
1.0 0.44 0 -1.5 5.5e-08 
1.0 0.46 0 -1.5 5.5e-08 
1.0 0.48 0 -1.5 5.5e-08 
1.0 0.5 0 -1.5 5.5e-08 
1.0 0.52 0 -1.5 5.5e-08 
1.0 0.54 0 -1.5 5.5e-08 
1.0 0.56 0 -1.5 5.5e-08 
1.0 0.58 0 -1.5 5.5e-08 
1.0 0.6 0 -1.5 5.5e-08 
1.0 0.62 0 -1.5 5.5e-08 
1.0 0.64 0 -1.5 5.5e-08 
1.0 0.66 0 -1.5 5.5e-08 
1.0 0.68 0 -1.5 5.5e-08 
1.0 0.7 0 -1.5 5.5e-08 
1.0 0.72 0 -1.5 5.5e-08 
1.0 0.74 0 -1.5 5.5e-08 
1.0 0.76 0 -1.5 5.5e-08 
1.0 0.78 0 -1.5 5.5e-08 
1.0 0.8 0 -1.5 5.5e-08 
1.0 0.82 0 -1.5 5.5e-08 
1.0 0.84 0 -1.5 5.5e-08 
1.0 0.86 0 -1.5 5.5e-08 
1.0 0.88 0 -1.5 5.5e-08 
1.0 0.9 0 -1.5 5.5e-08 
1.0 0.92 0 -1.5 5.5e-08 
1.0 0.94 0 -1.5 5.5e-08 
1.0 0.96 0 -1.5 5.5e-08 
1.0 0.98 0 -1.5 5.5e-08 
1.0 1.0 0 -1.5 5.5e-08 
1.0 1.02 0 -1.5 5.5e-08 
1.0 1.04 0 -1.5 5.5e-08 
1.0 1.06 0 -1.5 5.5e-08 
1.0 1.08 0 -1.5 5.5e-08 
1.0 1.1 0 -1.5 5.5e-08 
1.0 1.12 0 -1.5 5.5e-08 
1.0 1.14 0 -1.5 5.5e-08 
1.0 1.16 0 -1.5 5.5e-08 
1.0 1.18 0 -1.5 5.5e-08 
1.0 1.2 0 -1.5 5.5e-08 
1.0 1.22 0 -1.5 5.5e-08 
1.0 1.24 0 -1.5 5.5e-08 
1.0 1.26 0 -1.5 5.5e-08 
1.0 1.28 0 -1.5 5.5e-08 
1.0 1.3 0 -1.5 5.5e-08 
1.0 1.32 0 -1.5 5.5e-08 
1.0 1.34 0 -1.5 5.5e-08 
1.0 1.36 0 -1.5 5.5e-08 
1.0 1.38 0 -1.5 5.5e-08 
1.0 1.4 0 -1.5 5.5e-08 
1.0 1.42 0 -1.5 5.5e-08 
1.0 1.44 0 -1.5 5.5e-08 
1.0 1.46 0 -1.5 5.5e-08 
1.0 1.48 0 -1.5 5.5e-08 
1.0 -1.5 0 -2.0 5.5e-08 
1.0 -1.48 0 -2.0 5.5e-08 
1.0 -1.46 0 -2.0 5.5e-08 
1.0 -1.44 0 -2.0 5.5e-08 
1.0 -1.42 0 -2.0 5.5e-08 
1.0 -1.4 0 -2.0 5.5e-08 
1.0 -1.38 0 -2.0 5.5e-08 
1.0 -1.36 0 -2.0 5.5e-08 
1.0 -1.34 0 -2.0 5.5e-08 
1.0 -1.32 0 -2.0 5.5e-08 
1.0 -1.3 0 -2.0 5.5e-08 
1.0 -1.28 0 -2.0 5.5e-08 
1.0 -1.26 0 -2.0 5.5e-08 
1.0 -1.24 0 -2.0 5.5e-08 
1.0 -1.22 0 -2.0 5.5e-08 
1.0 -1.2 0 -2.0 5.5e-08 
1.0 -1.18 0 -2.0 5.5e-08 
1.0 -1.16 0 -2.0 5.5e-08 
1.0 -1.14 0 -2.0 5.5e-08 
1.0 -1.12 0 -2.0 5.5e-08 
1.0 -1.1 0 -2.0 5.5e-08 
1.0 -1.08 0 -2.0 5.5e-08 
1.0 -1.06 0 -2.0 5.5e-08 
1.0 -1.04 0 -2.0 5.5e-08 
1.0 -1.02 0 -2.0 5.5e-08 
1.0 -1.0 0 -2.0 5.5e-08 
1.0 -0.98 0 -2.0 5.5e-08 
1.0 -0.96 0 -2.0 5.5e-08 
1.0 -0.94 0 -2.0 5.5e-08 
1.0 -0.92 0 -2.0 5.5e-08 
1.0 -0.9 0 -2.0 5.5e-08 
1.0 -0.88 0 -2.0 5.5e-08 
1.0 -0.86 0 -2.0 5.5e-08 
1.0 -0.84 0 -2.0 5.5e-08 
1.0 -0.82 0 -2.0 5.5e-08 
1.0 -0.8 0 -2.0 5.5e-08 
1.0 -0.78 0 -2.0 5.5e-08 
1.0 -0.76 0 -2.0 5.5e-08 
1.0 -0.74 0 -2.0 5.5e-08 
1.0 -0.72 0 -2.0 5.5e-08 
1.0 -0.7 0 -2.0 5.5e-08 
1.0 -0.68 0 -2.0 5.5e-08 
1.0 -0.66 0 -2.0 5.5e-08 
1.0 -0.64 0 -2.0 5.5e-08 
1.0 -0.62 0 -2.0 5.5e-08 
1.0 -0.6 0 -2.0 5.5e-08 
1.0 -0.58 0 -2.0 5.5e-08 
1.0 -0.56 0 -2.0 5.5e-08 
1.0 -0.54 0 -2.0 5.5e-08 
1.0 -0.52 0 -2.0 5.5e-08 
1.0 -0.5 0 -2.0 5.5e-08 
1.0 -0.48 0 -2.0 5.5e-08 
1.0 -0.46 0 -2.0 5.5e-08 
1.0 -0.44 0 -2.0 5.5e-08 
1.0 -0.42 0 -2.0 5.5e-08 
1.0 -0.4 0 -2.0 5.5e-08 
1.0 -0.38 0 -2.0 5.5e-08 
1.0 -0.36 0 -2.0 5.5e-08 
1.0 -0.34 0 -2.0 5.5e-08 
1.0 -0.32 0 -2.0 5.5e-08 
1.0 -0.3 0 -2.0 5.5e-08 
1.0 -0.28 0 -2.0 5.5e-08 
1.0 -0.26 0 -2.0 5.5e-08 
1.0 -0.24 0 -2.0 5.5e-08 
1.0 -0.22 0 -2.0 5.5e-08 
1.0 -0.2 0 -2.0 5.5e-08 
1.0 -0.18 0 -2.0 5.5e-08 
1.0 -0.16 0 -2.0 5.5e-08 
1.0 -0.14 0 -2.0 5.5e-08 
1.0 -0.12 0 -2.0 5.5e-08 
1.0 -0.1 0 -2.0 5.5e-08 
1.0 -0.08 0 -2.0 5.5e-08 
1.0 -0.06 0 -2.0 5.5e-08 
1.0 -0.04 0 -2.0 5.5e-08 
1.0 -0.02 0 -2.0 5.5e-08 
1.0 1.33226762955e-15 0 -2.0 5.5e-08 
1.0 0.02 0 -2.0 5.5e-08 
1.0 0.04 0 -2.0 5.5e-08 
1.0 0.06 0 -2.0 5.5e-08 
1.0 0.08 0 -2.0 5.5e-08 
1.0 0.1 0 -2.0 5.5e-08 
1.0 0.12 0 -2.0 5.5e-08 
1.0 0.14 0 -2.0 5.5e-08 
1.0 0.16 0 -2.0 5.5e-08 
1.0 0.18 0 -2.0 5.5e-08 
1.0 0.2 0 -2.0 5.5e-08 
1.0 0.22 0 -2.0 5.5e-08 
1.0 0.24 0 -2.0 5.5e-08 
1.0 0.26 0 -2.0 5.5e-08 
1.0 0.28 0 -2.0 5.5e-08 
1.0 0.3 0 -2.0 5.5e-08 
1.0 0.32 0 -2.0 5.5e-08 
1.0 0.34 0 -2.0 5.5e-08 
1.0 0.36 0 -2.0 5.5e-08 
1.0 0.38 0 -2.0 5.5e-08 
1.0 0.4 0 -2.0 5.5e-08 
1.0 0.42 0 -2.0 5.5e-08 
1.0 0.44 0 -2.0 5.5e-08 
1.0 0.46 0 -2.0 5.5e-08 
1.0 0.48 0 -2.0 5.5e-08 
1.0 0.5 0 -2.0 5.5e-08 
1.0 0.52 0 -2.0 5.5e-08 
1.0 0.54 0 -2.0 5.5e-08 
1.0 0.56 0 -2.0 5.5e-08 
1.0 0.58 0 -2.0 5.5e-08 
1.0 0.6 0 -2.0 5.5e-08 
1.0 0.62 0 -2.0 5.5e-08 
1.0 0.64 0 -2.0 5.5e-08 
1.0 0.66 0 -2.0 5.5e-08 
1.0 0.68 0 -2.0 5.5e-08 
1.0 0.7 0 -2.0 5.5e-08 
1.0 0.72 0 -2.0 5.5e-08 
1.0 0.74 0 -2.0 5.5e-08 
1.0 0.76 0 -2.0 5.5e-08 
1.0 0.78 0 -2.0 5.5e-08 
1.0 0.8 0 -2.0 5.5e-08 
1.0 0.82 0 -2.0 5.5e-08 
1.0 0.84 0 -2.0 5.5e-08 
1.0 0.86 0 -2.0 5.5e-08 
1.0 0.88 0 -2.0 5.5e-08 
1.0 0.9 0 -2.0 5.5e-08 
1.0 0.92 0 -2.0 5.5e-08 
1.0 0.94 0 -2.0 5.5e-08 
1.0 0.96 0 -2.0 5.5e-08 
1.0 0.98 0 -2.0 5.5e-08 
1.0 1.0 0 -2.0 5.5e-08 
1.0 1.02 0 -2.0 5.5e-08 
1.0 1.04 0 -2.0 5.5e-08 
1.0 1.06 0 -2.0 5.5e-08 
1.0 1.08 0 -2.0 5.5e-08 
1.0 1.1 0 -2.0 5.5e-08 
1.0 1.12 0 -2.0 5.5e-08 
1.0 1.14 0 -2.0 5.5e-08 
1.0 1.16 0 -2.0 5.5e-08 
1.0 1.18 0 -2.0 5.5e-08 
1.0 1.2 0 -2.0 5.5e-08 
1.0 1.22 0 -2.0 5.5e-08 
1.0 1.24 0 -2.0 5.5e-08 
1.0 1.26 0 -2.0 5.5e-08 
1.0 1.28 0 -2.0 5.5e-08 
1.0 1.3 0 -2.0 5.5e-08 
1.0 1.32 0 -2.0 5.5e-08 
1.0 1.34 0 -2.0 5.5e-08 
1.0 1.36 0 -2.0 5.5e-08 
1.0 1.38 0 -2.0 5.5e-08 
1.0 1.4 0 -2.0 5.5e-08 
1.0 1.42 0 -2.0 5.5e-08 
1.0 1.44 0 -2.0 5.5e-08 
1.0 1.46 0 -2.0 5.5e-08 
1.0 1.48 0 -2.0 5.5e-08 
1.0 -1.5 0 -2.5 5.5e-08 
1.0 -1.48 0 -2.5 5.5e-08 
1.0 -1.46 0 -2.5 5.5e-08 
1.0 -1.44 0 -2.5 5.5e-08 
1.0 -1.42 0 -2.5 5.5e-08 
1.0 -1.4 0 -2.5 5.5e-08 
1.0 -1.38 0 -2.5 5.5e-08 
1.0 -1.36 0 -2.5 5.5e-08 
1.0 -1.34 0 -2.5 5.5e-08 
1.0 -1.32 0 -2.5 5.5e-08 
1.0 -1.3 0 -2.5 5.5e-08 
1.0 -1.28 0 -2.5 5.5e-08 
1.0 -1.26 0 -2.5 5.5e-08 
1.0 -1.24 0 -2.5 5.5e-08 
1.0 -1.22 0 -2.5 5.5e-08 
1.0 -1.2 0 -2.5 5.5e-08 
1.0 -1.18 0 -2.5 5.5e-08 
1.0 -1.16 0 -2.5 5.5e-08 
1.0 -1.14 0 -2.5 5.5e-08 
1.0 -1.12 0 -2.5 5.5e-08 
1.0 -1.1 0 -2.5 5.5e-08 
1.0 -1.08 0 -2.5 5.5e-08 
1.0 -1.06 0 -2.5 5.5e-08 
1.0 -1.04 0 -2.5 5.5e-08 
1.0 -1.02 0 -2.5 5.5e-08 
1.0 -1.0 0 -2.5 5.5e-08 
1.0 -0.98 0 -2.5 5.5e-08 
1.0 -0.96 0 -2.5 5.5e-08 
1.0 -0.94 0 -2.5 5.5e-08 
1.0 -0.92 0 -2.5 5.5e-08 
1.0 -0.9 0 -2.5 5.5e-08 
1.0 -0.88 0 -2.5 5.5e-08 
1.0 -0.86 0 -2.5 5.5e-08 
1.0 -0.84 0 -2.5 5.5e-08 
1.0 -0.82 0 -2.5 5.5e-08 
1.0 -0.8 0 -2.5 5.5e-08 
1.0 -0.78 0 -2.5 5.5e-08 
1.0 -0.76 0 -2.5 5.5e-08 
1.0 -0.74 0 -2.5 5.5e-08 
1.0 -0.72 0 -2.5 5.5e-08 
1.0 -0.7 0 -2.5 5.5e-08 
1.0 -0.68 0 -2.5 5.5e-08 
1.0 -0.66 0 -2.5 5.5e-08 
1.0 -0.64 0 -2.5 5.5e-08 
1.0 -0.62 0 -2.5 5.5e-08 
1.0 -0.6 0 -2.5 5.5e-08 
1.0 -0.58 0 -2.5 5.5e-08 
1.0 -0.56 0 -2.5 5.5e-08 
1.0 -0.54 0 -2.5 5.5e-08 
1.0 -0.52 0 -2.5 5.5e-08 
1.0 -0.5 0 -2.5 5.5e-08 
1.0 -0.48 0 -2.5 5.5e-08 
1.0 -0.46 0 -2.5 5.5e-08 
1.0 -0.44 0 -2.5 5.5e-08 
1.0 -0.42 0 -2.5 5.5e-08 
1.0 -0.4 0 -2.5 5.5e-08 
1.0 -0.38 0 -2.5 5.5e-08 
1.0 -0.36 0 -2.5 5.5e-08 
1.0 -0.34 0 -2.5 5.5e-08 
1.0 -0.32 0 -2.5 5.5e-08 
1.0 -0.3 0 -2.5 5.5e-08 
1.0 -0.28 0 -2.5 5.5e-08 
1.0 -0.26 0 -2.5 5.5e-08 
1.0 -0.24 0 -2.5 5.5e-08 
1.0 -0.22 0 -2.5 5.5e-08 
1.0 -0.2 0 -2.5 5.5e-08 
1.0 -0.18 0 -2.5 5.5e-08 
1.0 -0.16 0 -2.5 5.5e-08 
1.0 -0.14 0 -2.5 5.5e-08 
1.0 -0.12 0 -2.5 5.5e-08 
1.0 -0.1 0 -2.5 5.5e-08 
1.0 -0.08 0 -2.5 5.5e-08 
1.0 -0.06 0 -2.5 5.5e-08 
1.0 -0.04 0 -2.5 5.5e-08 
1.0 -0.02 0 -2.5 5.5e-08 
1.0 1.33226762955e-15 0 -2.5 5.5e-08 
1.0 0.02 0 -2.5 5.5e-08 
1.0 0.04 0 -2.5 5.5e-08 
1.0 0.06 0 -2.5 5.5e-08 
1.0 0.08 0 -2.5 5.5e-08 
1.0 0.1 0 -2.5 5.5e-08 
1.0 0.12 0 -2.5 5.5e-08 
1.0 0.14 0 -2.5 5.5e-08 
1.0 0.16 0 -2.5 5.5e-08 
1.0 0.18 0 -2.5 5.5e-08 
1.0 0.2 0 -2.5 5.5e-08 
1.0 0.22 0 -2.5 5.5e-08 
1.0 0.24 0 -2.5 5.5e-08 
1.0 0.26 0 -2.5 5.5e-08 
1.0 0.28 0 -2.5 5.5e-08 
1.0 0.3 0 -2.5 5.5e-08 
1.0 0.32 0 -2.5 5.5e-08 
1.0 0.34 0 -2.5 5.5e-08 
1.0 0.36 0 -2.5 5.5e-08 
1.0 0.38 0 -2.5 5.5e-08 
1.0 0.4 0 -2.5 5.5e-08 
1.0 0.42 0 -2.5 5.5e-08 
1.0 0.44 0 -2.5 5.5e-08 
1.0 0.46 0 -2.5 5.5e-08 
1.0 0.48 0 -2.5 5.5e-08 
1.0 0.5 0 -2.5 5.5e-08 
1.0 0.52 0 -2.5 5.5e-08 
1.0 0.54 0 -2.5 5.5e-08 
1.0 0.56 0 -2.5 5.5e-08 
1.0 0.58 0 -2.5 5.5e-08 
1.0 0.6 0 -2.5 5.5e-08 
1.0 0.62 0 -2.5 5.5e-08 
1.0 0.64 0 -2.5 5.5e-08 
1.0 0.66 0 -2.5 5.5e-08 
1.0 0.68 0 -2.5 5.5e-08 
1.0 0.7 0 -2.5 5.5e-08 
1.0 0.72 0 -2.5 5.5e-08 
1.0 0.74 0 -2.5 5.5e-08 
1.0 0.76 0 -2.5 5.5e-08 
1.0 0.78 0 -2.5 5.5e-08 
1.0 0.8 0 -2.5 5.5e-08 
1.0 0.82 0 -2.5 5.5e-08 
1.0 0.84 0 -2.5 5.5e-08 
1.0 0.86 0 -2.5 5.5e-08 
1.0 0.88 0 -2.5 5.5e-08 
1.0 0.9 0 -2.5 5.5e-08 
1.0 0.92 0 -2.5 5.5e-08 
1.0 0.94 0 -2.5 5.5e-08 
1.0 0.96 0 -2.5 5.5e-08 
1.0 0.98 0 -2.5 5.5e-08 
1.0 1.0 0 -2.5 5.5e-08 
1.0 1.02 0 -2.5 5.5e-08 
1.0 1.04 0 -2.5 5.5e-08 
1.0 1.06 0 -2.5 5.5e-08 
1.0 1.08 0 -2.5 5.5e-08 
1.0 1.1 0 -2.5 5.5e-08 
1.0 1.12 0 -2.5 5.5e-08 
1.0 1.14 0 -2.5 5.5e-08 
1.0 1.16 0 -2.5 5.5e-08 
1.0 1.18 0 -2.5 5.5e-08 
1.0 1.2 0 -2.5 5.5e-08 
1.0 1.22 0 -2.5 5.5e-08 
1.0 1.24 0 -2.5 5.5e-08 
1.0 1.26 0 -2.5 5.5e-08 
1.0 1.28 0 -2.5 5.5e-08 
1.0 1.3 0 -2.5 5.5e-08 
1.0 1.32 0 -2.5 5.5e-08 
1.0 1.34 0 -2.5 5.5e-08 
1.0 1.36 0 -2.5 5.5e-08 
1.0 1.38 0 -2.5 5.5e-08 
1.0 1.4 0 -2.5 5.5e-08 
1.0 1.42 0 -2.5 5.5e-08 
1.0 1.44 0 -2.5 5.5e-08 
1.0 1.46 0 -2.5 5.5e-08 
1.0 1.48 0 -2.5 5.5e-08 
1.0 -1.5 0 -3.0 5.5e-08 
1.0 -1.48 0 -3.0 5.5e-08 
1.0 -1.46 0 -3.0 5.5e-08 
1.0 -1.44 0 -3.0 5.5e-08 
1.0 -1.42 0 -3.0 5.5e-08 
1.0 -1.4 0 -3.0 5.5e-08 
1.0 -1.38 0 -3.0 5.5e-08 
1.0 -1.36 0 -3.0 5.5e-08 
1.0 -1.34 0 -3.0 5.5e-08 
1.0 -1.32 0 -3.0 5.5e-08 
1.0 -1.3 0 -3.0 5.5e-08 
1.0 -1.28 0 -3.0 5.5e-08 
1.0 -1.26 0 -3.0 5.5e-08 
1.0 -1.24 0 -3.0 5.5e-08 
1.0 -1.22 0 -3.0 5.5e-08 
1.0 -1.2 0 -3.0 5.5e-08 
1.0 -1.18 0 -3.0 5.5e-08 
1.0 -1.16 0 -3.0 5.5e-08 
1.0 -1.14 0 -3.0 5.5e-08 
1.0 -1.12 0 -3.0 5.5e-08 
1.0 -1.1 0 -3.0 5.5e-08 
1.0 -1.08 0 -3.0 5.5e-08 
1.0 -1.06 0 -3.0 5.5e-08 
1.0 -1.04 0 -3.0 5.5e-08 
1.0 -1.02 0 -3.0 5.5e-08 
1.0 -1.0 0 -3.0 5.5e-08 
1.0 -0.98 0 -3.0 5.5e-08 
1.0 -0.96 0 -3.0 5.5e-08 
1.0 -0.94 0 -3.0 5.5e-08 
1.0 -0.92 0 -3.0 5.5e-08 
1.0 -0.9 0 -3.0 5.5e-08 
1.0 -0.88 0 -3.0 5.5e-08 
1.0 -0.86 0 -3.0 5.5e-08 
1.0 -0.84 0 -3.0 5.5e-08 
1.0 -0.82 0 -3.0 5.5e-08 
1.0 -0.8 0 -3.0 5.5e-08 
1.0 -0.78 0 -3.0 5.5e-08 
1.0 -0.76 0 -3.0 5.5e-08 
1.0 -0.74 0 -3.0 5.5e-08 
1.0 -0.72 0 -3.0 5.5e-08 
1.0 -0.7 0 -3.0 5.5e-08 
1.0 -0.68 0 -3.0 5.5e-08 
1.0 -0.66 0 -3.0 5.5e-08 
1.0 -0.64 0 -3.0 5.5e-08 
1.0 -0.62 0 -3.0 5.5e-08 
1.0 -0.6 0 -3.0 5.5e-08 
1.0 -0.58 0 -3.0 5.5e-08 
1.0 -0.56 0 -3.0 5.5e-08 
1.0 -0.54 0 -3.0 5.5e-08 
1.0 -0.52 0 -3.0 5.5e-08 
1.0 -0.5 0 -3.0 5.5e-08 
1.0 -0.48 0 -3.0 5.5e-08 
1.0 -0.46 0 -3.0 5.5e-08 
1.0 -0.44 0 -3.0 5.5e-08 
1.0 -0.42 0 -3.0 5.5e-08 
1.0 -0.4 0 -3.0 5.5e-08 
1.0 -0.38 0 -3.0 5.5e-08 
1.0 -0.36 0 -3.0 5.5e-08 
1.0 -0.34 0 -3.0 5.5e-08 
1.0 -0.32 0 -3.0 5.5e-08 
1.0 -0.3 0 -3.0 5.5e-08 
1.0 -0.28 0 -3.0 5.5e-08 
1.0 -0.26 0 -3.0 5.5e-08 
1.0 -0.24 0 -3.0 5.5e-08 
1.0 -0.22 0 -3.0 5.5e-08 
1.0 -0.2 0 -3.0 5.5e-08 
1.0 -0.18 0 -3.0 5.5e-08 
1.0 -0.16 0 -3.0 5.5e-08 
1.0 -0.14 0 -3.0 5.5e-08 
1.0 -0.12 0 -3.0 5.5e-08 
1.0 -0.1 0 -3.0 5.5e-08 
1.0 -0.08 0 -3.0 5.5e-08 
1.0 -0.06 0 -3.0 5.5e-08 
1.0 -0.04 0 -3.0 5.5e-08 
1.0 -0.02 0 -3.0 5.5e-08 
1.0 1.33226762955e-15 0 -3.0 5.5e-08 
1.0 0.02 0 -3.0 5.5e-08 
1.0 0.04 0 -3.0 5.5e-08 
1.0 0.06 0 -3.0 5.5e-08 
1.0 0.08 0 -3.0 5.5e-08 
1.0 0.1 0 -3.0 5.5e-08 
1.0 0.12 0 -3.0 5.5e-08 
1.0 0.14 0 -3.0 5.5e-08 
1.0 0.16 0 -3.0 5.5e-08 
1.0 0.18 0 -3.0 5.5e-08 
1.0 0.2 0 -3.0 5.5e-08 
1.0 0.22 0 -3.0 5.5e-08 
1.0 0.24 0 -3.0 5.5e-08 
1.0 0.26 0 -3.0 5.5e-08 
1.0 0.28 0 -3.0 5.5e-08 
1.0 0.3 0 -3.0 5.5e-08 
1.0 0.32 0 -3.0 5.5e-08 
1.0 0.34 0 -3.0 5.5e-08 
1.0 0.36 0 -3.0 5.5e-08 
1.0 0.38 0 -3.0 5.5e-08 
1.0 0.4 0 -3.0 5.5e-08 
1.0 0.42 0 -3.0 5.5e-08 
1.0 0.44 0 -3.0 5.5e-08 
1.0 0.46 0 -3.0 5.5e-08 
1.0 0.48 0 -3.0 5.5e-08 
1.0 0.5 0 -3.0 5.5e-08 
1.0 0.52 0 -3.0 5.5e-08 
1.0 0.54 0 -3.0 5.5e-08 
1.0 0.56 0 -3.0 5.5e-08 
1.0 0.58 0 -3.0 5.5e-08 
1.0 0.6 0 -3.0 5.5e-08 
1.0 0.62 0 -3.0 5.5e-08 
1.0 0.64 0 -3.0 5.5e-08 
1.0 0.66 0 -3.0 5.5e-08 
1.0 0.68 0 -3.0 5.5e-08 
1.0 0.7 0 -3.0 5.5e-08 
1.0 0.72 0 -3.0 5.5e-08 
1.0 0.74 0 -3.0 5.5e-08 
1.0 0.76 0 -3.0 5.5e-08 
1.0 0.78 0 -3.0 5.5e-08 
1.0 0.8 0 -3.0 5.5e-08 
1.0 0.82 0 -3.0 5.5e-08 
1.0 0.84 0 -3.0 5.5e-08 
1.0 0.86 0 -3.0 5.5e-08 
1.0 0.88 0 -3.0 5.5e-08 
1.0 0.9 0 -3.0 5.5e-08 
1.0 0.92 0 -3.0 5.5e-08 
1.0 0.94 0 -3.0 5.5e-08 
1.0 0.96 0 -3.0 5.5e-08 
1.0 0.98 0 -3.0 5.5e-08 
1.0 1.0 0 -3.0 5.5e-08 
1.0 1.02 0 -3.0 5.5e-08 
1.0 1.04 0 -3.0 5.5e-08 
1.0 1.06 0 -3.0 5.5e-08 
1.0 1.08 0 -3.0 5.5e-08 
1.0 1.1 0 -3.0 5.5e-08 
1.0 1.12 0 -3.0 5.5e-08 
1.0 1.14 0 -3.0 5.5e-08 
1.0 1.16 0 -3.0 5.5e-08 
1.0 1.18 0 -3.0 5.5e-08 
1.0 1.2 0 -3.0 5.5e-08 
1.0 1.22 0 -3.0 5.5e-08 
1.0 1.24 0 -3.0 5.5e-08 
1.0 1.26 0 -3.0 5.5e-08 
1.0 1.28 0 -3.0 5.5e-08 
1.0 1.3 0 -3.0 5.5e-08 
1.0 1.32 0 -3.0 5.5e-08 
1.0 1.34 0 -3.0 5.5e-08 
1.0 1.36 0 -3.0 5.5e-08 
1.0 1.38 0 -3.0 5.5e-08 
1.0 1.4 0 -3.0 5.5e-08 
1.0 1.42 0 -3.0 5.5e-08 
1.0 1.44 0 -3.0 5.5e-08 
1.0 1.46 0 -3.0 5.5e-08 
1.0 1.48 0 -3.0 5.5e-08 
1.0 -1.5 0 -3.5 5.5e-08 
1.0 -1.48 0 -3.5 5.5e-08 
1.0 -1.46 0 -3.5 5.5e-08 
1.0 -1.44 0 -3.5 5.5e-08 
1.0 -1.42 0 -3.5 5.5e-08 
1.0 -1.4 0 -3.5 5.5e-08 
1.0 -1.38 0 -3.5 5.5e-08 
1.0 -1.36 0 -3.5 5.5e-08 
1.0 -1.34 0 -3.5 5.5e-08 
1.0 -1.32 0 -3.5 5.5e-08 
1.0 -1.3 0 -3.5 5.5e-08 
1.0 -1.28 0 -3.5 5.5e-08 
1.0 -1.26 0 -3.5 5.5e-08 
1.0 -1.24 0 -3.5 5.5e-08 
1.0 -1.22 0 -3.5 5.5e-08 
1.0 -1.2 0 -3.5 5.5e-08 
1.0 -1.18 0 -3.5 5.5e-08 
1.0 -1.16 0 -3.5 5.5e-08 
1.0 -1.14 0 -3.5 5.5e-08 
1.0 -1.12 0 -3.5 5.5e-08 
1.0 -1.1 0 -3.5 5.5e-08 
1.0 -1.08 0 -3.5 5.5e-08 
1.0 -1.06 0 -3.5 5.5e-08 
1.0 -1.04 0 -3.5 5.5e-08 
1.0 -1.02 0 -3.5 5.5e-08 
1.0 -1.0 0 -3.5 5.5e-08 
1.0 -0.98 0 -3.5 5.5e-08 
1.0 -0.96 0 -3.5 5.5e-08 
1.0 -0.94 0 -3.5 5.5e-08 
1.0 -0.92 0 -3.5 5.5e-08 
1.0 -0.9 0 -3.5 5.5e-08 
1.0 -0.88 0 -3.5 5.5e-08 
1.0 -0.86 0 -3.5 5.5e-08 
1.0 -0.84 0 -3.5 5.5e-08 
1.0 -0.82 0 -3.5 5.5e-08 
1.0 -0.8 0 -3.5 5.5e-08 
1.0 -0.78 0 -3.5 5.5e-08 
1.0 -0.76 0 -3.5 5.5e-08 
1.0 -0.74 0 -3.5 5.5e-08 
1.0 -0.72 0 -3.5 5.5e-08 
1.0 -0.7 0 -3.5 5.5e-08 
1.0 -0.68 0 -3.5 5.5e-08 
1.0 -0.66 0 -3.5 5.5e-08 
1.0 -0.64 0 -3.5 5.5e-08 
1.0 -0.62 0 -3.5 5.5e-08 
1.0 -0.6 0 -3.5 5.5e-08 
1.0 -0.58 0 -3.5 5.5e-08 
1.0 -0.56 0 -3.5 5.5e-08 
1.0 -0.54 0 -3.5 5.5e-08 
1.0 -0.52 0 -3.5 5.5e-08 
1.0 -0.5 0 -3.5 5.5e-08 
1.0 -0.48 0 -3.5 5.5e-08 
1.0 -0.46 0 -3.5 5.5e-08 
1.0 -0.44 0 -3.5 5.5e-08 
1.0 -0.42 0 -3.5 5.5e-08 
1.0 -0.4 0 -3.5 5.5e-08 
1.0 -0.38 0 -3.5 5.5e-08 
1.0 -0.36 0 -3.5 5.5e-08 
1.0 -0.34 0 -3.5 5.5e-08 
1.0 -0.32 0 -3.5 5.5e-08 
1.0 -0.3 0 -3.5 5.5e-08 
1.0 -0.28 0 -3.5 5.5e-08 
1.0 -0.26 0 -3.5 5.5e-08 
1.0 -0.24 0 -3.5 5.5e-08 
1.0 -0.22 0 -3.5 5.5e-08 
1.0 -0.2 0 -3.5 5.5e-08 
1.0 -0.18 0 -3.5 5.5e-08 
1.0 -0.16 0 -3.5 5.5e-08 
1.0 -0.14 0 -3.5 5.5e-08 
1.0 -0.12 0 -3.5 5.5e-08 
1.0 -0.1 0 -3.5 5.5e-08 
1.0 -0.08 0 -3.5 5.5e-08 
1.0 -0.06 0 -3.5 5.5e-08 
1.0 -0.04 0 -3.5 5.5e-08 
1.0 -0.02 0 -3.5 5.5e-08 
1.0 1.33226762955e-15 0 -3.5 5.5e-08 
1.0 0.02 0 -3.5 5.5e-08 
1.0 0.04 0 -3.5 5.5e-08 
1.0 0.06 0 -3.5 5.5e-08 
1.0 0.08 0 -3.5 5.5e-08 
1.0 0.1 0 -3.5 5.5e-08 
1.0 0.12 0 -3.5 5.5e-08 
1.0 0.14 0 -3.5 5.5e-08 
1.0 0.16 0 -3.5 5.5e-08 
1.0 0.18 0 -3.5 5.5e-08 
1.0 0.2 0 -3.5 5.5e-08 
1.0 0.22 0 -3.5 5.5e-08 
1.0 0.24 0 -3.5 5.5e-08 
1.0 0.26 0 -3.5 5.5e-08 
1.0 0.28 0 -3.5 5.5e-08 
1.0 0.3 0 -3.5 5.5e-08 
1.0 0.32 0 -3.5 5.5e-08 
1.0 0.34 0 -3.5 5.5e-08 
1.0 0.36 0 -3.5 5.5e-08 
1.0 0.38 0 -3.5 5.5e-08 
1.0 0.4 0 -3.5 5.5e-08 
1.0 0.42 0 -3.5 5.5e-08 
1.0 0.44 0 -3.5 5.5e-08 
1.0 0.46 0 -3.5 5.5e-08 
1.0 0.48 0 -3.5 5.5e-08 
1.0 0.5 0 -3.5 5.5e-08 
1.0 0.52 0 -3.5 5.5e-08 
1.0 0.54 0 -3.5 5.5e-08 
1.0 0.56 0 -3.5 5.5e-08 
1.0 0.58 0 -3.5 5.5e-08 
1.0 0.6 0 -3.5 5.5e-08 
1.0 0.62 0 -3.5 5.5e-08 
1.0 0.64 0 -3.5 5.5e-08 
1.0 0.66 0 -3.5 5.5e-08 
1.0 0.68 0 -3.5 5.5e-08 
1.0 0.7 0 -3.5 5.5e-08 
1.0 0.72 0 -3.5 5.5e-08 
1.0 0.74 0 -3.5 5.5e-08 
1.0 0.76 0 -3.5 5.5e-08 
1.0 0.78 0 -3.5 5.5e-08 
1.0 0.8 0 -3.5 5.5e-08 
1.0 0.82 0 -3.5 5.5e-08 
1.0 0.84 0 -3.5 5.5e-08 
1.0 0.86 0 -3.5 5.5e-08 
1.0 0.88 0 -3.5 5.5e-08 
1.0 0.9 0 -3.5 5.5e-08 
1.0 0.92 0 -3.5 5.5e-08 
1.0 0.94 0 -3.5 5.5e-08 
1.0 0.96 0 -3.5 5.5e-08 
1.0 0.98 0 -3.5 5.5e-08 
1.0 1.0 0 -3.5 5.5e-08 
1.0 1.02 0 -3.5 5.5e-08 
1.0 1.04 0 -3.5 5.5e-08 
1.0 1.06 0 -3.5 5.5e-08 
1.0 1.08 0 -3.5 5.5e-08 
1.0 1.1 0 -3.5 5.5e-08 
1.0 1.12 0 -3.5 5.5e-08 
1.0 1.14 0 -3.5 5.5e-08 
1.0 1.16 0 -3.5 5.5e-08 
1.0 1.18 0 -3.5 5.5e-08 
1.0 1.2 0 -3.5 5.5e-08 
1.0 1.22 0 -3.5 5.5e-08 
1.0 1.24 0 -3.5 5.5e-08 
1.0 1.26 0 -3.5 5.5e-08 
1.0 1.28 0 -3.5 5.5e-08 
1.0 1.3 0 -3.5 5.5e-08 
1.0 1.32 0 -3.5 5.5e-08 
1.0 1.34 0 -3.5 5.5e-08 
1.0 1.36 0 -3.5 5.5e-08 
1.0 1.38 0 -3.5 5.5e-08 
1.0 1.4 0 -3.5 5.5e-08 
1.0 1.42 0 -3.5 5.5e-08 
1.0 1.44 0 -3.5 5.5e-08 
1.0 1.46 0 -3.5 5.5e-08 
1.0 1.48 0 -3.5 5.5e-08 
1.0 -1.5 0 -4.0 5.5e-08 
1.0 -1.48 0 -4.0 5.5e-08 
1.0 -1.46 0 -4.0 5.5e-08 
1.0 -1.44 0 -4.0 5.5e-08 
1.0 -1.42 0 -4.0 5.5e-08 
1.0 -1.4 0 -4.0 5.5e-08 
1.0 -1.38 0 -4.0 5.5e-08 
1.0 -1.36 0 -4.0 5.5e-08 
1.0 -1.34 0 -4.0 5.5e-08 
1.0 -1.32 0 -4.0 5.5e-08 
1.0 -1.3 0 -4.0 5.5e-08 
1.0 -1.28 0 -4.0 5.5e-08 
1.0 -1.26 0 -4.0 5.5e-08 
1.0 -1.24 0 -4.0 5.5e-08 
1.0 -1.22 0 -4.0 5.5e-08 
1.0 -1.2 0 -4.0 5.5e-08 
1.0 -1.18 0 -4.0 5.5e-08 
1.0 -1.16 0 -4.0 5.5e-08 
1.0 -1.14 0 -4.0 5.5e-08 
1.0 -1.12 0 -4.0 5.5e-08 
1.0 -1.1 0 -4.0 5.5e-08 
1.0 -1.08 0 -4.0 5.5e-08 
1.0 -1.06 0 -4.0 5.5e-08 
1.0 -1.04 0 -4.0 5.5e-08 
1.0 -1.02 0 -4.0 5.5e-08 
1.0 -1.0 0 -4.0 5.5e-08 
1.0 -0.98 0 -4.0 5.5e-08 
1.0 -0.96 0 -4.0 5.5e-08 
1.0 -0.94 0 -4.0 5.5e-08 
1.0 -0.92 0 -4.0 5.5e-08 
1.0 -0.9 0 -4.0 5.5e-08 
1.0 -0.88 0 -4.0 5.5e-08 
1.0 -0.86 0 -4.0 5.5e-08 
1.0 -0.84 0 -4.0 5.5e-08 
1.0 -0.82 0 -4.0 5.5e-08 
1.0 -0.8 0 -4.0 5.5e-08 
1.0 -0.78 0 -4.0 5.5e-08 
1.0 -0.76 0 -4.0 5.5e-08 
1.0 -0.74 0 -4.0 5.5e-08 
1.0 -0.72 0 -4.0 5.5e-08 
1.0 -0.7 0 -4.0 5.5e-08 
1.0 -0.68 0 -4.0 5.5e-08 
1.0 -0.66 0 -4.0 5.5e-08 
1.0 -0.64 0 -4.0 5.5e-08 
1.0 -0.62 0 -4.0 5.5e-08 
1.0 -0.6 0 -4.0 5.5e-08 
1.0 -0.58 0 -4.0 5.5e-08 
1.0 -0.56 0 -4.0 5.5e-08 
1.0 -0.54 0 -4.0 5.5e-08 
1.0 -0.52 0 -4.0 5.5e-08 
1.0 -0.5 0 -4.0 5.5e-08 
1.0 -0.48 0 -4.0 5.5e-08 
1.0 -0.46 0 -4.0 5.5e-08 
1.0 -0.44 0 -4.0 5.5e-08 
1.0 -0.42 0 -4.0 5.5e-08 
1.0 -0.4 0 -4.0 5.5e-08 
1.0 -0.38 0 -4.0 5.5e-08 
1.0 -0.36 0 -4.0 5.5e-08 
1.0 -0.34 0 -4.0 5.5e-08 
1.0 -0.32 0 -4.0 5.5e-08 
1.0 -0.3 0 -4.0 5.5e-08 
1.0 -0.28 0 -4.0 5.5e-08 
1.0 -0.26 0 -4.0 5.5e-08 
1.0 -0.24 0 -4.0 5.5e-08 
1.0 -0.22 0 -4.0 5.5e-08 
1.0 -0.2 0 -4.0 5.5e-08 
1.0 -0.18 0 -4.0 5.5e-08 
1.0 -0.16 0 -4.0 5.5e-08 
1.0 -0.14 0 -4.0 5.5e-08 
1.0 -0.12 0 -4.0 5.5e-08 
1.0 -0.1 0 -4.0 5.5e-08 
1.0 -0.08 0 -4.0 5.5e-08 
1.0 -0.06 0 -4.0 5.5e-08 
1.0 -0.04 0 -4.0 5.5e-08 
1.0 -0.02 0 -4.0 5.5e-08 
1.0 1.33226762955e-15 0 -4.0 5.5e-08 
1.0 0.02 0 -4.0 5.5e-08 
1.0 0.04 0 -4.0 5.5e-08 
1.0 0.06 0 -4.0 5.5e-08 
1.0 0.08 0 -4.0 5.5e-08 
1.0 0.1 0 -4.0 5.5e-08 
1.0 0.12 0 -4.0 5.5e-08 
1.0 0.14 0 -4.0 5.5e-08 
1.0 0.16 0 -4.0 5.5e-08 
1.0 0.18 0 -4.0 5.5e-08 
1.0 0.2 0 -4.0 5.5e-08 
1.0 0.22 0 -4.0 5.5e-08 
1.0 0.24 0 -4.0 5.5e-08 
1.0 0.26 0 -4.0 5.5e-08 
1.0 0.28 0 -4.0 5.5e-08 
1.0 0.3 0 -4.0 5.5e-08 
1.0 0.32 0 -4.0 5.5e-08 
1.0 0.34 0 -4.0 5.5e-08 
1.0 0.36 0 -4.0 5.5e-08 
1.0 0.38 0 -4.0 5.5e-08 
1.0 0.4 0 -4.0 5.5e-08 
1.0 0.42 0 -4.0 5.5e-08 
1.0 0.44 0 -4.0 5.5e-08 
1.0 0.46 0 -4.0 5.5e-08 
1.0 0.48 0 -4.0 5.5e-08 
1.0 0.5 0 -4.0 5.5e-08 
1.0 0.52 0 -4.0 5.5e-08 
1.0 0.54 0 -4.0 5.5e-08 
1.0 0.56 0 -4.0 5.5e-08 
1.0 0.58 0 -4.0 5.5e-08 
1.0 0.6 0 -4.0 5.5e-08 
1.0 0.62 0 -4.0 5.5e-08 
1.0 0.64 0 -4.0 5.5e-08 
1.0 0.66 0 -4.0 5.5e-08 
1.0 0.68 0 -4.0 5.5e-08 
1.0 0.7 0 -4.0 5.5e-08 
1.0 0.72 0 -4.0 5.5e-08 
1.0 0.74 0 -4.0 5.5e-08 
1.0 0.76 0 -4.0 5.5e-08 
1.0 0.78 0 -4.0 5.5e-08 
1.0 0.8 0 -4.0 5.5e-08 
1.0 0.82 0 -4.0 5.5e-08 
1.0 0.84 0 -4.0 5.5e-08 
1.0 0.86 0 -4.0 5.5e-08 
1.0 0.88 0 -4.0 5.5e-08 
1.0 0.9 0 -4.0 5.5e-08 
1.0 0.92 0 -4.0 5.5e-08 
1.0 0.94 0 -4.0 5.5e-08 
1.0 0.96 0 -4.0 5.5e-08 
1.0 0.98 0 -4.0 5.5e-08 
1.0 1.0 0 -4.0 5.5e-08 
1.0 1.02 0 -4.0 5.5e-08 
1.0 1.04 0 -4.0 5.5e-08 
1.0 1.06 0 -4.0 5.5e-08 
1.0 1.08 0 -4.0 5.5e-08 
1.0 1.1 0 -4.0 5.5e-08 
1.0 1.12 0 -4.0 5.5e-08 
1.0 1.14 0 -4.0 5.5e-08 
1.0 1.16 0 -4.0 5.5e-08 
1.0 1.18 0 -4.0 5.5e-08 
1.0 1.2 0 -4.0 5.5e-08 
1.0 1.22 0 -4.0 5.5e-08 
1.0 1.24 0 -4.0 5.5e-08 
1.0 1.26 0 -4.0 5.5e-08 
1.0 1.28 0 -4.0 5.5e-08 
1.0 1.3 0 -4.0 5.5e-08 
1.0 1.32 0 -4.0 5.5e-08 
1.0 1.34 0 -4.0 5.5e-08 
1.0 1.36 0 -4.0 5.5e-08 
1.0 1.38 0 -4.0 5.5e-08 
1.0 1.4 0 -4.0 5.5e-08 
1.0 1.42 0 -4.0 5.5e-08 
1.0 1.44 0 -4.0 5.5e-08 
1.0 1.46 0 -4.0 5.5e-08 
1.0 1.48 0 -4.0 5.5e-08 
1.0 -1.5 0 -4.5 5.5e-08 
1.0 -1.48 0 -4.5 5.5e-08 
1.0 -1.46 0 -4.5 5.5e-08 
1.0 -1.44 0 -4.5 5.5e-08 
1.0 -1.42 0 -4.5 5.5e-08 
1.0 -1.4 0 -4.5 5.5e-08 
1.0 -1.38 0 -4.5 5.5e-08 
1.0 -1.36 0 -4.5 5.5e-08 
1.0 -1.34 0 -4.5 5.5e-08 
1.0 -1.32 0 -4.5 5.5e-08 
1.0 -1.3 0 -4.5 5.5e-08 
1.0 -1.28 0 -4.5 5.5e-08 
1.0 -1.26 0 -4.5 5.5e-08 
1.0 -1.24 0 -4.5 5.5e-08 
1.0 -1.22 0 -4.5 5.5e-08 
1.0 -1.2 0 -4.5 5.5e-08 
1.0 -1.18 0 -4.5 5.5e-08 
1.0 -1.16 0 -4.5 5.5e-08 
1.0 -1.14 0 -4.5 5.5e-08 
1.0 -1.12 0 -4.5 5.5e-08 
1.0 -1.1 0 -4.5 5.5e-08 
1.0 -1.08 0 -4.5 5.5e-08 
1.0 -1.06 0 -4.5 5.5e-08 
1.0 -1.04 0 -4.5 5.5e-08 
1.0 -1.02 0 -4.5 5.5e-08 
1.0 -1.0 0 -4.5 5.5e-08 
1.0 -0.98 0 -4.5 5.5e-08 
1.0 -0.96 0 -4.5 5.5e-08 
1.0 -0.94 0 -4.5 5.5e-08 
1.0 -0.92 0 -4.5 5.5e-08 
1.0 -0.9 0 -4.5 5.5e-08 
1.0 -0.88 0 -4.5 5.5e-08 
1.0 -0.86 0 -4.5 5.5e-08 
1.0 -0.84 0 -4.5 5.5e-08 
1.0 -0.82 0 -4.5 5.5e-08 
1.0 -0.8 0 -4.5 5.5e-08 
1.0 -0.78 0 -4.5 5.5e-08 
1.0 -0.76 0 -4.5 5.5e-08 
1.0 -0.74 0 -4.5 5.5e-08 
1.0 -0.72 0 -4.5 5.5e-08 
1.0 -0.7 0 -4.5 5.5e-08 
1.0 -0.68 0 -4.5 5.5e-08 
1.0 -0.66 0 -4.5 5.5e-08 
1.0 -0.64 0 -4.5 5.5e-08 
1.0 -0.62 0 -4.5 5.5e-08 
1.0 -0.6 0 -4.5 5.5e-08 
1.0 -0.58 0 -4.5 5.5e-08 
1.0 -0.56 0 -4.5 5.5e-08 
1.0 -0.54 0 -4.5 5.5e-08 
1.0 -0.52 0 -4.5 5.5e-08 
1.0 -0.5 0 -4.5 5.5e-08 
1.0 -0.48 0 -4.5 5.5e-08 
1.0 -0.46 0 -4.5 5.5e-08 
1.0 -0.44 0 -4.5 5.5e-08 
1.0 -0.42 0 -4.5 5.5e-08 
1.0 -0.4 0 -4.5 5.5e-08 
1.0 -0.38 0 -4.5 5.5e-08 
1.0 -0.36 0 -4.5 5.5e-08 
1.0 -0.34 0 -4.5 5.5e-08 
1.0 -0.32 0 -4.5 5.5e-08 
1.0 -0.3 0 -4.5 5.5e-08 
1.0 -0.28 0 -4.5 5.5e-08 
1.0 -0.26 0 -4.5 5.5e-08 
1.0 -0.24 0 -4.5 5.5e-08 
1.0 -0.22 0 -4.5 5.5e-08 
1.0 -0.2 0 -4.5 5.5e-08 
1.0 -0.18 0 -4.5 5.5e-08 
1.0 -0.16 0 -4.5 5.5e-08 
1.0 -0.14 0 -4.5 5.5e-08 
1.0 -0.12 0 -4.5 5.5e-08 
1.0 -0.1 0 -4.5 5.5e-08 
1.0 -0.08 0 -4.5 5.5e-08 
1.0 -0.06 0 -4.5 5.5e-08 
1.0 -0.04 0 -4.5 5.5e-08 
1.0 -0.02 0 -4.5 5.5e-08 
1.0 1.33226762955e-15 0 -4.5 5.5e-08 
1.0 0.02 0 -4.5 5.5e-08 
1.0 0.04 0 -4.5 5.5e-08 
1.0 0.06 0 -4.5 5.5e-08 
1.0 0.08 0 -4.5 5.5e-08 
1.0 0.1 0 -4.5 5.5e-08 
1.0 0.12 0 -4.5 5.5e-08 
1.0 0.14 0 -4.5 5.5e-08 
1.0 0.16 0 -4.5 5.5e-08 
1.0 0.18 0 -4.5 5.5e-08 
1.0 0.2 0 -4.5 5.5e-08 
1.0 0.22 0 -4.5 5.5e-08 
1.0 0.24 0 -4.5 5.5e-08 
1.0 0.26 0 -4.5 5.5e-08 
1.0 0.28 0 -4.5 5.5e-08 
1.0 0.3 0 -4.5 5.5e-08 
1.0 0.32 0 -4.5 5.5e-08 
1.0 0.34 0 -4.5 5.5e-08 
1.0 0.36 0 -4.5 5.5e-08 
1.0 0.38 0 -4.5 5.5e-08 
1.0 0.4 0 -4.5 5.5e-08 
1.0 0.42 0 -4.5 5.5e-08 
1.0 0.44 0 -4.5 5.5e-08 
1.0 0.46 0 -4.5 5.5e-08 
1.0 0.48 0 -4.5 5.5e-08 
1.0 0.5 0 -4.5 5.5e-08 
1.0 0.52 0 -4.5 5.5e-08 
1.0 0.54 0 -4.5 5.5e-08 
1.0 0.56 0 -4.5 5.5e-08 
1.0 0.58 0 -4.5 5.5e-08 
1.0 0.6 0 -4.5 5.5e-08 
1.0 0.62 0 -4.5 5.5e-08 
1.0 0.64 0 -4.5 5.5e-08 
1.0 0.66 0 -4.5 5.5e-08 
1.0 0.68 0 -4.5 5.5e-08 
1.0 0.7 0 -4.5 5.5e-08 
1.0 0.72 0 -4.5 5.5e-08 
1.0 0.74 0 -4.5 5.5e-08 
1.0 0.76 0 -4.5 5.5e-08 
1.0 0.78 0 -4.5 5.5e-08 
1.0 0.8 0 -4.5 5.5e-08 
1.0 0.82 0 -4.5 5.5e-08 
1.0 0.84 0 -4.5 5.5e-08 
1.0 0.86 0 -4.5 5.5e-08 
1.0 0.88 0 -4.5 5.5e-08 
1.0 0.9 0 -4.5 5.5e-08 
1.0 0.92 0 -4.5 5.5e-08 
1.0 0.94 0 -4.5 5.5e-08 
1.0 0.96 0 -4.5 5.5e-08 
1.0 0.98 0 -4.5 5.5e-08 
1.0 1.0 0 -4.5 5.5e-08 
1.0 1.02 0 -4.5 5.5e-08 
1.0 1.04 0 -4.5 5.5e-08 
1.0 1.06 0 -4.5 5.5e-08 
1.0 1.08 0 -4.5 5.5e-08 
1.0 1.1 0 -4.5 5.5e-08 
1.0 1.12 0 -4.5 5.5e-08 
1.0 1.14 0 -4.5 5.5e-08 
1.0 1.16 0 -4.5 5.5e-08 
1.0 1.18 0 -4.5 5.5e-08 
1.0 1.2 0 -4.5 5.5e-08 
1.0 1.22 0 -4.5 5.5e-08 
1.0 1.24 0 -4.5 5.5e-08 
1.0 1.26 0 -4.5 5.5e-08 
1.0 1.28 0 -4.5 5.5e-08 
1.0 1.3 0 -4.5 5.5e-08 
1.0 1.32 0 -4.5 5.5e-08 
1.0 1.34 0 -4.5 5.5e-08 
1.0 1.36 0 -4.5 5.5e-08 
1.0 1.38 0 -4.5 5.5e-08 
1.0 1.4 0 -4.5 5.5e-08 
1.0 1.42 0 -4.5 5.5e-08 
1.0 1.44 0 -4.5 5.5e-08 
1.0 1.46 0 -4.5 5.5e-08 
1.0 1.48 0 -4.5 5.5e-08 
1.0 -1.5 0 -5.0 5.5e-08 
1.0 -1.48 0 -5.0 5.5e-08 
1.0 -1.46 0 -5.0 5.5e-08 
1.0 -1.44 0 -5.0 5.5e-08 
1.0 -1.42 0 -5.0 5.5e-08 
1.0 -1.4 0 -5.0 5.5e-08 
1.0 -1.38 0 -5.0 5.5e-08 
1.0 -1.36 0 -5.0 5.5e-08 
1.0 -1.34 0 -5.0 5.5e-08 
1.0 -1.32 0 -5.0 5.5e-08 
1.0 -1.3 0 -5.0 5.5e-08 
1.0 -1.28 0 -5.0 5.5e-08 
1.0 -1.26 0 -5.0 5.5e-08 
1.0 -1.24 0 -5.0 5.5e-08 
1.0 -1.22 0 -5.0 5.5e-08 
1.0 -1.2 0 -5.0 5.5e-08 
1.0 -1.18 0 -5.0 5.5e-08 
1.0 -1.16 0 -5.0 5.5e-08 
1.0 -1.14 0 -5.0 5.5e-08 
1.0 -1.12 0 -5.0 5.5e-08 
1.0 -1.1 0 -5.0 5.5e-08 
1.0 -1.08 0 -5.0 5.5e-08 
1.0 -1.06 0 -5.0 5.5e-08 
1.0 -1.04 0 -5.0 5.5e-08 
1.0 -1.02 0 -5.0 5.5e-08 
1.0 -1.0 0 -5.0 5.5e-08 
1.0 -0.98 0 -5.0 5.5e-08 
1.0 -0.96 0 -5.0 5.5e-08 
1.0 -0.94 0 -5.0 5.5e-08 
1.0 -0.92 0 -5.0 5.5e-08 
1.0 -0.9 0 -5.0 5.5e-08 
1.0 -0.88 0 -5.0 5.5e-08 
1.0 -0.86 0 -5.0 5.5e-08 
1.0 -0.84 0 -5.0 5.5e-08 
1.0 -0.82 0 -5.0 5.5e-08 
1.0 -0.8 0 -5.0 5.5e-08 
1.0 -0.78 0 -5.0 5.5e-08 
1.0 -0.76 0 -5.0 5.5e-08 
1.0 -0.74 0 -5.0 5.5e-08 
1.0 -0.72 0 -5.0 5.5e-08 
1.0 -0.7 0 -5.0 5.5e-08 
1.0 -0.68 0 -5.0 5.5e-08 
1.0 -0.66 0 -5.0 5.5e-08 
1.0 -0.64 0 -5.0 5.5e-08 
1.0 -0.62 0 -5.0 5.5e-08 
1.0 -0.6 0 -5.0 5.5e-08 
1.0 -0.58 0 -5.0 5.5e-08 
1.0 -0.56 0 -5.0 5.5e-08 
1.0 -0.54 0 -5.0 5.5e-08 
1.0 -0.52 0 -5.0 5.5e-08 
1.0 -0.5 0 -5.0 5.5e-08 
1.0 -0.48 0 -5.0 5.5e-08 
1.0 -0.46 0 -5.0 5.5e-08 
1.0 -0.44 0 -5.0 5.5e-08 
1.0 -0.42 0 -5.0 5.5e-08 
1.0 -0.4 0 -5.0 5.5e-08 
1.0 -0.38 0 -5.0 5.5e-08 
1.0 -0.36 0 -5.0 5.5e-08 
1.0 -0.34 0 -5.0 5.5e-08 
1.0 -0.32 0 -5.0 5.5e-08 
1.0 -0.3 0 -5.0 5.5e-08 
1.0 -0.28 0 -5.0 5.5e-08 
1.0 -0.26 0 -5.0 5.5e-08 
1.0 -0.24 0 -5.0 5.5e-08 
1.0 -0.22 0 -5.0 5.5e-08 
1.0 -0.2 0 -5.0 5.5e-08 
1.0 -0.18 0 -5.0 5.5e-08 
1.0 -0.16 0 -5.0 5.5e-08 
1.0 -0.14 0 -5.0 5.5e-08 
1.0 -0.12 0 -5.0 5.5e-08 
1.0 -0.1 0 -5.0 5.5e-08 
1.0 -0.08 0 -5.0 5.5e-08 
1.0 -0.06 0 -5.0 5.5e-08 
1.0 -0.04 0 -5.0 5.5e-08 
1.0 -0.02 0 -5.0 5.5e-08 
1.0 1.33226762955e-15 0 -5.0 5.5e-08 
1.0 0.02 0 -5.0 5.5e-08 
1.0 0.04 0 -5.0 5.5e-08 
1.0 0.06 0 -5.0 5.5e-08 
1.0 0.08 0 -5.0 5.5e-08 
1.0 0.1 0 -5.0 5.5e-08 
1.0 0.12 0 -5.0 5.5e-08 
1.0 0.14 0 -5.0 5.5e-08 
1.0 0.16 0 -5.0 5.5e-08 
1.0 0.18 0 -5.0 5.5e-08 
1.0 0.2 0 -5.0 5.5e-08 
1.0 0.22 0 -5.0 5.5e-08 
1.0 0.24 0 -5.0 5.5e-08 
1.0 0.26 0 -5.0 5.5e-08 
1.0 0.28 0 -5.0 5.5e-08 
1.0 0.3 0 -5.0 5.5e-08 
1.0 0.32 0 -5.0 5.5e-08 
1.0 0.34 0 -5.0 5.5e-08 
1.0 0.36 0 -5.0 5.5e-08 
1.0 0.38 0 -5.0 5.5e-08 
1.0 0.4 0 -5.0 5.5e-08 
1.0 0.42 0 -5.0 5.5e-08 
1.0 0.44 0 -5.0 5.5e-08 
1.0 0.46 0 -5.0 5.5e-08 
1.0 0.48 0 -5.0 5.5e-08 
1.0 0.5 0 -5.0 5.5e-08 
1.0 0.52 0 -5.0 5.5e-08 
1.0 0.54 0 -5.0 5.5e-08 
1.0 0.56 0 -5.0 5.5e-08 
1.0 0.58 0 -5.0 5.5e-08 
1.0 0.6 0 -5.0 5.5e-08 
1.0 0.62 0 -5.0 5.5e-08 
1.0 0.64 0 -5.0 5.5e-08 
1.0 0.66 0 -5.0 5.5e-08 
1.0 0.68 0 -5.0 5.5e-08 
1.0 0.7 0 -5.0 5.5e-08 
1.0 0.72 0 -5.0 5.5e-08 
1.0 0.74 0 -5.0 5.5e-08 
1.0 0.76 0 -5.0 5.5e-08 
1.0 0.78 0 -5.0 5.5e-08 
1.0 0.8 0 -5.0 5.5e-08 
1.0 0.82 0 -5.0 5.5e-08 
1.0 0.84 0 -5.0 5.5e-08 
1.0 0.86 0 -5.0 5.5e-08 
1.0 0.88 0 -5.0 5.5e-08 
1.0 0.9 0 -5.0 5.5e-08 
1.0 0.92 0 -5.0 5.5e-08 
1.0 0.94 0 -5.0 5.5e-08 
1.0 0.96 0 -5.0 5.5e-08 
1.0 0.98 0 -5.0 5.5e-08 
1.0 1.0 0 -5.0 5.5e-08 
1.0 1.02 0 -5.0 5.5e-08 
1.0 1.04 0 -5.0 5.5e-08 
1.0 1.06 0 -5.0 5.5e-08 
1.0 1.08 0 -5.0 5.5e-08 
1.0 1.1 0 -5.0 5.5e-08 
1.0 1.12 0 -5.0 5.5e-08 
1.0 1.14 0 -5.0 5.5e-08 
1.0 1.16 0 -5.0 5.5e-08 
1.0 1.18 0 -5.0 5.5e-08 
1.0 1.2 0 -5.0 5.5e-08 
1.0 1.22 0 -5.0 5.5e-08 
1.0 1.24 0 -5.0 5.5e-08 
1.0 1.26 0 -5.0 5.5e-08 
1.0 1.28 0 -5.0 5.5e-08 
1.0 1.3 0 -5.0 5.5e-08 
1.0 1.32 0 -5.0 5.5e-08 
1.0 1.34 0 -5.0 5.5e-08 
1.0 1.36 0 -5.0 5.5e-08 
1.0 1.38 0 -5.0 5.5e-08 
1.0 1.4 0 -5.0 5.5e-08 
1.0 1.42 0 -5.0 5.5e-08 
1.0 1.44 0 -5.0 5.5e-08 
1.0 1.46 0 -5.0 5.5e-08 
1.0 1.48 0 -5.0 5.5e-08 
.ENDDATA 
.dc sweep DATA = datadc 
.print dc X1:IDS X1:qicore X1:xg1 X1:xg2 
.end