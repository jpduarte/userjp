*script to generate hspice simulation using cmdp, Juan Duarte 
*Date: 04/24/2015, time: 20:14:59

.option abstol=1e-6 reltol=1e-6 post ingold 
.option measform=1 
.temp 27 

.hdl "/users/jpduarte/BSIM_CM_Matlab/BSIM_model_development_v2/DM_Verilog_Hspice/Models_Verilog/BSIMIMGref/code/bsimimg.va" 
.include "/users/jpduarte/BSIM_CM_Matlab/BSIM_model_development_v2/DM_Verilog_Hspice/Models_Verilog/BSIMIMG/benchmark_tests/modelcard.pmos" 

.PARAM Vd_value = 0 
.PARAM Vgf_value = 0 
.PARAM Vs_value = 0 
.PARAM Vgb_value = 0 
.PARAM L_value = 1e-06 

Vd Vd 0.0 dc = Vd_value 
Vgf Vgf 0.0 dc = Vgf_value 
Vs Vs 0.0 dc = Vs_value 
Vgb Vgb 0.0 dc = Vgb_value 

X1 Vd Vgf Vs Vgb pmos1 L = 'L_value'

.DATA datadc Vd_value Vgf_value Vs_value Vgb_value L_value 
0.0 -1.0 1 1 1e-06 
0.95 -1.0 1 1 1e-06 
0.0 -0.979797979798 1 1 1e-06 
0.95 -0.979797979798 1 1 1e-06 
0.0 -0.959595959596 1 1 1e-06 
0.95 -0.959595959596 1 1 1e-06 
0.0 -0.939393939394 1 1 1e-06 
0.95 -0.939393939394 1 1 1e-06 
0.0 -0.919191919192 1 1 1e-06 
0.95 -0.919191919192 1 1 1e-06 
0.0 -0.89898989899 1 1 1e-06 
0.95 -0.89898989899 1 1 1e-06 
0.0 -0.878787878788 1 1 1e-06 
0.95 -0.878787878788 1 1 1e-06 
0.0 -0.858585858586 1 1 1e-06 
0.95 -0.858585858586 1 1 1e-06 
0.0 -0.838383838384 1 1 1e-06 
0.95 -0.838383838384 1 1 1e-06 
0.0 -0.818181818182 1 1 1e-06 
0.95 -0.818181818182 1 1 1e-06 
0.0 -0.79797979798 1 1 1e-06 
0.95 -0.79797979798 1 1 1e-06 
0.0 -0.777777777778 1 1 1e-06 
0.95 -0.777777777778 1 1 1e-06 
0.0 -0.757575757576 1 1 1e-06 
0.95 -0.757575757576 1 1 1e-06 
0.0 -0.737373737374 1 1 1e-06 
0.95 -0.737373737374 1 1 1e-06 
0.0 -0.717171717172 1 1 1e-06 
0.95 -0.717171717172 1 1 1e-06 
0.0 -0.69696969697 1 1 1e-06 
0.95 -0.69696969697 1 1 1e-06 
0.0 -0.676767676768 1 1 1e-06 
0.95 -0.676767676768 1 1 1e-06 
0.0 -0.656565656566 1 1 1e-06 
0.95 -0.656565656566 1 1 1e-06 
0.0 -0.636363636364 1 1 1e-06 
0.95 -0.636363636364 1 1 1e-06 
0.0 -0.616161616162 1 1 1e-06 
0.95 -0.616161616162 1 1 1e-06 
0.0 -0.59595959596 1 1 1e-06 
0.95 -0.59595959596 1 1 1e-06 
0.0 -0.575757575758 1 1 1e-06 
0.95 -0.575757575758 1 1 1e-06 
0.0 -0.555555555556 1 1 1e-06 
0.95 -0.555555555556 1 1 1e-06 
0.0 -0.535353535354 1 1 1e-06 
0.95 -0.535353535354 1 1 1e-06 
0.0 -0.515151515152 1 1 1e-06 
0.95 -0.515151515152 1 1 1e-06 
0.0 -0.494949494949 1 1 1e-06 
0.95 -0.494949494949 1 1 1e-06 
0.0 -0.474747474747 1 1 1e-06 
0.95 -0.474747474747 1 1 1e-06 
0.0 -0.454545454545 1 1 1e-06 
0.95 -0.454545454545 1 1 1e-06 
0.0 -0.434343434343 1 1 1e-06 
0.95 -0.434343434343 1 1 1e-06 
0.0 -0.414141414141 1 1 1e-06 
0.95 -0.414141414141 1 1 1e-06 
0.0 -0.393939393939 1 1 1e-06 
0.95 -0.393939393939 1 1 1e-06 
0.0 -0.373737373737 1 1 1e-06 
0.95 -0.373737373737 1 1 1e-06 
0.0 -0.353535353535 1 1 1e-06 
0.95 -0.353535353535 1 1 1e-06 
0.0 -0.333333333333 1 1 1e-06 
0.95 -0.333333333333 1 1 1e-06 
0.0 -0.313131313131 1 1 1e-06 
0.95 -0.313131313131 1 1 1e-06 
0.0 -0.292929292929 1 1 1e-06 
0.95 -0.292929292929 1 1 1e-06 
0.0 -0.272727272727 1 1 1e-06 
0.95 -0.272727272727 1 1 1e-06 
0.0 -0.252525252525 1 1 1e-06 
0.95 -0.252525252525 1 1 1e-06 
0.0 -0.232323232323 1 1 1e-06 
0.95 -0.232323232323 1 1 1e-06 
0.0 -0.212121212121 1 1 1e-06 
0.95 -0.212121212121 1 1 1e-06 
0.0 -0.191919191919 1 1 1e-06 
0.95 -0.191919191919 1 1 1e-06 
0.0 -0.171717171717 1 1 1e-06 
0.95 -0.171717171717 1 1 1e-06 
0.0 -0.151515151515 1 1 1e-06 
0.95 -0.151515151515 1 1 1e-06 
0.0 -0.131313131313 1 1 1e-06 
0.95 -0.131313131313 1 1 1e-06 
0.0 -0.111111111111 1 1 1e-06 
0.95 -0.111111111111 1 1 1e-06 
0.0 -0.0909090909091 1 1 1e-06 
0.95 -0.0909090909091 1 1 1e-06 
0.0 -0.0707070707071 1 1 1e-06 
0.95 -0.0707070707071 1 1 1e-06 
0.0 -0.0505050505051 1 1 1e-06 
0.95 -0.0505050505051 1 1 1e-06 
0.0 -0.030303030303 1 1 1e-06 
0.95 -0.030303030303 1 1 1e-06 
0.0 -0.010101010101 1 1 1e-06 
0.95 -0.010101010101 1 1 1e-06 
0.0 0.010101010101 1 1 1e-06 
0.95 0.010101010101 1 1 1e-06 
0.0 0.030303030303 1 1 1e-06 
0.95 0.030303030303 1 1 1e-06 
0.0 0.0505050505051 1 1 1e-06 
0.95 0.0505050505051 1 1 1e-06 
0.0 0.0707070707071 1 1 1e-06 
0.95 0.0707070707071 1 1 1e-06 
0.0 0.0909090909091 1 1 1e-06 
0.95 0.0909090909091 1 1 1e-06 
0.0 0.111111111111 1 1 1e-06 
0.95 0.111111111111 1 1 1e-06 
0.0 0.131313131313 1 1 1e-06 
0.95 0.131313131313 1 1 1e-06 
0.0 0.151515151515 1 1 1e-06 
0.95 0.151515151515 1 1 1e-06 
0.0 0.171717171717 1 1 1e-06 
0.95 0.171717171717 1 1 1e-06 
0.0 0.191919191919 1 1 1e-06 
0.95 0.191919191919 1 1 1e-06 
0.0 0.212121212121 1 1 1e-06 
0.95 0.212121212121 1 1 1e-06 
0.0 0.232323232323 1 1 1e-06 
0.95 0.232323232323 1 1 1e-06 
0.0 0.252525252525 1 1 1e-06 
0.95 0.252525252525 1 1 1e-06 
0.0 0.272727272727 1 1 1e-06 
0.95 0.272727272727 1 1 1e-06 
0.0 0.292929292929 1 1 1e-06 
0.95 0.292929292929 1 1 1e-06 
0.0 0.313131313131 1 1 1e-06 
0.95 0.313131313131 1 1 1e-06 
0.0 0.333333333333 1 1 1e-06 
0.95 0.333333333333 1 1 1e-06 
0.0 0.353535353535 1 1 1e-06 
0.95 0.353535353535 1 1 1e-06 
0.0 0.373737373737 1 1 1e-06 
0.95 0.373737373737 1 1 1e-06 
0.0 0.393939393939 1 1 1e-06 
0.95 0.393939393939 1 1 1e-06 
0.0 0.414141414141 1 1 1e-06 
0.95 0.414141414141 1 1 1e-06 
0.0 0.434343434343 1 1 1e-06 
0.95 0.434343434343 1 1 1e-06 
0.0 0.454545454545 1 1 1e-06 
0.95 0.454545454545 1 1 1e-06 
0.0 0.474747474747 1 1 1e-06 
0.95 0.474747474747 1 1 1e-06 
0.0 0.494949494949 1 1 1e-06 
0.95 0.494949494949 1 1 1e-06 
0.0 0.515151515152 1 1 1e-06 
0.95 0.515151515152 1 1 1e-06 
0.0 0.535353535354 1 1 1e-06 
0.95 0.535353535354 1 1 1e-06 
0.0 0.555555555556 1 1 1e-06 
0.95 0.555555555556 1 1 1e-06 
0.0 0.575757575758 1 1 1e-06 
0.95 0.575757575758 1 1 1e-06 
0.0 0.59595959596 1 1 1e-06 
0.95 0.59595959596 1 1 1e-06 
0.0 0.616161616162 1 1 1e-06 
0.95 0.616161616162 1 1 1e-06 
0.0 0.636363636364 1 1 1e-06 
0.95 0.636363636364 1 1 1e-06 
0.0 0.656565656566 1 1 1e-06 
0.95 0.656565656566 1 1 1e-06 
0.0 0.676767676768 1 1 1e-06 
0.95 0.676767676768 1 1 1e-06 
0.0 0.69696969697 1 1 1e-06 
0.95 0.69696969697 1 1 1e-06 
0.0 0.717171717172 1 1 1e-06 
0.95 0.717171717172 1 1 1e-06 
0.0 0.737373737374 1 1 1e-06 
0.95 0.737373737374 1 1 1e-06 
0.0 0.757575757576 1 1 1e-06 
0.95 0.757575757576 1 1 1e-06 
0.0 0.777777777778 1 1 1e-06 
0.95 0.777777777778 1 1 1e-06 
0.0 0.79797979798 1 1 1e-06 
0.95 0.79797979798 1 1 1e-06 
0.0 0.818181818182 1 1 1e-06 
0.95 0.818181818182 1 1 1e-06 
0.0 0.838383838384 1 1 1e-06 
0.95 0.838383838384 1 1 1e-06 
0.0 0.858585858586 1 1 1e-06 
0.95 0.858585858586 1 1 1e-06 
0.0 0.878787878788 1 1 1e-06 
0.95 0.878787878788 1 1 1e-06 
0.0 0.89898989899 1 1 1e-06 
0.95 0.89898989899 1 1 1e-06 
0.0 0.919191919192 1 1 1e-06 
0.95 0.919191919192 1 1 1e-06 
0.0 0.939393939394 1 1 1e-06 
0.95 0.939393939394 1 1 1e-06 
0.0 0.959595959596 1 1 1e-06 
0.95 0.959595959596 1 1 1e-06 
0.0 0.979797979798 1 1 1e-06 
0.95 0.979797979798 1 1 1e-06 
0.0 1.0 1 1 1e-06 
0.95 1.0 1 1 1e-06 
.ENDDATA 
.dc sweep DATA = datadc 
.print dc X1:IDS X1:qtotd X1:qtots X1:vbgs 
.end