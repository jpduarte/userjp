*script to generate hspice simulation using cmdp, Juan Duarte 
*Date: 09/22/2015, time: 20:17:46

.option abstol=1e-6 reltol=1e-6 post ingold 
.option measform=1 
.temp 27 

.hdl "/users/jpduarte/research/BSIMIMG/code/bsimimg.va" 
.include "/users/jpduarte/research/userjp/project2/modelcards/leapmodelcard.nmos" 

.PARAM Vd_value = 0 
.PARAM Vgf_value = 0 
.PARAM Vs_value = 0 
.PARAM Vgb_value = 0 
.PARAM L_value = 1e-06 

Vd Vd 0.0 dc = Vd_value 
Vgf Vgf 0.0 dc = Vgf_value 
Vs Vs 0.0 dc = Vs_value 
Vgb Vgb 0.0 dc = Vgb_value 

X1 Vd Vgf Vs Vgb nmos1 L = 'L_value'

.DATA datadc Vd_value Vgf_value Vs_value Vgb_value L_value 
0.5 -2.0 0 -2.0 1e-06 
0.555555555556 -2.0 0 -2.0 1e-06 
0.611111111111 -2.0 0 -2.0 1e-06 
0.666666666667 -2.0 0 -2.0 1e-06 
0.722222222222 -2.0 0 -2.0 1e-06 
0.777777777778 -2.0 0 -2.0 1e-06 
0.833333333333 -2.0 0 -2.0 1e-06 
0.888888888889 -2.0 0 -2.0 1e-06 
0.944444444444 -2.0 0 -2.0 1e-06 
1.0 -2.0 0 -2.0 1e-06 
0.5 -1.9595959596 0 -2.0 1e-06 
0.555555555556 -1.9595959596 0 -2.0 1e-06 
0.611111111111 -1.9595959596 0 -2.0 1e-06 
0.666666666667 -1.9595959596 0 -2.0 1e-06 
0.722222222222 -1.9595959596 0 -2.0 1e-06 
0.777777777778 -1.9595959596 0 -2.0 1e-06 
0.833333333333 -1.9595959596 0 -2.0 1e-06 
0.888888888889 -1.9595959596 0 -2.0 1e-06 
0.944444444444 -1.9595959596 0 -2.0 1e-06 
1.0 -1.9595959596 0 -2.0 1e-06 
0.5 -1.91919191919 0 -2.0 1e-06 
0.555555555556 -1.91919191919 0 -2.0 1e-06 
0.611111111111 -1.91919191919 0 -2.0 1e-06 
0.666666666667 -1.91919191919 0 -2.0 1e-06 
0.722222222222 -1.91919191919 0 -2.0 1e-06 
0.777777777778 -1.91919191919 0 -2.0 1e-06 
0.833333333333 -1.91919191919 0 -2.0 1e-06 
0.888888888889 -1.91919191919 0 -2.0 1e-06 
0.944444444444 -1.91919191919 0 -2.0 1e-06 
1.0 -1.91919191919 0 -2.0 1e-06 
0.5 -1.87878787879 0 -2.0 1e-06 
0.555555555556 -1.87878787879 0 -2.0 1e-06 
0.611111111111 -1.87878787879 0 -2.0 1e-06 
0.666666666667 -1.87878787879 0 -2.0 1e-06 
0.722222222222 -1.87878787879 0 -2.0 1e-06 
0.777777777778 -1.87878787879 0 -2.0 1e-06 
0.833333333333 -1.87878787879 0 -2.0 1e-06 
0.888888888889 -1.87878787879 0 -2.0 1e-06 
0.944444444444 -1.87878787879 0 -2.0 1e-06 
1.0 -1.87878787879 0 -2.0 1e-06 
0.5 -1.83838383838 0 -2.0 1e-06 
0.555555555556 -1.83838383838 0 -2.0 1e-06 
0.611111111111 -1.83838383838 0 -2.0 1e-06 
0.666666666667 -1.83838383838 0 -2.0 1e-06 
0.722222222222 -1.83838383838 0 -2.0 1e-06 
0.777777777778 -1.83838383838 0 -2.0 1e-06 
0.833333333333 -1.83838383838 0 -2.0 1e-06 
0.888888888889 -1.83838383838 0 -2.0 1e-06 
0.944444444444 -1.83838383838 0 -2.0 1e-06 
1.0 -1.83838383838 0 -2.0 1e-06 
0.5 -1.79797979798 0 -2.0 1e-06 
0.555555555556 -1.79797979798 0 -2.0 1e-06 
0.611111111111 -1.79797979798 0 -2.0 1e-06 
0.666666666667 -1.79797979798 0 -2.0 1e-06 
0.722222222222 -1.79797979798 0 -2.0 1e-06 
0.777777777778 -1.79797979798 0 -2.0 1e-06 
0.833333333333 -1.79797979798 0 -2.0 1e-06 
0.888888888889 -1.79797979798 0 -2.0 1e-06 
0.944444444444 -1.79797979798 0 -2.0 1e-06 
1.0 -1.79797979798 0 -2.0 1e-06 
0.5 -1.75757575758 0 -2.0 1e-06 
0.555555555556 -1.75757575758 0 -2.0 1e-06 
0.611111111111 -1.75757575758 0 -2.0 1e-06 
0.666666666667 -1.75757575758 0 -2.0 1e-06 
0.722222222222 -1.75757575758 0 -2.0 1e-06 
0.777777777778 -1.75757575758 0 -2.0 1e-06 
0.833333333333 -1.75757575758 0 -2.0 1e-06 
0.888888888889 -1.75757575758 0 -2.0 1e-06 
0.944444444444 -1.75757575758 0 -2.0 1e-06 
1.0 -1.75757575758 0 -2.0 1e-06 
0.5 -1.71717171717 0 -2.0 1e-06 
0.555555555556 -1.71717171717 0 -2.0 1e-06 
0.611111111111 -1.71717171717 0 -2.0 1e-06 
0.666666666667 -1.71717171717 0 -2.0 1e-06 
0.722222222222 -1.71717171717 0 -2.0 1e-06 
0.777777777778 -1.71717171717 0 -2.0 1e-06 
0.833333333333 -1.71717171717 0 -2.0 1e-06 
0.888888888889 -1.71717171717 0 -2.0 1e-06 
0.944444444444 -1.71717171717 0 -2.0 1e-06 
1.0 -1.71717171717 0 -2.0 1e-06 
0.5 -1.67676767677 0 -2.0 1e-06 
0.555555555556 -1.67676767677 0 -2.0 1e-06 
0.611111111111 -1.67676767677 0 -2.0 1e-06 
0.666666666667 -1.67676767677 0 -2.0 1e-06 
0.722222222222 -1.67676767677 0 -2.0 1e-06 
0.777777777778 -1.67676767677 0 -2.0 1e-06 
0.833333333333 -1.67676767677 0 -2.0 1e-06 
0.888888888889 -1.67676767677 0 -2.0 1e-06 
0.944444444444 -1.67676767677 0 -2.0 1e-06 
1.0 -1.67676767677 0 -2.0 1e-06 
0.5 -1.63636363636 0 -2.0 1e-06 
0.555555555556 -1.63636363636 0 -2.0 1e-06 
0.611111111111 -1.63636363636 0 -2.0 1e-06 
0.666666666667 -1.63636363636 0 -2.0 1e-06 
0.722222222222 -1.63636363636 0 -2.0 1e-06 
0.777777777778 -1.63636363636 0 -2.0 1e-06 
0.833333333333 -1.63636363636 0 -2.0 1e-06 
0.888888888889 -1.63636363636 0 -2.0 1e-06 
0.944444444444 -1.63636363636 0 -2.0 1e-06 
1.0 -1.63636363636 0 -2.0 1e-06 
0.5 -1.59595959596 0 -2.0 1e-06 
0.555555555556 -1.59595959596 0 -2.0 1e-06 
0.611111111111 -1.59595959596 0 -2.0 1e-06 
0.666666666667 -1.59595959596 0 -2.0 1e-06 
0.722222222222 -1.59595959596 0 -2.0 1e-06 
0.777777777778 -1.59595959596 0 -2.0 1e-06 
0.833333333333 -1.59595959596 0 -2.0 1e-06 
0.888888888889 -1.59595959596 0 -2.0 1e-06 
0.944444444444 -1.59595959596 0 -2.0 1e-06 
1.0 -1.59595959596 0 -2.0 1e-06 
0.5 -1.55555555556 0 -2.0 1e-06 
0.555555555556 -1.55555555556 0 -2.0 1e-06 
0.611111111111 -1.55555555556 0 -2.0 1e-06 
0.666666666667 -1.55555555556 0 -2.0 1e-06 
0.722222222222 -1.55555555556 0 -2.0 1e-06 
0.777777777778 -1.55555555556 0 -2.0 1e-06 
0.833333333333 -1.55555555556 0 -2.0 1e-06 
0.888888888889 -1.55555555556 0 -2.0 1e-06 
0.944444444444 -1.55555555556 0 -2.0 1e-06 
1.0 -1.55555555556 0 -2.0 1e-06 
0.5 -1.51515151515 0 -2.0 1e-06 
0.555555555556 -1.51515151515 0 -2.0 1e-06 
0.611111111111 -1.51515151515 0 -2.0 1e-06 
0.666666666667 -1.51515151515 0 -2.0 1e-06 
0.722222222222 -1.51515151515 0 -2.0 1e-06 
0.777777777778 -1.51515151515 0 -2.0 1e-06 
0.833333333333 -1.51515151515 0 -2.0 1e-06 
0.888888888889 -1.51515151515 0 -2.0 1e-06 
0.944444444444 -1.51515151515 0 -2.0 1e-06 
1.0 -1.51515151515 0 -2.0 1e-06 
0.5 -1.47474747475 0 -2.0 1e-06 
0.555555555556 -1.47474747475 0 -2.0 1e-06 
0.611111111111 -1.47474747475 0 -2.0 1e-06 
0.666666666667 -1.47474747475 0 -2.0 1e-06 
0.722222222222 -1.47474747475 0 -2.0 1e-06 
0.777777777778 -1.47474747475 0 -2.0 1e-06 
0.833333333333 -1.47474747475 0 -2.0 1e-06 
0.888888888889 -1.47474747475 0 -2.0 1e-06 
0.944444444444 -1.47474747475 0 -2.0 1e-06 
1.0 -1.47474747475 0 -2.0 1e-06 
0.5 -1.43434343434 0 -2.0 1e-06 
0.555555555556 -1.43434343434 0 -2.0 1e-06 
0.611111111111 -1.43434343434 0 -2.0 1e-06 
0.666666666667 -1.43434343434 0 -2.0 1e-06 
0.722222222222 -1.43434343434 0 -2.0 1e-06 
0.777777777778 -1.43434343434 0 -2.0 1e-06 
0.833333333333 -1.43434343434 0 -2.0 1e-06 
0.888888888889 -1.43434343434 0 -2.0 1e-06 
0.944444444444 -1.43434343434 0 -2.0 1e-06 
1.0 -1.43434343434 0 -2.0 1e-06 
0.5 -1.39393939394 0 -2.0 1e-06 
0.555555555556 -1.39393939394 0 -2.0 1e-06 
0.611111111111 -1.39393939394 0 -2.0 1e-06 
0.666666666667 -1.39393939394 0 -2.0 1e-06 
0.722222222222 -1.39393939394 0 -2.0 1e-06 
0.777777777778 -1.39393939394 0 -2.0 1e-06 
0.833333333333 -1.39393939394 0 -2.0 1e-06 
0.888888888889 -1.39393939394 0 -2.0 1e-06 
0.944444444444 -1.39393939394 0 -2.0 1e-06 
1.0 -1.39393939394 0 -2.0 1e-06 
0.5 -1.35353535354 0 -2.0 1e-06 
0.555555555556 -1.35353535354 0 -2.0 1e-06 
0.611111111111 -1.35353535354 0 -2.0 1e-06 
0.666666666667 -1.35353535354 0 -2.0 1e-06 
0.722222222222 -1.35353535354 0 -2.0 1e-06 
0.777777777778 -1.35353535354 0 -2.0 1e-06 
0.833333333333 -1.35353535354 0 -2.0 1e-06 
0.888888888889 -1.35353535354 0 -2.0 1e-06 
0.944444444444 -1.35353535354 0 -2.0 1e-06 
1.0 -1.35353535354 0 -2.0 1e-06 
0.5 -1.31313131313 0 -2.0 1e-06 
0.555555555556 -1.31313131313 0 -2.0 1e-06 
0.611111111111 -1.31313131313 0 -2.0 1e-06 
0.666666666667 -1.31313131313 0 -2.0 1e-06 
0.722222222222 -1.31313131313 0 -2.0 1e-06 
0.777777777778 -1.31313131313 0 -2.0 1e-06 
0.833333333333 -1.31313131313 0 -2.0 1e-06 
0.888888888889 -1.31313131313 0 -2.0 1e-06 
0.944444444444 -1.31313131313 0 -2.0 1e-06 
1.0 -1.31313131313 0 -2.0 1e-06 
0.5 -1.27272727273 0 -2.0 1e-06 
0.555555555556 -1.27272727273 0 -2.0 1e-06 
0.611111111111 -1.27272727273 0 -2.0 1e-06 
0.666666666667 -1.27272727273 0 -2.0 1e-06 
0.722222222222 -1.27272727273 0 -2.0 1e-06 
0.777777777778 -1.27272727273 0 -2.0 1e-06 
0.833333333333 -1.27272727273 0 -2.0 1e-06 
0.888888888889 -1.27272727273 0 -2.0 1e-06 
0.944444444444 -1.27272727273 0 -2.0 1e-06 
1.0 -1.27272727273 0 -2.0 1e-06 
0.5 -1.23232323232 0 -2.0 1e-06 
0.555555555556 -1.23232323232 0 -2.0 1e-06 
0.611111111111 -1.23232323232 0 -2.0 1e-06 
0.666666666667 -1.23232323232 0 -2.0 1e-06 
0.722222222222 -1.23232323232 0 -2.0 1e-06 
0.777777777778 -1.23232323232 0 -2.0 1e-06 
0.833333333333 -1.23232323232 0 -2.0 1e-06 
0.888888888889 -1.23232323232 0 -2.0 1e-06 
0.944444444444 -1.23232323232 0 -2.0 1e-06 
1.0 -1.23232323232 0 -2.0 1e-06 
0.5 -1.19191919192 0 -2.0 1e-06 
0.555555555556 -1.19191919192 0 -2.0 1e-06 
0.611111111111 -1.19191919192 0 -2.0 1e-06 
0.666666666667 -1.19191919192 0 -2.0 1e-06 
0.722222222222 -1.19191919192 0 -2.0 1e-06 
0.777777777778 -1.19191919192 0 -2.0 1e-06 
0.833333333333 -1.19191919192 0 -2.0 1e-06 
0.888888888889 -1.19191919192 0 -2.0 1e-06 
0.944444444444 -1.19191919192 0 -2.0 1e-06 
1.0 -1.19191919192 0 -2.0 1e-06 
0.5 -1.15151515152 0 -2.0 1e-06 
0.555555555556 -1.15151515152 0 -2.0 1e-06 
0.611111111111 -1.15151515152 0 -2.0 1e-06 
0.666666666667 -1.15151515152 0 -2.0 1e-06 
0.722222222222 -1.15151515152 0 -2.0 1e-06 
0.777777777778 -1.15151515152 0 -2.0 1e-06 
0.833333333333 -1.15151515152 0 -2.0 1e-06 
0.888888888889 -1.15151515152 0 -2.0 1e-06 
0.944444444444 -1.15151515152 0 -2.0 1e-06 
1.0 -1.15151515152 0 -2.0 1e-06 
0.5 -1.11111111111 0 -2.0 1e-06 
0.555555555556 -1.11111111111 0 -2.0 1e-06 
0.611111111111 -1.11111111111 0 -2.0 1e-06 
0.666666666667 -1.11111111111 0 -2.0 1e-06 
0.722222222222 -1.11111111111 0 -2.0 1e-06 
0.777777777778 -1.11111111111 0 -2.0 1e-06 
0.833333333333 -1.11111111111 0 -2.0 1e-06 
0.888888888889 -1.11111111111 0 -2.0 1e-06 
0.944444444444 -1.11111111111 0 -2.0 1e-06 
1.0 -1.11111111111 0 -2.0 1e-06 
0.5 -1.07070707071 0 -2.0 1e-06 
0.555555555556 -1.07070707071 0 -2.0 1e-06 
0.611111111111 -1.07070707071 0 -2.0 1e-06 
0.666666666667 -1.07070707071 0 -2.0 1e-06 
0.722222222222 -1.07070707071 0 -2.0 1e-06 
0.777777777778 -1.07070707071 0 -2.0 1e-06 
0.833333333333 -1.07070707071 0 -2.0 1e-06 
0.888888888889 -1.07070707071 0 -2.0 1e-06 
0.944444444444 -1.07070707071 0 -2.0 1e-06 
1.0 -1.07070707071 0 -2.0 1e-06 
0.5 -1.0303030303 0 -2.0 1e-06 
0.555555555556 -1.0303030303 0 -2.0 1e-06 
0.611111111111 -1.0303030303 0 -2.0 1e-06 
0.666666666667 -1.0303030303 0 -2.0 1e-06 
0.722222222222 -1.0303030303 0 -2.0 1e-06 
0.777777777778 -1.0303030303 0 -2.0 1e-06 
0.833333333333 -1.0303030303 0 -2.0 1e-06 
0.888888888889 -1.0303030303 0 -2.0 1e-06 
0.944444444444 -1.0303030303 0 -2.0 1e-06 
1.0 -1.0303030303 0 -2.0 1e-06 
0.5 -0.989898989899 0 -2.0 1e-06 
0.555555555556 -0.989898989899 0 -2.0 1e-06 
0.611111111111 -0.989898989899 0 -2.0 1e-06 
0.666666666667 -0.989898989899 0 -2.0 1e-06 
0.722222222222 -0.989898989899 0 -2.0 1e-06 
0.777777777778 -0.989898989899 0 -2.0 1e-06 
0.833333333333 -0.989898989899 0 -2.0 1e-06 
0.888888888889 -0.989898989899 0 -2.0 1e-06 
0.944444444444 -0.989898989899 0 -2.0 1e-06 
1.0 -0.989898989899 0 -2.0 1e-06 
0.5 -0.949494949495 0 -2.0 1e-06 
0.555555555556 -0.949494949495 0 -2.0 1e-06 
0.611111111111 -0.949494949495 0 -2.0 1e-06 
0.666666666667 -0.949494949495 0 -2.0 1e-06 
0.722222222222 -0.949494949495 0 -2.0 1e-06 
0.777777777778 -0.949494949495 0 -2.0 1e-06 
0.833333333333 -0.949494949495 0 -2.0 1e-06 
0.888888888889 -0.949494949495 0 -2.0 1e-06 
0.944444444444 -0.949494949495 0 -2.0 1e-06 
1.0 -0.949494949495 0 -2.0 1e-06 
0.5 -0.909090909091 0 -2.0 1e-06 
0.555555555556 -0.909090909091 0 -2.0 1e-06 
0.611111111111 -0.909090909091 0 -2.0 1e-06 
0.666666666667 -0.909090909091 0 -2.0 1e-06 
0.722222222222 -0.909090909091 0 -2.0 1e-06 
0.777777777778 -0.909090909091 0 -2.0 1e-06 
0.833333333333 -0.909090909091 0 -2.0 1e-06 
0.888888888889 -0.909090909091 0 -2.0 1e-06 
0.944444444444 -0.909090909091 0 -2.0 1e-06 
1.0 -0.909090909091 0 -2.0 1e-06 
0.5 -0.868686868687 0 -2.0 1e-06 
0.555555555556 -0.868686868687 0 -2.0 1e-06 
0.611111111111 -0.868686868687 0 -2.0 1e-06 
0.666666666667 -0.868686868687 0 -2.0 1e-06 
0.722222222222 -0.868686868687 0 -2.0 1e-06 
0.777777777778 -0.868686868687 0 -2.0 1e-06 
0.833333333333 -0.868686868687 0 -2.0 1e-06 
0.888888888889 -0.868686868687 0 -2.0 1e-06 
0.944444444444 -0.868686868687 0 -2.0 1e-06 
1.0 -0.868686868687 0 -2.0 1e-06 
0.5 -0.828282828283 0 -2.0 1e-06 
0.555555555556 -0.828282828283 0 -2.0 1e-06 
0.611111111111 -0.828282828283 0 -2.0 1e-06 
0.666666666667 -0.828282828283 0 -2.0 1e-06 
0.722222222222 -0.828282828283 0 -2.0 1e-06 
0.777777777778 -0.828282828283 0 -2.0 1e-06 
0.833333333333 -0.828282828283 0 -2.0 1e-06 
0.888888888889 -0.828282828283 0 -2.0 1e-06 
0.944444444444 -0.828282828283 0 -2.0 1e-06 
1.0 -0.828282828283 0 -2.0 1e-06 
0.5 -0.787878787879 0 -2.0 1e-06 
0.555555555556 -0.787878787879 0 -2.0 1e-06 
0.611111111111 -0.787878787879 0 -2.0 1e-06 
0.666666666667 -0.787878787879 0 -2.0 1e-06 
0.722222222222 -0.787878787879 0 -2.0 1e-06 
0.777777777778 -0.787878787879 0 -2.0 1e-06 
0.833333333333 -0.787878787879 0 -2.0 1e-06 
0.888888888889 -0.787878787879 0 -2.0 1e-06 
0.944444444444 -0.787878787879 0 -2.0 1e-06 
1.0 -0.787878787879 0 -2.0 1e-06 
0.5 -0.747474747475 0 -2.0 1e-06 
0.555555555556 -0.747474747475 0 -2.0 1e-06 
0.611111111111 -0.747474747475 0 -2.0 1e-06 
0.666666666667 -0.747474747475 0 -2.0 1e-06 
0.722222222222 -0.747474747475 0 -2.0 1e-06 
0.777777777778 -0.747474747475 0 -2.0 1e-06 
0.833333333333 -0.747474747475 0 -2.0 1e-06 
0.888888888889 -0.747474747475 0 -2.0 1e-06 
0.944444444444 -0.747474747475 0 -2.0 1e-06 
1.0 -0.747474747475 0 -2.0 1e-06 
0.5 -0.707070707071 0 -2.0 1e-06 
0.555555555556 -0.707070707071 0 -2.0 1e-06 
0.611111111111 -0.707070707071 0 -2.0 1e-06 
0.666666666667 -0.707070707071 0 -2.0 1e-06 
0.722222222222 -0.707070707071 0 -2.0 1e-06 
0.777777777778 -0.707070707071 0 -2.0 1e-06 
0.833333333333 -0.707070707071 0 -2.0 1e-06 
0.888888888889 -0.707070707071 0 -2.0 1e-06 
0.944444444444 -0.707070707071 0 -2.0 1e-06 
1.0 -0.707070707071 0 -2.0 1e-06 
0.5 -0.666666666667 0 -2.0 1e-06 
0.555555555556 -0.666666666667 0 -2.0 1e-06 
0.611111111111 -0.666666666667 0 -2.0 1e-06 
0.666666666667 -0.666666666667 0 -2.0 1e-06 
0.722222222222 -0.666666666667 0 -2.0 1e-06 
0.777777777778 -0.666666666667 0 -2.0 1e-06 
0.833333333333 -0.666666666667 0 -2.0 1e-06 
0.888888888889 -0.666666666667 0 -2.0 1e-06 
0.944444444444 -0.666666666667 0 -2.0 1e-06 
1.0 -0.666666666667 0 -2.0 1e-06 
0.5 -0.626262626263 0 -2.0 1e-06 
0.555555555556 -0.626262626263 0 -2.0 1e-06 
0.611111111111 -0.626262626263 0 -2.0 1e-06 
0.666666666667 -0.626262626263 0 -2.0 1e-06 
0.722222222222 -0.626262626263 0 -2.0 1e-06 
0.777777777778 -0.626262626263 0 -2.0 1e-06 
0.833333333333 -0.626262626263 0 -2.0 1e-06 
0.888888888889 -0.626262626263 0 -2.0 1e-06 
0.944444444444 -0.626262626263 0 -2.0 1e-06 
1.0 -0.626262626263 0 -2.0 1e-06 
0.5 -0.585858585859 0 -2.0 1e-06 
0.555555555556 -0.585858585859 0 -2.0 1e-06 
0.611111111111 -0.585858585859 0 -2.0 1e-06 
0.666666666667 -0.585858585859 0 -2.0 1e-06 
0.722222222222 -0.585858585859 0 -2.0 1e-06 
0.777777777778 -0.585858585859 0 -2.0 1e-06 
0.833333333333 -0.585858585859 0 -2.0 1e-06 
0.888888888889 -0.585858585859 0 -2.0 1e-06 
0.944444444444 -0.585858585859 0 -2.0 1e-06 
1.0 -0.585858585859 0 -2.0 1e-06 
0.5 -0.545454545455 0 -2.0 1e-06 
0.555555555556 -0.545454545455 0 -2.0 1e-06 
0.611111111111 -0.545454545455 0 -2.0 1e-06 
0.666666666667 -0.545454545455 0 -2.0 1e-06 
0.722222222222 -0.545454545455 0 -2.0 1e-06 
0.777777777778 -0.545454545455 0 -2.0 1e-06 
0.833333333333 -0.545454545455 0 -2.0 1e-06 
0.888888888889 -0.545454545455 0 -2.0 1e-06 
0.944444444444 -0.545454545455 0 -2.0 1e-06 
1.0 -0.545454545455 0 -2.0 1e-06 
0.5 -0.505050505051 0 -2.0 1e-06 
0.555555555556 -0.505050505051 0 -2.0 1e-06 
0.611111111111 -0.505050505051 0 -2.0 1e-06 
0.666666666667 -0.505050505051 0 -2.0 1e-06 
0.722222222222 -0.505050505051 0 -2.0 1e-06 
0.777777777778 -0.505050505051 0 -2.0 1e-06 
0.833333333333 -0.505050505051 0 -2.0 1e-06 
0.888888888889 -0.505050505051 0 -2.0 1e-06 
0.944444444444 -0.505050505051 0 -2.0 1e-06 
1.0 -0.505050505051 0 -2.0 1e-06 
0.5 -0.464646464646 0 -2.0 1e-06 
0.555555555556 -0.464646464646 0 -2.0 1e-06 
0.611111111111 -0.464646464646 0 -2.0 1e-06 
0.666666666667 -0.464646464646 0 -2.0 1e-06 
0.722222222222 -0.464646464646 0 -2.0 1e-06 
0.777777777778 -0.464646464646 0 -2.0 1e-06 
0.833333333333 -0.464646464646 0 -2.0 1e-06 
0.888888888889 -0.464646464646 0 -2.0 1e-06 
0.944444444444 -0.464646464646 0 -2.0 1e-06 
1.0 -0.464646464646 0 -2.0 1e-06 
0.5 -0.424242424242 0 -2.0 1e-06 
0.555555555556 -0.424242424242 0 -2.0 1e-06 
0.611111111111 -0.424242424242 0 -2.0 1e-06 
0.666666666667 -0.424242424242 0 -2.0 1e-06 
0.722222222222 -0.424242424242 0 -2.0 1e-06 
0.777777777778 -0.424242424242 0 -2.0 1e-06 
0.833333333333 -0.424242424242 0 -2.0 1e-06 
0.888888888889 -0.424242424242 0 -2.0 1e-06 
0.944444444444 -0.424242424242 0 -2.0 1e-06 
1.0 -0.424242424242 0 -2.0 1e-06 
0.5 -0.383838383838 0 -2.0 1e-06 
0.555555555556 -0.383838383838 0 -2.0 1e-06 
0.611111111111 -0.383838383838 0 -2.0 1e-06 
0.666666666667 -0.383838383838 0 -2.0 1e-06 
0.722222222222 -0.383838383838 0 -2.0 1e-06 
0.777777777778 -0.383838383838 0 -2.0 1e-06 
0.833333333333 -0.383838383838 0 -2.0 1e-06 
0.888888888889 -0.383838383838 0 -2.0 1e-06 
0.944444444444 -0.383838383838 0 -2.0 1e-06 
1.0 -0.383838383838 0 -2.0 1e-06 
0.5 -0.343434343434 0 -2.0 1e-06 
0.555555555556 -0.343434343434 0 -2.0 1e-06 
0.611111111111 -0.343434343434 0 -2.0 1e-06 
0.666666666667 -0.343434343434 0 -2.0 1e-06 
0.722222222222 -0.343434343434 0 -2.0 1e-06 
0.777777777778 -0.343434343434 0 -2.0 1e-06 
0.833333333333 -0.343434343434 0 -2.0 1e-06 
0.888888888889 -0.343434343434 0 -2.0 1e-06 
0.944444444444 -0.343434343434 0 -2.0 1e-06 
1.0 -0.343434343434 0 -2.0 1e-06 
0.5 -0.30303030303 0 -2.0 1e-06 
0.555555555556 -0.30303030303 0 -2.0 1e-06 
0.611111111111 -0.30303030303 0 -2.0 1e-06 
0.666666666667 -0.30303030303 0 -2.0 1e-06 
0.722222222222 -0.30303030303 0 -2.0 1e-06 
0.777777777778 -0.30303030303 0 -2.0 1e-06 
0.833333333333 -0.30303030303 0 -2.0 1e-06 
0.888888888889 -0.30303030303 0 -2.0 1e-06 
0.944444444444 -0.30303030303 0 -2.0 1e-06 
1.0 -0.30303030303 0 -2.0 1e-06 
0.5 -0.262626262626 0 -2.0 1e-06 
0.555555555556 -0.262626262626 0 -2.0 1e-06 
0.611111111111 -0.262626262626 0 -2.0 1e-06 
0.666666666667 -0.262626262626 0 -2.0 1e-06 
0.722222222222 -0.262626262626 0 -2.0 1e-06 
0.777777777778 -0.262626262626 0 -2.0 1e-06 
0.833333333333 -0.262626262626 0 -2.0 1e-06 
0.888888888889 -0.262626262626 0 -2.0 1e-06 
0.944444444444 -0.262626262626 0 -2.0 1e-06 
1.0 -0.262626262626 0 -2.0 1e-06 
0.5 -0.222222222222 0 -2.0 1e-06 
0.555555555556 -0.222222222222 0 -2.0 1e-06 
0.611111111111 -0.222222222222 0 -2.0 1e-06 
0.666666666667 -0.222222222222 0 -2.0 1e-06 
0.722222222222 -0.222222222222 0 -2.0 1e-06 
0.777777777778 -0.222222222222 0 -2.0 1e-06 
0.833333333333 -0.222222222222 0 -2.0 1e-06 
0.888888888889 -0.222222222222 0 -2.0 1e-06 
0.944444444444 -0.222222222222 0 -2.0 1e-06 
1.0 -0.222222222222 0 -2.0 1e-06 
0.5 -0.181818181818 0 -2.0 1e-06 
0.555555555556 -0.181818181818 0 -2.0 1e-06 
0.611111111111 -0.181818181818 0 -2.0 1e-06 
0.666666666667 -0.181818181818 0 -2.0 1e-06 
0.722222222222 -0.181818181818 0 -2.0 1e-06 
0.777777777778 -0.181818181818 0 -2.0 1e-06 
0.833333333333 -0.181818181818 0 -2.0 1e-06 
0.888888888889 -0.181818181818 0 -2.0 1e-06 
0.944444444444 -0.181818181818 0 -2.0 1e-06 
1.0 -0.181818181818 0 -2.0 1e-06 
0.5 -0.141414141414 0 -2.0 1e-06 
0.555555555556 -0.141414141414 0 -2.0 1e-06 
0.611111111111 -0.141414141414 0 -2.0 1e-06 
0.666666666667 -0.141414141414 0 -2.0 1e-06 
0.722222222222 -0.141414141414 0 -2.0 1e-06 
0.777777777778 -0.141414141414 0 -2.0 1e-06 
0.833333333333 -0.141414141414 0 -2.0 1e-06 
0.888888888889 -0.141414141414 0 -2.0 1e-06 
0.944444444444 -0.141414141414 0 -2.0 1e-06 
1.0 -0.141414141414 0 -2.0 1e-06 
0.5 -0.10101010101 0 -2.0 1e-06 
0.555555555556 -0.10101010101 0 -2.0 1e-06 
0.611111111111 -0.10101010101 0 -2.0 1e-06 
0.666666666667 -0.10101010101 0 -2.0 1e-06 
0.722222222222 -0.10101010101 0 -2.0 1e-06 
0.777777777778 -0.10101010101 0 -2.0 1e-06 
0.833333333333 -0.10101010101 0 -2.0 1e-06 
0.888888888889 -0.10101010101 0 -2.0 1e-06 
0.944444444444 -0.10101010101 0 -2.0 1e-06 
1.0 -0.10101010101 0 -2.0 1e-06 
0.5 -0.0606060606061 0 -2.0 1e-06 
0.555555555556 -0.0606060606061 0 -2.0 1e-06 
0.611111111111 -0.0606060606061 0 -2.0 1e-06 
0.666666666667 -0.0606060606061 0 -2.0 1e-06 
0.722222222222 -0.0606060606061 0 -2.0 1e-06 
0.777777777778 -0.0606060606061 0 -2.0 1e-06 
0.833333333333 -0.0606060606061 0 -2.0 1e-06 
0.888888888889 -0.0606060606061 0 -2.0 1e-06 
0.944444444444 -0.0606060606061 0 -2.0 1e-06 
1.0 -0.0606060606061 0 -2.0 1e-06 
0.5 -0.020202020202 0 -2.0 1e-06 
0.555555555556 -0.020202020202 0 -2.0 1e-06 
0.611111111111 -0.020202020202 0 -2.0 1e-06 
0.666666666667 -0.020202020202 0 -2.0 1e-06 
0.722222222222 -0.020202020202 0 -2.0 1e-06 
0.777777777778 -0.020202020202 0 -2.0 1e-06 
0.833333333333 -0.020202020202 0 -2.0 1e-06 
0.888888888889 -0.020202020202 0 -2.0 1e-06 
0.944444444444 -0.020202020202 0 -2.0 1e-06 
1.0 -0.020202020202 0 -2.0 1e-06 
0.5 0.020202020202 0 -2.0 1e-06 
0.555555555556 0.020202020202 0 -2.0 1e-06 
0.611111111111 0.020202020202 0 -2.0 1e-06 
0.666666666667 0.020202020202 0 -2.0 1e-06 
0.722222222222 0.020202020202 0 -2.0 1e-06 
0.777777777778 0.020202020202 0 -2.0 1e-06 
0.833333333333 0.020202020202 0 -2.0 1e-06 
0.888888888889 0.020202020202 0 -2.0 1e-06 
0.944444444444 0.020202020202 0 -2.0 1e-06 
1.0 0.020202020202 0 -2.0 1e-06 
0.5 0.0606060606061 0 -2.0 1e-06 
0.555555555556 0.0606060606061 0 -2.0 1e-06 
0.611111111111 0.0606060606061 0 -2.0 1e-06 
0.666666666667 0.0606060606061 0 -2.0 1e-06 
0.722222222222 0.0606060606061 0 -2.0 1e-06 
0.777777777778 0.0606060606061 0 -2.0 1e-06 
0.833333333333 0.0606060606061 0 -2.0 1e-06 
0.888888888889 0.0606060606061 0 -2.0 1e-06 
0.944444444444 0.0606060606061 0 -2.0 1e-06 
1.0 0.0606060606061 0 -2.0 1e-06 
0.5 0.10101010101 0 -2.0 1e-06 
0.555555555556 0.10101010101 0 -2.0 1e-06 
0.611111111111 0.10101010101 0 -2.0 1e-06 
0.666666666667 0.10101010101 0 -2.0 1e-06 
0.722222222222 0.10101010101 0 -2.0 1e-06 
0.777777777778 0.10101010101 0 -2.0 1e-06 
0.833333333333 0.10101010101 0 -2.0 1e-06 
0.888888888889 0.10101010101 0 -2.0 1e-06 
0.944444444444 0.10101010101 0 -2.0 1e-06 
1.0 0.10101010101 0 -2.0 1e-06 
0.5 0.141414141414 0 -2.0 1e-06 
0.555555555556 0.141414141414 0 -2.0 1e-06 
0.611111111111 0.141414141414 0 -2.0 1e-06 
0.666666666667 0.141414141414 0 -2.0 1e-06 
0.722222222222 0.141414141414 0 -2.0 1e-06 
0.777777777778 0.141414141414 0 -2.0 1e-06 
0.833333333333 0.141414141414 0 -2.0 1e-06 
0.888888888889 0.141414141414 0 -2.0 1e-06 
0.944444444444 0.141414141414 0 -2.0 1e-06 
1.0 0.141414141414 0 -2.0 1e-06 
0.5 0.181818181818 0 -2.0 1e-06 
0.555555555556 0.181818181818 0 -2.0 1e-06 
0.611111111111 0.181818181818 0 -2.0 1e-06 
0.666666666667 0.181818181818 0 -2.0 1e-06 
0.722222222222 0.181818181818 0 -2.0 1e-06 
0.777777777778 0.181818181818 0 -2.0 1e-06 
0.833333333333 0.181818181818 0 -2.0 1e-06 
0.888888888889 0.181818181818 0 -2.0 1e-06 
0.944444444444 0.181818181818 0 -2.0 1e-06 
1.0 0.181818181818 0 -2.0 1e-06 
0.5 0.222222222222 0 -2.0 1e-06 
0.555555555556 0.222222222222 0 -2.0 1e-06 
0.611111111111 0.222222222222 0 -2.0 1e-06 
0.666666666667 0.222222222222 0 -2.0 1e-06 
0.722222222222 0.222222222222 0 -2.0 1e-06 
0.777777777778 0.222222222222 0 -2.0 1e-06 
0.833333333333 0.222222222222 0 -2.0 1e-06 
0.888888888889 0.222222222222 0 -2.0 1e-06 
0.944444444444 0.222222222222 0 -2.0 1e-06 
1.0 0.222222222222 0 -2.0 1e-06 
0.5 0.262626262626 0 -2.0 1e-06 
0.555555555556 0.262626262626 0 -2.0 1e-06 
0.611111111111 0.262626262626 0 -2.0 1e-06 
0.666666666667 0.262626262626 0 -2.0 1e-06 
0.722222222222 0.262626262626 0 -2.0 1e-06 
0.777777777778 0.262626262626 0 -2.0 1e-06 
0.833333333333 0.262626262626 0 -2.0 1e-06 
0.888888888889 0.262626262626 0 -2.0 1e-06 
0.944444444444 0.262626262626 0 -2.0 1e-06 
1.0 0.262626262626 0 -2.0 1e-06 
0.5 0.30303030303 0 -2.0 1e-06 
0.555555555556 0.30303030303 0 -2.0 1e-06 
0.611111111111 0.30303030303 0 -2.0 1e-06 
0.666666666667 0.30303030303 0 -2.0 1e-06 
0.722222222222 0.30303030303 0 -2.0 1e-06 
0.777777777778 0.30303030303 0 -2.0 1e-06 
0.833333333333 0.30303030303 0 -2.0 1e-06 
0.888888888889 0.30303030303 0 -2.0 1e-06 
0.944444444444 0.30303030303 0 -2.0 1e-06 
1.0 0.30303030303 0 -2.0 1e-06 
0.5 0.343434343434 0 -2.0 1e-06 
0.555555555556 0.343434343434 0 -2.0 1e-06 
0.611111111111 0.343434343434 0 -2.0 1e-06 
0.666666666667 0.343434343434 0 -2.0 1e-06 
0.722222222222 0.343434343434 0 -2.0 1e-06 
0.777777777778 0.343434343434 0 -2.0 1e-06 
0.833333333333 0.343434343434 0 -2.0 1e-06 
0.888888888889 0.343434343434 0 -2.0 1e-06 
0.944444444444 0.343434343434 0 -2.0 1e-06 
1.0 0.343434343434 0 -2.0 1e-06 
0.5 0.383838383838 0 -2.0 1e-06 
0.555555555556 0.383838383838 0 -2.0 1e-06 
0.611111111111 0.383838383838 0 -2.0 1e-06 
0.666666666667 0.383838383838 0 -2.0 1e-06 
0.722222222222 0.383838383838 0 -2.0 1e-06 
0.777777777778 0.383838383838 0 -2.0 1e-06 
0.833333333333 0.383838383838 0 -2.0 1e-06 
0.888888888889 0.383838383838 0 -2.0 1e-06 
0.944444444444 0.383838383838 0 -2.0 1e-06 
1.0 0.383838383838 0 -2.0 1e-06 
0.5 0.424242424242 0 -2.0 1e-06 
0.555555555556 0.424242424242 0 -2.0 1e-06 
0.611111111111 0.424242424242 0 -2.0 1e-06 
0.666666666667 0.424242424242 0 -2.0 1e-06 
0.722222222222 0.424242424242 0 -2.0 1e-06 
0.777777777778 0.424242424242 0 -2.0 1e-06 
0.833333333333 0.424242424242 0 -2.0 1e-06 
0.888888888889 0.424242424242 0 -2.0 1e-06 
0.944444444444 0.424242424242 0 -2.0 1e-06 
1.0 0.424242424242 0 -2.0 1e-06 
0.5 0.464646464646 0 -2.0 1e-06 
0.555555555556 0.464646464646 0 -2.0 1e-06 
0.611111111111 0.464646464646 0 -2.0 1e-06 
0.666666666667 0.464646464646 0 -2.0 1e-06 
0.722222222222 0.464646464646 0 -2.0 1e-06 
0.777777777778 0.464646464646 0 -2.0 1e-06 
0.833333333333 0.464646464646 0 -2.0 1e-06 
0.888888888889 0.464646464646 0 -2.0 1e-06 
0.944444444444 0.464646464646 0 -2.0 1e-06 
1.0 0.464646464646 0 -2.0 1e-06 
0.5 0.505050505051 0 -2.0 1e-06 
0.555555555556 0.505050505051 0 -2.0 1e-06 
0.611111111111 0.505050505051 0 -2.0 1e-06 
0.666666666667 0.505050505051 0 -2.0 1e-06 
0.722222222222 0.505050505051 0 -2.0 1e-06 
0.777777777778 0.505050505051 0 -2.0 1e-06 
0.833333333333 0.505050505051 0 -2.0 1e-06 
0.888888888889 0.505050505051 0 -2.0 1e-06 
0.944444444444 0.505050505051 0 -2.0 1e-06 
1.0 0.505050505051 0 -2.0 1e-06 
0.5 0.545454545455 0 -2.0 1e-06 
0.555555555556 0.545454545455 0 -2.0 1e-06 
0.611111111111 0.545454545455 0 -2.0 1e-06 
0.666666666667 0.545454545455 0 -2.0 1e-06 
0.722222222222 0.545454545455 0 -2.0 1e-06 
0.777777777778 0.545454545455 0 -2.0 1e-06 
0.833333333333 0.545454545455 0 -2.0 1e-06 
0.888888888889 0.545454545455 0 -2.0 1e-06 
0.944444444444 0.545454545455 0 -2.0 1e-06 
1.0 0.545454545455 0 -2.0 1e-06 
0.5 0.585858585859 0 -2.0 1e-06 
0.555555555556 0.585858585859 0 -2.0 1e-06 
0.611111111111 0.585858585859 0 -2.0 1e-06 
0.666666666667 0.585858585859 0 -2.0 1e-06 
0.722222222222 0.585858585859 0 -2.0 1e-06 
0.777777777778 0.585858585859 0 -2.0 1e-06 
0.833333333333 0.585858585859 0 -2.0 1e-06 
0.888888888889 0.585858585859 0 -2.0 1e-06 
0.944444444444 0.585858585859 0 -2.0 1e-06 
1.0 0.585858585859 0 -2.0 1e-06 
0.5 0.626262626263 0 -2.0 1e-06 
0.555555555556 0.626262626263 0 -2.0 1e-06 
0.611111111111 0.626262626263 0 -2.0 1e-06 
0.666666666667 0.626262626263 0 -2.0 1e-06 
0.722222222222 0.626262626263 0 -2.0 1e-06 
0.777777777778 0.626262626263 0 -2.0 1e-06 
0.833333333333 0.626262626263 0 -2.0 1e-06 
0.888888888889 0.626262626263 0 -2.0 1e-06 
0.944444444444 0.626262626263 0 -2.0 1e-06 
1.0 0.626262626263 0 -2.0 1e-06 
0.5 0.666666666667 0 -2.0 1e-06 
0.555555555556 0.666666666667 0 -2.0 1e-06 
0.611111111111 0.666666666667 0 -2.0 1e-06 
0.666666666667 0.666666666667 0 -2.0 1e-06 
0.722222222222 0.666666666667 0 -2.0 1e-06 
0.777777777778 0.666666666667 0 -2.0 1e-06 
0.833333333333 0.666666666667 0 -2.0 1e-06 
0.888888888889 0.666666666667 0 -2.0 1e-06 
0.944444444444 0.666666666667 0 -2.0 1e-06 
1.0 0.666666666667 0 -2.0 1e-06 
0.5 0.707070707071 0 -2.0 1e-06 
0.555555555556 0.707070707071 0 -2.0 1e-06 
0.611111111111 0.707070707071 0 -2.0 1e-06 
0.666666666667 0.707070707071 0 -2.0 1e-06 
0.722222222222 0.707070707071 0 -2.0 1e-06 
0.777777777778 0.707070707071 0 -2.0 1e-06 
0.833333333333 0.707070707071 0 -2.0 1e-06 
0.888888888889 0.707070707071 0 -2.0 1e-06 
0.944444444444 0.707070707071 0 -2.0 1e-06 
1.0 0.707070707071 0 -2.0 1e-06 
0.5 0.747474747475 0 -2.0 1e-06 
0.555555555556 0.747474747475 0 -2.0 1e-06 
0.611111111111 0.747474747475 0 -2.0 1e-06 
0.666666666667 0.747474747475 0 -2.0 1e-06 
0.722222222222 0.747474747475 0 -2.0 1e-06 
0.777777777778 0.747474747475 0 -2.0 1e-06 
0.833333333333 0.747474747475 0 -2.0 1e-06 
0.888888888889 0.747474747475 0 -2.0 1e-06 
0.944444444444 0.747474747475 0 -2.0 1e-06 
1.0 0.747474747475 0 -2.0 1e-06 
0.5 0.787878787879 0 -2.0 1e-06 
0.555555555556 0.787878787879 0 -2.0 1e-06 
0.611111111111 0.787878787879 0 -2.0 1e-06 
0.666666666667 0.787878787879 0 -2.0 1e-06 
0.722222222222 0.787878787879 0 -2.0 1e-06 
0.777777777778 0.787878787879 0 -2.0 1e-06 
0.833333333333 0.787878787879 0 -2.0 1e-06 
0.888888888889 0.787878787879 0 -2.0 1e-06 
0.944444444444 0.787878787879 0 -2.0 1e-06 
1.0 0.787878787879 0 -2.0 1e-06 
0.5 0.828282828283 0 -2.0 1e-06 
0.555555555556 0.828282828283 0 -2.0 1e-06 
0.611111111111 0.828282828283 0 -2.0 1e-06 
0.666666666667 0.828282828283 0 -2.0 1e-06 
0.722222222222 0.828282828283 0 -2.0 1e-06 
0.777777777778 0.828282828283 0 -2.0 1e-06 
0.833333333333 0.828282828283 0 -2.0 1e-06 
0.888888888889 0.828282828283 0 -2.0 1e-06 
0.944444444444 0.828282828283 0 -2.0 1e-06 
1.0 0.828282828283 0 -2.0 1e-06 
0.5 0.868686868687 0 -2.0 1e-06 
0.555555555556 0.868686868687 0 -2.0 1e-06 
0.611111111111 0.868686868687 0 -2.0 1e-06 
0.666666666667 0.868686868687 0 -2.0 1e-06 
0.722222222222 0.868686868687 0 -2.0 1e-06 
0.777777777778 0.868686868687 0 -2.0 1e-06 
0.833333333333 0.868686868687 0 -2.0 1e-06 
0.888888888889 0.868686868687 0 -2.0 1e-06 
0.944444444444 0.868686868687 0 -2.0 1e-06 
1.0 0.868686868687 0 -2.0 1e-06 
0.5 0.909090909091 0 -2.0 1e-06 
0.555555555556 0.909090909091 0 -2.0 1e-06 
0.611111111111 0.909090909091 0 -2.0 1e-06 
0.666666666667 0.909090909091 0 -2.0 1e-06 
0.722222222222 0.909090909091 0 -2.0 1e-06 
0.777777777778 0.909090909091 0 -2.0 1e-06 
0.833333333333 0.909090909091 0 -2.0 1e-06 
0.888888888889 0.909090909091 0 -2.0 1e-06 
0.944444444444 0.909090909091 0 -2.0 1e-06 
1.0 0.909090909091 0 -2.0 1e-06 
0.5 0.949494949495 0 -2.0 1e-06 
0.555555555556 0.949494949495 0 -2.0 1e-06 
0.611111111111 0.949494949495 0 -2.0 1e-06 
0.666666666667 0.949494949495 0 -2.0 1e-06 
0.722222222222 0.949494949495 0 -2.0 1e-06 
0.777777777778 0.949494949495 0 -2.0 1e-06 
0.833333333333 0.949494949495 0 -2.0 1e-06 
0.888888888889 0.949494949495 0 -2.0 1e-06 
0.944444444444 0.949494949495 0 -2.0 1e-06 
1.0 0.949494949495 0 -2.0 1e-06 
0.5 0.989898989899 0 -2.0 1e-06 
0.555555555556 0.989898989899 0 -2.0 1e-06 
0.611111111111 0.989898989899 0 -2.0 1e-06 
0.666666666667 0.989898989899 0 -2.0 1e-06 
0.722222222222 0.989898989899 0 -2.0 1e-06 
0.777777777778 0.989898989899 0 -2.0 1e-06 
0.833333333333 0.989898989899 0 -2.0 1e-06 
0.888888888889 0.989898989899 0 -2.0 1e-06 
0.944444444444 0.989898989899 0 -2.0 1e-06 
1.0 0.989898989899 0 -2.0 1e-06 
0.5 1.0303030303 0 -2.0 1e-06 
0.555555555556 1.0303030303 0 -2.0 1e-06 
0.611111111111 1.0303030303 0 -2.0 1e-06 
0.666666666667 1.0303030303 0 -2.0 1e-06 
0.722222222222 1.0303030303 0 -2.0 1e-06 
0.777777777778 1.0303030303 0 -2.0 1e-06 
0.833333333333 1.0303030303 0 -2.0 1e-06 
0.888888888889 1.0303030303 0 -2.0 1e-06 
0.944444444444 1.0303030303 0 -2.0 1e-06 
1.0 1.0303030303 0 -2.0 1e-06 
0.5 1.07070707071 0 -2.0 1e-06 
0.555555555556 1.07070707071 0 -2.0 1e-06 
0.611111111111 1.07070707071 0 -2.0 1e-06 
0.666666666667 1.07070707071 0 -2.0 1e-06 
0.722222222222 1.07070707071 0 -2.0 1e-06 
0.777777777778 1.07070707071 0 -2.0 1e-06 
0.833333333333 1.07070707071 0 -2.0 1e-06 
0.888888888889 1.07070707071 0 -2.0 1e-06 
0.944444444444 1.07070707071 0 -2.0 1e-06 
1.0 1.07070707071 0 -2.0 1e-06 
0.5 1.11111111111 0 -2.0 1e-06 
0.555555555556 1.11111111111 0 -2.0 1e-06 
0.611111111111 1.11111111111 0 -2.0 1e-06 
0.666666666667 1.11111111111 0 -2.0 1e-06 
0.722222222222 1.11111111111 0 -2.0 1e-06 
0.777777777778 1.11111111111 0 -2.0 1e-06 
0.833333333333 1.11111111111 0 -2.0 1e-06 
0.888888888889 1.11111111111 0 -2.0 1e-06 
0.944444444444 1.11111111111 0 -2.0 1e-06 
1.0 1.11111111111 0 -2.0 1e-06 
0.5 1.15151515152 0 -2.0 1e-06 
0.555555555556 1.15151515152 0 -2.0 1e-06 
0.611111111111 1.15151515152 0 -2.0 1e-06 
0.666666666667 1.15151515152 0 -2.0 1e-06 
0.722222222222 1.15151515152 0 -2.0 1e-06 
0.777777777778 1.15151515152 0 -2.0 1e-06 
0.833333333333 1.15151515152 0 -2.0 1e-06 
0.888888888889 1.15151515152 0 -2.0 1e-06 
0.944444444444 1.15151515152 0 -2.0 1e-06 
1.0 1.15151515152 0 -2.0 1e-06 
0.5 1.19191919192 0 -2.0 1e-06 
0.555555555556 1.19191919192 0 -2.0 1e-06 
0.611111111111 1.19191919192 0 -2.0 1e-06 
0.666666666667 1.19191919192 0 -2.0 1e-06 
0.722222222222 1.19191919192 0 -2.0 1e-06 
0.777777777778 1.19191919192 0 -2.0 1e-06 
0.833333333333 1.19191919192 0 -2.0 1e-06 
0.888888888889 1.19191919192 0 -2.0 1e-06 
0.944444444444 1.19191919192 0 -2.0 1e-06 
1.0 1.19191919192 0 -2.0 1e-06 
0.5 1.23232323232 0 -2.0 1e-06 
0.555555555556 1.23232323232 0 -2.0 1e-06 
0.611111111111 1.23232323232 0 -2.0 1e-06 
0.666666666667 1.23232323232 0 -2.0 1e-06 
0.722222222222 1.23232323232 0 -2.0 1e-06 
0.777777777778 1.23232323232 0 -2.0 1e-06 
0.833333333333 1.23232323232 0 -2.0 1e-06 
0.888888888889 1.23232323232 0 -2.0 1e-06 
0.944444444444 1.23232323232 0 -2.0 1e-06 
1.0 1.23232323232 0 -2.0 1e-06 
0.5 1.27272727273 0 -2.0 1e-06 
0.555555555556 1.27272727273 0 -2.0 1e-06 
0.611111111111 1.27272727273 0 -2.0 1e-06 
0.666666666667 1.27272727273 0 -2.0 1e-06 
0.722222222222 1.27272727273 0 -2.0 1e-06 
0.777777777778 1.27272727273 0 -2.0 1e-06 
0.833333333333 1.27272727273 0 -2.0 1e-06 
0.888888888889 1.27272727273 0 -2.0 1e-06 
0.944444444444 1.27272727273 0 -2.0 1e-06 
1.0 1.27272727273 0 -2.0 1e-06 
0.5 1.31313131313 0 -2.0 1e-06 
0.555555555556 1.31313131313 0 -2.0 1e-06 
0.611111111111 1.31313131313 0 -2.0 1e-06 
0.666666666667 1.31313131313 0 -2.0 1e-06 
0.722222222222 1.31313131313 0 -2.0 1e-06 
0.777777777778 1.31313131313 0 -2.0 1e-06 
0.833333333333 1.31313131313 0 -2.0 1e-06 
0.888888888889 1.31313131313 0 -2.0 1e-06 
0.944444444444 1.31313131313 0 -2.0 1e-06 
1.0 1.31313131313 0 -2.0 1e-06 
0.5 1.35353535354 0 -2.0 1e-06 
0.555555555556 1.35353535354 0 -2.0 1e-06 
0.611111111111 1.35353535354 0 -2.0 1e-06 
0.666666666667 1.35353535354 0 -2.0 1e-06 
0.722222222222 1.35353535354 0 -2.0 1e-06 
0.777777777778 1.35353535354 0 -2.0 1e-06 
0.833333333333 1.35353535354 0 -2.0 1e-06 
0.888888888889 1.35353535354 0 -2.0 1e-06 
0.944444444444 1.35353535354 0 -2.0 1e-06 
1.0 1.35353535354 0 -2.0 1e-06 
0.5 1.39393939394 0 -2.0 1e-06 
0.555555555556 1.39393939394 0 -2.0 1e-06 
0.611111111111 1.39393939394 0 -2.0 1e-06 
0.666666666667 1.39393939394 0 -2.0 1e-06 
0.722222222222 1.39393939394 0 -2.0 1e-06 
0.777777777778 1.39393939394 0 -2.0 1e-06 
0.833333333333 1.39393939394 0 -2.0 1e-06 
0.888888888889 1.39393939394 0 -2.0 1e-06 
0.944444444444 1.39393939394 0 -2.0 1e-06 
1.0 1.39393939394 0 -2.0 1e-06 
0.5 1.43434343434 0 -2.0 1e-06 
0.555555555556 1.43434343434 0 -2.0 1e-06 
0.611111111111 1.43434343434 0 -2.0 1e-06 
0.666666666667 1.43434343434 0 -2.0 1e-06 
0.722222222222 1.43434343434 0 -2.0 1e-06 
0.777777777778 1.43434343434 0 -2.0 1e-06 
0.833333333333 1.43434343434 0 -2.0 1e-06 
0.888888888889 1.43434343434 0 -2.0 1e-06 
0.944444444444 1.43434343434 0 -2.0 1e-06 
1.0 1.43434343434 0 -2.0 1e-06 
0.5 1.47474747475 0 -2.0 1e-06 
0.555555555556 1.47474747475 0 -2.0 1e-06 
0.611111111111 1.47474747475 0 -2.0 1e-06 
0.666666666667 1.47474747475 0 -2.0 1e-06 
0.722222222222 1.47474747475 0 -2.0 1e-06 
0.777777777778 1.47474747475 0 -2.0 1e-06 
0.833333333333 1.47474747475 0 -2.0 1e-06 
0.888888888889 1.47474747475 0 -2.0 1e-06 
0.944444444444 1.47474747475 0 -2.0 1e-06 
1.0 1.47474747475 0 -2.0 1e-06 
0.5 1.51515151515 0 -2.0 1e-06 
0.555555555556 1.51515151515 0 -2.0 1e-06 
0.611111111111 1.51515151515 0 -2.0 1e-06 
0.666666666667 1.51515151515 0 -2.0 1e-06 
0.722222222222 1.51515151515 0 -2.0 1e-06 
0.777777777778 1.51515151515 0 -2.0 1e-06 
0.833333333333 1.51515151515 0 -2.0 1e-06 
0.888888888889 1.51515151515 0 -2.0 1e-06 
0.944444444444 1.51515151515 0 -2.0 1e-06 
1.0 1.51515151515 0 -2.0 1e-06 
0.5 1.55555555556 0 -2.0 1e-06 
0.555555555556 1.55555555556 0 -2.0 1e-06 
0.611111111111 1.55555555556 0 -2.0 1e-06 
0.666666666667 1.55555555556 0 -2.0 1e-06 
0.722222222222 1.55555555556 0 -2.0 1e-06 
0.777777777778 1.55555555556 0 -2.0 1e-06 
0.833333333333 1.55555555556 0 -2.0 1e-06 
0.888888888889 1.55555555556 0 -2.0 1e-06 
0.944444444444 1.55555555556 0 -2.0 1e-06 
1.0 1.55555555556 0 -2.0 1e-06 
0.5 1.59595959596 0 -2.0 1e-06 
0.555555555556 1.59595959596 0 -2.0 1e-06 
0.611111111111 1.59595959596 0 -2.0 1e-06 
0.666666666667 1.59595959596 0 -2.0 1e-06 
0.722222222222 1.59595959596 0 -2.0 1e-06 
0.777777777778 1.59595959596 0 -2.0 1e-06 
0.833333333333 1.59595959596 0 -2.0 1e-06 
0.888888888889 1.59595959596 0 -2.0 1e-06 
0.944444444444 1.59595959596 0 -2.0 1e-06 
1.0 1.59595959596 0 -2.0 1e-06 
0.5 1.63636363636 0 -2.0 1e-06 
0.555555555556 1.63636363636 0 -2.0 1e-06 
0.611111111111 1.63636363636 0 -2.0 1e-06 
0.666666666667 1.63636363636 0 -2.0 1e-06 
0.722222222222 1.63636363636 0 -2.0 1e-06 
0.777777777778 1.63636363636 0 -2.0 1e-06 
0.833333333333 1.63636363636 0 -2.0 1e-06 
0.888888888889 1.63636363636 0 -2.0 1e-06 
0.944444444444 1.63636363636 0 -2.0 1e-06 
1.0 1.63636363636 0 -2.0 1e-06 
0.5 1.67676767677 0 -2.0 1e-06 
0.555555555556 1.67676767677 0 -2.0 1e-06 
0.611111111111 1.67676767677 0 -2.0 1e-06 
0.666666666667 1.67676767677 0 -2.0 1e-06 
0.722222222222 1.67676767677 0 -2.0 1e-06 
0.777777777778 1.67676767677 0 -2.0 1e-06 
0.833333333333 1.67676767677 0 -2.0 1e-06 
0.888888888889 1.67676767677 0 -2.0 1e-06 
0.944444444444 1.67676767677 0 -2.0 1e-06 
1.0 1.67676767677 0 -2.0 1e-06 
0.5 1.71717171717 0 -2.0 1e-06 
0.555555555556 1.71717171717 0 -2.0 1e-06 
0.611111111111 1.71717171717 0 -2.0 1e-06 
0.666666666667 1.71717171717 0 -2.0 1e-06 
0.722222222222 1.71717171717 0 -2.0 1e-06 
0.777777777778 1.71717171717 0 -2.0 1e-06 
0.833333333333 1.71717171717 0 -2.0 1e-06 
0.888888888889 1.71717171717 0 -2.0 1e-06 
0.944444444444 1.71717171717 0 -2.0 1e-06 
1.0 1.71717171717 0 -2.0 1e-06 
0.5 1.75757575758 0 -2.0 1e-06 
0.555555555556 1.75757575758 0 -2.0 1e-06 
0.611111111111 1.75757575758 0 -2.0 1e-06 
0.666666666667 1.75757575758 0 -2.0 1e-06 
0.722222222222 1.75757575758 0 -2.0 1e-06 
0.777777777778 1.75757575758 0 -2.0 1e-06 
0.833333333333 1.75757575758 0 -2.0 1e-06 
0.888888888889 1.75757575758 0 -2.0 1e-06 
0.944444444444 1.75757575758 0 -2.0 1e-06 
1.0 1.75757575758 0 -2.0 1e-06 
0.5 1.79797979798 0 -2.0 1e-06 
0.555555555556 1.79797979798 0 -2.0 1e-06 
0.611111111111 1.79797979798 0 -2.0 1e-06 
0.666666666667 1.79797979798 0 -2.0 1e-06 
0.722222222222 1.79797979798 0 -2.0 1e-06 
0.777777777778 1.79797979798 0 -2.0 1e-06 
0.833333333333 1.79797979798 0 -2.0 1e-06 
0.888888888889 1.79797979798 0 -2.0 1e-06 
0.944444444444 1.79797979798 0 -2.0 1e-06 
1.0 1.79797979798 0 -2.0 1e-06 
0.5 1.83838383838 0 -2.0 1e-06 
0.555555555556 1.83838383838 0 -2.0 1e-06 
0.611111111111 1.83838383838 0 -2.0 1e-06 
0.666666666667 1.83838383838 0 -2.0 1e-06 
0.722222222222 1.83838383838 0 -2.0 1e-06 
0.777777777778 1.83838383838 0 -2.0 1e-06 
0.833333333333 1.83838383838 0 -2.0 1e-06 
0.888888888889 1.83838383838 0 -2.0 1e-06 
0.944444444444 1.83838383838 0 -2.0 1e-06 
1.0 1.83838383838 0 -2.0 1e-06 
0.5 1.87878787879 0 -2.0 1e-06 
0.555555555556 1.87878787879 0 -2.0 1e-06 
0.611111111111 1.87878787879 0 -2.0 1e-06 
0.666666666667 1.87878787879 0 -2.0 1e-06 
0.722222222222 1.87878787879 0 -2.0 1e-06 
0.777777777778 1.87878787879 0 -2.0 1e-06 
0.833333333333 1.87878787879 0 -2.0 1e-06 
0.888888888889 1.87878787879 0 -2.0 1e-06 
0.944444444444 1.87878787879 0 -2.0 1e-06 
1.0 1.87878787879 0 -2.0 1e-06 
0.5 1.91919191919 0 -2.0 1e-06 
0.555555555556 1.91919191919 0 -2.0 1e-06 
0.611111111111 1.91919191919 0 -2.0 1e-06 
0.666666666667 1.91919191919 0 -2.0 1e-06 
0.722222222222 1.91919191919 0 -2.0 1e-06 
0.777777777778 1.91919191919 0 -2.0 1e-06 
0.833333333333 1.91919191919 0 -2.0 1e-06 
0.888888888889 1.91919191919 0 -2.0 1e-06 
0.944444444444 1.91919191919 0 -2.0 1e-06 
1.0 1.91919191919 0 -2.0 1e-06 
0.5 1.9595959596 0 -2.0 1e-06 
0.555555555556 1.9595959596 0 -2.0 1e-06 
0.611111111111 1.9595959596 0 -2.0 1e-06 
0.666666666667 1.9595959596 0 -2.0 1e-06 
0.722222222222 1.9595959596 0 -2.0 1e-06 
0.777777777778 1.9595959596 0 -2.0 1e-06 
0.833333333333 1.9595959596 0 -2.0 1e-06 
0.888888888889 1.9595959596 0 -2.0 1e-06 
0.944444444444 1.9595959596 0 -2.0 1e-06 
1.0 1.9595959596 0 -2.0 1e-06 
0.5 2.0 0 -2.0 1e-06 
0.555555555556 2.0 0 -2.0 1e-06 
0.611111111111 2.0 0 -2.0 1e-06 
0.666666666667 2.0 0 -2.0 1e-06 
0.722222222222 2.0 0 -2.0 1e-06 
0.777777777778 2.0 0 -2.0 1e-06 
0.833333333333 2.0 0 -2.0 1e-06 
0.888888888889 2.0 0 -2.0 1e-06 
0.944444444444 2.0 0 -2.0 1e-06 
1.0 2.0 0 -2.0 1e-06 
0.5 -2.0 0 -1.6 1e-06 
0.555555555556 -2.0 0 -1.6 1e-06 
0.611111111111 -2.0 0 -1.6 1e-06 
0.666666666667 -2.0 0 -1.6 1e-06 
0.722222222222 -2.0 0 -1.6 1e-06 
0.777777777778 -2.0 0 -1.6 1e-06 
0.833333333333 -2.0 0 -1.6 1e-06 
0.888888888889 -2.0 0 -1.6 1e-06 
0.944444444444 -2.0 0 -1.6 1e-06 
1.0 -2.0 0 -1.6 1e-06 
0.5 -1.9595959596 0 -1.6 1e-06 
0.555555555556 -1.9595959596 0 -1.6 1e-06 
0.611111111111 -1.9595959596 0 -1.6 1e-06 
0.666666666667 -1.9595959596 0 -1.6 1e-06 
0.722222222222 -1.9595959596 0 -1.6 1e-06 
0.777777777778 -1.9595959596 0 -1.6 1e-06 
0.833333333333 -1.9595959596 0 -1.6 1e-06 
0.888888888889 -1.9595959596 0 -1.6 1e-06 
0.944444444444 -1.9595959596 0 -1.6 1e-06 
1.0 -1.9595959596 0 -1.6 1e-06 
0.5 -1.91919191919 0 -1.6 1e-06 
0.555555555556 -1.91919191919 0 -1.6 1e-06 
0.611111111111 -1.91919191919 0 -1.6 1e-06 
0.666666666667 -1.91919191919 0 -1.6 1e-06 
0.722222222222 -1.91919191919 0 -1.6 1e-06 
0.777777777778 -1.91919191919 0 -1.6 1e-06 
0.833333333333 -1.91919191919 0 -1.6 1e-06 
0.888888888889 -1.91919191919 0 -1.6 1e-06 
0.944444444444 -1.91919191919 0 -1.6 1e-06 
1.0 -1.91919191919 0 -1.6 1e-06 
0.5 -1.87878787879 0 -1.6 1e-06 
0.555555555556 -1.87878787879 0 -1.6 1e-06 
0.611111111111 -1.87878787879 0 -1.6 1e-06 
0.666666666667 -1.87878787879 0 -1.6 1e-06 
0.722222222222 -1.87878787879 0 -1.6 1e-06 
0.777777777778 -1.87878787879 0 -1.6 1e-06 
0.833333333333 -1.87878787879 0 -1.6 1e-06 
0.888888888889 -1.87878787879 0 -1.6 1e-06 
0.944444444444 -1.87878787879 0 -1.6 1e-06 
1.0 -1.87878787879 0 -1.6 1e-06 
0.5 -1.83838383838 0 -1.6 1e-06 
0.555555555556 -1.83838383838 0 -1.6 1e-06 
0.611111111111 -1.83838383838 0 -1.6 1e-06 
0.666666666667 -1.83838383838 0 -1.6 1e-06 
0.722222222222 -1.83838383838 0 -1.6 1e-06 
0.777777777778 -1.83838383838 0 -1.6 1e-06 
0.833333333333 -1.83838383838 0 -1.6 1e-06 
0.888888888889 -1.83838383838 0 -1.6 1e-06 
0.944444444444 -1.83838383838 0 -1.6 1e-06 
1.0 -1.83838383838 0 -1.6 1e-06 
0.5 -1.79797979798 0 -1.6 1e-06 
0.555555555556 -1.79797979798 0 -1.6 1e-06 
0.611111111111 -1.79797979798 0 -1.6 1e-06 
0.666666666667 -1.79797979798 0 -1.6 1e-06 
0.722222222222 -1.79797979798 0 -1.6 1e-06 
0.777777777778 -1.79797979798 0 -1.6 1e-06 
0.833333333333 -1.79797979798 0 -1.6 1e-06 
0.888888888889 -1.79797979798 0 -1.6 1e-06 
0.944444444444 -1.79797979798 0 -1.6 1e-06 
1.0 -1.79797979798 0 -1.6 1e-06 
0.5 -1.75757575758 0 -1.6 1e-06 
0.555555555556 -1.75757575758 0 -1.6 1e-06 
0.611111111111 -1.75757575758 0 -1.6 1e-06 
0.666666666667 -1.75757575758 0 -1.6 1e-06 
0.722222222222 -1.75757575758 0 -1.6 1e-06 
0.777777777778 -1.75757575758 0 -1.6 1e-06 
0.833333333333 -1.75757575758 0 -1.6 1e-06 
0.888888888889 -1.75757575758 0 -1.6 1e-06 
0.944444444444 -1.75757575758 0 -1.6 1e-06 
1.0 -1.75757575758 0 -1.6 1e-06 
0.5 -1.71717171717 0 -1.6 1e-06 
0.555555555556 -1.71717171717 0 -1.6 1e-06 
0.611111111111 -1.71717171717 0 -1.6 1e-06 
0.666666666667 -1.71717171717 0 -1.6 1e-06 
0.722222222222 -1.71717171717 0 -1.6 1e-06 
0.777777777778 -1.71717171717 0 -1.6 1e-06 
0.833333333333 -1.71717171717 0 -1.6 1e-06 
0.888888888889 -1.71717171717 0 -1.6 1e-06 
0.944444444444 -1.71717171717 0 -1.6 1e-06 
1.0 -1.71717171717 0 -1.6 1e-06 
0.5 -1.67676767677 0 -1.6 1e-06 
0.555555555556 -1.67676767677 0 -1.6 1e-06 
0.611111111111 -1.67676767677 0 -1.6 1e-06 
0.666666666667 -1.67676767677 0 -1.6 1e-06 
0.722222222222 -1.67676767677 0 -1.6 1e-06 
0.777777777778 -1.67676767677 0 -1.6 1e-06 
0.833333333333 -1.67676767677 0 -1.6 1e-06 
0.888888888889 -1.67676767677 0 -1.6 1e-06 
0.944444444444 -1.67676767677 0 -1.6 1e-06 
1.0 -1.67676767677 0 -1.6 1e-06 
0.5 -1.63636363636 0 -1.6 1e-06 
0.555555555556 -1.63636363636 0 -1.6 1e-06 
0.611111111111 -1.63636363636 0 -1.6 1e-06 
0.666666666667 -1.63636363636 0 -1.6 1e-06 
0.722222222222 -1.63636363636 0 -1.6 1e-06 
0.777777777778 -1.63636363636 0 -1.6 1e-06 
0.833333333333 -1.63636363636 0 -1.6 1e-06 
0.888888888889 -1.63636363636 0 -1.6 1e-06 
0.944444444444 -1.63636363636 0 -1.6 1e-06 
1.0 -1.63636363636 0 -1.6 1e-06 
0.5 -1.59595959596 0 -1.6 1e-06 
0.555555555556 -1.59595959596 0 -1.6 1e-06 
0.611111111111 -1.59595959596 0 -1.6 1e-06 
0.666666666667 -1.59595959596 0 -1.6 1e-06 
0.722222222222 -1.59595959596 0 -1.6 1e-06 
0.777777777778 -1.59595959596 0 -1.6 1e-06 
0.833333333333 -1.59595959596 0 -1.6 1e-06 
0.888888888889 -1.59595959596 0 -1.6 1e-06 
0.944444444444 -1.59595959596 0 -1.6 1e-06 
1.0 -1.59595959596 0 -1.6 1e-06 
0.5 -1.55555555556 0 -1.6 1e-06 
0.555555555556 -1.55555555556 0 -1.6 1e-06 
0.611111111111 -1.55555555556 0 -1.6 1e-06 
0.666666666667 -1.55555555556 0 -1.6 1e-06 
0.722222222222 -1.55555555556 0 -1.6 1e-06 
0.777777777778 -1.55555555556 0 -1.6 1e-06 
0.833333333333 -1.55555555556 0 -1.6 1e-06 
0.888888888889 -1.55555555556 0 -1.6 1e-06 
0.944444444444 -1.55555555556 0 -1.6 1e-06 
1.0 -1.55555555556 0 -1.6 1e-06 
0.5 -1.51515151515 0 -1.6 1e-06 
0.555555555556 -1.51515151515 0 -1.6 1e-06 
0.611111111111 -1.51515151515 0 -1.6 1e-06 
0.666666666667 -1.51515151515 0 -1.6 1e-06 
0.722222222222 -1.51515151515 0 -1.6 1e-06 
0.777777777778 -1.51515151515 0 -1.6 1e-06 
0.833333333333 -1.51515151515 0 -1.6 1e-06 
0.888888888889 -1.51515151515 0 -1.6 1e-06 
0.944444444444 -1.51515151515 0 -1.6 1e-06 
1.0 -1.51515151515 0 -1.6 1e-06 
0.5 -1.47474747475 0 -1.6 1e-06 
0.555555555556 -1.47474747475 0 -1.6 1e-06 
0.611111111111 -1.47474747475 0 -1.6 1e-06 
0.666666666667 -1.47474747475 0 -1.6 1e-06 
0.722222222222 -1.47474747475 0 -1.6 1e-06 
0.777777777778 -1.47474747475 0 -1.6 1e-06 
0.833333333333 -1.47474747475 0 -1.6 1e-06 
0.888888888889 -1.47474747475 0 -1.6 1e-06 
0.944444444444 -1.47474747475 0 -1.6 1e-06 
1.0 -1.47474747475 0 -1.6 1e-06 
0.5 -1.43434343434 0 -1.6 1e-06 
0.555555555556 -1.43434343434 0 -1.6 1e-06 
0.611111111111 -1.43434343434 0 -1.6 1e-06 
0.666666666667 -1.43434343434 0 -1.6 1e-06 
0.722222222222 -1.43434343434 0 -1.6 1e-06 
0.777777777778 -1.43434343434 0 -1.6 1e-06 
0.833333333333 -1.43434343434 0 -1.6 1e-06 
0.888888888889 -1.43434343434 0 -1.6 1e-06 
0.944444444444 -1.43434343434 0 -1.6 1e-06 
1.0 -1.43434343434 0 -1.6 1e-06 
0.5 -1.39393939394 0 -1.6 1e-06 
0.555555555556 -1.39393939394 0 -1.6 1e-06 
0.611111111111 -1.39393939394 0 -1.6 1e-06 
0.666666666667 -1.39393939394 0 -1.6 1e-06 
0.722222222222 -1.39393939394 0 -1.6 1e-06 
0.777777777778 -1.39393939394 0 -1.6 1e-06 
0.833333333333 -1.39393939394 0 -1.6 1e-06 
0.888888888889 -1.39393939394 0 -1.6 1e-06 
0.944444444444 -1.39393939394 0 -1.6 1e-06 
1.0 -1.39393939394 0 -1.6 1e-06 
0.5 -1.35353535354 0 -1.6 1e-06 
0.555555555556 -1.35353535354 0 -1.6 1e-06 
0.611111111111 -1.35353535354 0 -1.6 1e-06 
0.666666666667 -1.35353535354 0 -1.6 1e-06 
0.722222222222 -1.35353535354 0 -1.6 1e-06 
0.777777777778 -1.35353535354 0 -1.6 1e-06 
0.833333333333 -1.35353535354 0 -1.6 1e-06 
0.888888888889 -1.35353535354 0 -1.6 1e-06 
0.944444444444 -1.35353535354 0 -1.6 1e-06 
1.0 -1.35353535354 0 -1.6 1e-06 
0.5 -1.31313131313 0 -1.6 1e-06 
0.555555555556 -1.31313131313 0 -1.6 1e-06 
0.611111111111 -1.31313131313 0 -1.6 1e-06 
0.666666666667 -1.31313131313 0 -1.6 1e-06 
0.722222222222 -1.31313131313 0 -1.6 1e-06 
0.777777777778 -1.31313131313 0 -1.6 1e-06 
0.833333333333 -1.31313131313 0 -1.6 1e-06 
0.888888888889 -1.31313131313 0 -1.6 1e-06 
0.944444444444 -1.31313131313 0 -1.6 1e-06 
1.0 -1.31313131313 0 -1.6 1e-06 
0.5 -1.27272727273 0 -1.6 1e-06 
0.555555555556 -1.27272727273 0 -1.6 1e-06 
0.611111111111 -1.27272727273 0 -1.6 1e-06 
0.666666666667 -1.27272727273 0 -1.6 1e-06 
0.722222222222 -1.27272727273 0 -1.6 1e-06 
0.777777777778 -1.27272727273 0 -1.6 1e-06 
0.833333333333 -1.27272727273 0 -1.6 1e-06 
0.888888888889 -1.27272727273 0 -1.6 1e-06 
0.944444444444 -1.27272727273 0 -1.6 1e-06 
1.0 -1.27272727273 0 -1.6 1e-06 
0.5 -1.23232323232 0 -1.6 1e-06 
0.555555555556 -1.23232323232 0 -1.6 1e-06 
0.611111111111 -1.23232323232 0 -1.6 1e-06 
0.666666666667 -1.23232323232 0 -1.6 1e-06 
0.722222222222 -1.23232323232 0 -1.6 1e-06 
0.777777777778 -1.23232323232 0 -1.6 1e-06 
0.833333333333 -1.23232323232 0 -1.6 1e-06 
0.888888888889 -1.23232323232 0 -1.6 1e-06 
0.944444444444 -1.23232323232 0 -1.6 1e-06 
1.0 -1.23232323232 0 -1.6 1e-06 
0.5 -1.19191919192 0 -1.6 1e-06 
0.555555555556 -1.19191919192 0 -1.6 1e-06 
0.611111111111 -1.19191919192 0 -1.6 1e-06 
0.666666666667 -1.19191919192 0 -1.6 1e-06 
0.722222222222 -1.19191919192 0 -1.6 1e-06 
0.777777777778 -1.19191919192 0 -1.6 1e-06 
0.833333333333 -1.19191919192 0 -1.6 1e-06 
0.888888888889 -1.19191919192 0 -1.6 1e-06 
0.944444444444 -1.19191919192 0 -1.6 1e-06 
1.0 -1.19191919192 0 -1.6 1e-06 
0.5 -1.15151515152 0 -1.6 1e-06 
0.555555555556 -1.15151515152 0 -1.6 1e-06 
0.611111111111 -1.15151515152 0 -1.6 1e-06 
0.666666666667 -1.15151515152 0 -1.6 1e-06 
0.722222222222 -1.15151515152 0 -1.6 1e-06 
0.777777777778 -1.15151515152 0 -1.6 1e-06 
0.833333333333 -1.15151515152 0 -1.6 1e-06 
0.888888888889 -1.15151515152 0 -1.6 1e-06 
0.944444444444 -1.15151515152 0 -1.6 1e-06 
1.0 -1.15151515152 0 -1.6 1e-06 
0.5 -1.11111111111 0 -1.6 1e-06 
0.555555555556 -1.11111111111 0 -1.6 1e-06 
0.611111111111 -1.11111111111 0 -1.6 1e-06 
0.666666666667 -1.11111111111 0 -1.6 1e-06 
0.722222222222 -1.11111111111 0 -1.6 1e-06 
0.777777777778 -1.11111111111 0 -1.6 1e-06 
0.833333333333 -1.11111111111 0 -1.6 1e-06 
0.888888888889 -1.11111111111 0 -1.6 1e-06 
0.944444444444 -1.11111111111 0 -1.6 1e-06 
1.0 -1.11111111111 0 -1.6 1e-06 
0.5 -1.07070707071 0 -1.6 1e-06 
0.555555555556 -1.07070707071 0 -1.6 1e-06 
0.611111111111 -1.07070707071 0 -1.6 1e-06 
0.666666666667 -1.07070707071 0 -1.6 1e-06 
0.722222222222 -1.07070707071 0 -1.6 1e-06 
0.777777777778 -1.07070707071 0 -1.6 1e-06 
0.833333333333 -1.07070707071 0 -1.6 1e-06 
0.888888888889 -1.07070707071 0 -1.6 1e-06 
0.944444444444 -1.07070707071 0 -1.6 1e-06 
1.0 -1.07070707071 0 -1.6 1e-06 
0.5 -1.0303030303 0 -1.6 1e-06 
0.555555555556 -1.0303030303 0 -1.6 1e-06 
0.611111111111 -1.0303030303 0 -1.6 1e-06 
0.666666666667 -1.0303030303 0 -1.6 1e-06 
0.722222222222 -1.0303030303 0 -1.6 1e-06 
0.777777777778 -1.0303030303 0 -1.6 1e-06 
0.833333333333 -1.0303030303 0 -1.6 1e-06 
0.888888888889 -1.0303030303 0 -1.6 1e-06 
0.944444444444 -1.0303030303 0 -1.6 1e-06 
1.0 -1.0303030303 0 -1.6 1e-06 
0.5 -0.989898989899 0 -1.6 1e-06 
0.555555555556 -0.989898989899 0 -1.6 1e-06 
0.611111111111 -0.989898989899 0 -1.6 1e-06 
0.666666666667 -0.989898989899 0 -1.6 1e-06 
0.722222222222 -0.989898989899 0 -1.6 1e-06 
0.777777777778 -0.989898989899 0 -1.6 1e-06 
0.833333333333 -0.989898989899 0 -1.6 1e-06 
0.888888888889 -0.989898989899 0 -1.6 1e-06 
0.944444444444 -0.989898989899 0 -1.6 1e-06 
1.0 -0.989898989899 0 -1.6 1e-06 
0.5 -0.949494949495 0 -1.6 1e-06 
0.555555555556 -0.949494949495 0 -1.6 1e-06 
0.611111111111 -0.949494949495 0 -1.6 1e-06 
0.666666666667 -0.949494949495 0 -1.6 1e-06 
0.722222222222 -0.949494949495 0 -1.6 1e-06 
0.777777777778 -0.949494949495 0 -1.6 1e-06 
0.833333333333 -0.949494949495 0 -1.6 1e-06 
0.888888888889 -0.949494949495 0 -1.6 1e-06 
0.944444444444 -0.949494949495 0 -1.6 1e-06 
1.0 -0.949494949495 0 -1.6 1e-06 
0.5 -0.909090909091 0 -1.6 1e-06 
0.555555555556 -0.909090909091 0 -1.6 1e-06 
0.611111111111 -0.909090909091 0 -1.6 1e-06 
0.666666666667 -0.909090909091 0 -1.6 1e-06 
0.722222222222 -0.909090909091 0 -1.6 1e-06 
0.777777777778 -0.909090909091 0 -1.6 1e-06 
0.833333333333 -0.909090909091 0 -1.6 1e-06 
0.888888888889 -0.909090909091 0 -1.6 1e-06 
0.944444444444 -0.909090909091 0 -1.6 1e-06 
1.0 -0.909090909091 0 -1.6 1e-06 
0.5 -0.868686868687 0 -1.6 1e-06 
0.555555555556 -0.868686868687 0 -1.6 1e-06 
0.611111111111 -0.868686868687 0 -1.6 1e-06 
0.666666666667 -0.868686868687 0 -1.6 1e-06 
0.722222222222 -0.868686868687 0 -1.6 1e-06 
0.777777777778 -0.868686868687 0 -1.6 1e-06 
0.833333333333 -0.868686868687 0 -1.6 1e-06 
0.888888888889 -0.868686868687 0 -1.6 1e-06 
0.944444444444 -0.868686868687 0 -1.6 1e-06 
1.0 -0.868686868687 0 -1.6 1e-06 
0.5 -0.828282828283 0 -1.6 1e-06 
0.555555555556 -0.828282828283 0 -1.6 1e-06 
0.611111111111 -0.828282828283 0 -1.6 1e-06 
0.666666666667 -0.828282828283 0 -1.6 1e-06 
0.722222222222 -0.828282828283 0 -1.6 1e-06 
0.777777777778 -0.828282828283 0 -1.6 1e-06 
0.833333333333 -0.828282828283 0 -1.6 1e-06 
0.888888888889 -0.828282828283 0 -1.6 1e-06 
0.944444444444 -0.828282828283 0 -1.6 1e-06 
1.0 -0.828282828283 0 -1.6 1e-06 
0.5 -0.787878787879 0 -1.6 1e-06 
0.555555555556 -0.787878787879 0 -1.6 1e-06 
0.611111111111 -0.787878787879 0 -1.6 1e-06 
0.666666666667 -0.787878787879 0 -1.6 1e-06 
0.722222222222 -0.787878787879 0 -1.6 1e-06 
0.777777777778 -0.787878787879 0 -1.6 1e-06 
0.833333333333 -0.787878787879 0 -1.6 1e-06 
0.888888888889 -0.787878787879 0 -1.6 1e-06 
0.944444444444 -0.787878787879 0 -1.6 1e-06 
1.0 -0.787878787879 0 -1.6 1e-06 
0.5 -0.747474747475 0 -1.6 1e-06 
0.555555555556 -0.747474747475 0 -1.6 1e-06 
0.611111111111 -0.747474747475 0 -1.6 1e-06 
0.666666666667 -0.747474747475 0 -1.6 1e-06 
0.722222222222 -0.747474747475 0 -1.6 1e-06 
0.777777777778 -0.747474747475 0 -1.6 1e-06 
0.833333333333 -0.747474747475 0 -1.6 1e-06 
0.888888888889 -0.747474747475 0 -1.6 1e-06 
0.944444444444 -0.747474747475 0 -1.6 1e-06 
1.0 -0.747474747475 0 -1.6 1e-06 
0.5 -0.707070707071 0 -1.6 1e-06 
0.555555555556 -0.707070707071 0 -1.6 1e-06 
0.611111111111 -0.707070707071 0 -1.6 1e-06 
0.666666666667 -0.707070707071 0 -1.6 1e-06 
0.722222222222 -0.707070707071 0 -1.6 1e-06 
0.777777777778 -0.707070707071 0 -1.6 1e-06 
0.833333333333 -0.707070707071 0 -1.6 1e-06 
0.888888888889 -0.707070707071 0 -1.6 1e-06 
0.944444444444 -0.707070707071 0 -1.6 1e-06 
1.0 -0.707070707071 0 -1.6 1e-06 
0.5 -0.666666666667 0 -1.6 1e-06 
0.555555555556 -0.666666666667 0 -1.6 1e-06 
0.611111111111 -0.666666666667 0 -1.6 1e-06 
0.666666666667 -0.666666666667 0 -1.6 1e-06 
0.722222222222 -0.666666666667 0 -1.6 1e-06 
0.777777777778 -0.666666666667 0 -1.6 1e-06 
0.833333333333 -0.666666666667 0 -1.6 1e-06 
0.888888888889 -0.666666666667 0 -1.6 1e-06 
0.944444444444 -0.666666666667 0 -1.6 1e-06 
1.0 -0.666666666667 0 -1.6 1e-06 
0.5 -0.626262626263 0 -1.6 1e-06 
0.555555555556 -0.626262626263 0 -1.6 1e-06 
0.611111111111 -0.626262626263 0 -1.6 1e-06 
0.666666666667 -0.626262626263 0 -1.6 1e-06 
0.722222222222 -0.626262626263 0 -1.6 1e-06 
0.777777777778 -0.626262626263 0 -1.6 1e-06 
0.833333333333 -0.626262626263 0 -1.6 1e-06 
0.888888888889 -0.626262626263 0 -1.6 1e-06 
0.944444444444 -0.626262626263 0 -1.6 1e-06 
1.0 -0.626262626263 0 -1.6 1e-06 
0.5 -0.585858585859 0 -1.6 1e-06 
0.555555555556 -0.585858585859 0 -1.6 1e-06 
0.611111111111 -0.585858585859 0 -1.6 1e-06 
0.666666666667 -0.585858585859 0 -1.6 1e-06 
0.722222222222 -0.585858585859 0 -1.6 1e-06 
0.777777777778 -0.585858585859 0 -1.6 1e-06 
0.833333333333 -0.585858585859 0 -1.6 1e-06 
0.888888888889 -0.585858585859 0 -1.6 1e-06 
0.944444444444 -0.585858585859 0 -1.6 1e-06 
1.0 -0.585858585859 0 -1.6 1e-06 
0.5 -0.545454545455 0 -1.6 1e-06 
0.555555555556 -0.545454545455 0 -1.6 1e-06 
0.611111111111 -0.545454545455 0 -1.6 1e-06 
0.666666666667 -0.545454545455 0 -1.6 1e-06 
0.722222222222 -0.545454545455 0 -1.6 1e-06 
0.777777777778 -0.545454545455 0 -1.6 1e-06 
0.833333333333 -0.545454545455 0 -1.6 1e-06 
0.888888888889 -0.545454545455 0 -1.6 1e-06 
0.944444444444 -0.545454545455 0 -1.6 1e-06 
1.0 -0.545454545455 0 -1.6 1e-06 
0.5 -0.505050505051 0 -1.6 1e-06 
0.555555555556 -0.505050505051 0 -1.6 1e-06 
0.611111111111 -0.505050505051 0 -1.6 1e-06 
0.666666666667 -0.505050505051 0 -1.6 1e-06 
0.722222222222 -0.505050505051 0 -1.6 1e-06 
0.777777777778 -0.505050505051 0 -1.6 1e-06 
0.833333333333 -0.505050505051 0 -1.6 1e-06 
0.888888888889 -0.505050505051 0 -1.6 1e-06 
0.944444444444 -0.505050505051 0 -1.6 1e-06 
1.0 -0.505050505051 0 -1.6 1e-06 
0.5 -0.464646464646 0 -1.6 1e-06 
0.555555555556 -0.464646464646 0 -1.6 1e-06 
0.611111111111 -0.464646464646 0 -1.6 1e-06 
0.666666666667 -0.464646464646 0 -1.6 1e-06 
0.722222222222 -0.464646464646 0 -1.6 1e-06 
0.777777777778 -0.464646464646 0 -1.6 1e-06 
0.833333333333 -0.464646464646 0 -1.6 1e-06 
0.888888888889 -0.464646464646 0 -1.6 1e-06 
0.944444444444 -0.464646464646 0 -1.6 1e-06 
1.0 -0.464646464646 0 -1.6 1e-06 
0.5 -0.424242424242 0 -1.6 1e-06 
0.555555555556 -0.424242424242 0 -1.6 1e-06 
0.611111111111 -0.424242424242 0 -1.6 1e-06 
0.666666666667 -0.424242424242 0 -1.6 1e-06 
0.722222222222 -0.424242424242 0 -1.6 1e-06 
0.777777777778 -0.424242424242 0 -1.6 1e-06 
0.833333333333 -0.424242424242 0 -1.6 1e-06 
0.888888888889 -0.424242424242 0 -1.6 1e-06 
0.944444444444 -0.424242424242 0 -1.6 1e-06 
1.0 -0.424242424242 0 -1.6 1e-06 
0.5 -0.383838383838 0 -1.6 1e-06 
0.555555555556 -0.383838383838 0 -1.6 1e-06 
0.611111111111 -0.383838383838 0 -1.6 1e-06 
0.666666666667 -0.383838383838 0 -1.6 1e-06 
0.722222222222 -0.383838383838 0 -1.6 1e-06 
0.777777777778 -0.383838383838 0 -1.6 1e-06 
0.833333333333 -0.383838383838 0 -1.6 1e-06 
0.888888888889 -0.383838383838 0 -1.6 1e-06 
0.944444444444 -0.383838383838 0 -1.6 1e-06 
1.0 -0.383838383838 0 -1.6 1e-06 
0.5 -0.343434343434 0 -1.6 1e-06 
0.555555555556 -0.343434343434 0 -1.6 1e-06 
0.611111111111 -0.343434343434 0 -1.6 1e-06 
0.666666666667 -0.343434343434 0 -1.6 1e-06 
0.722222222222 -0.343434343434 0 -1.6 1e-06 
0.777777777778 -0.343434343434 0 -1.6 1e-06 
0.833333333333 -0.343434343434 0 -1.6 1e-06 
0.888888888889 -0.343434343434 0 -1.6 1e-06 
0.944444444444 -0.343434343434 0 -1.6 1e-06 
1.0 -0.343434343434 0 -1.6 1e-06 
0.5 -0.30303030303 0 -1.6 1e-06 
0.555555555556 -0.30303030303 0 -1.6 1e-06 
0.611111111111 -0.30303030303 0 -1.6 1e-06 
0.666666666667 -0.30303030303 0 -1.6 1e-06 
0.722222222222 -0.30303030303 0 -1.6 1e-06 
0.777777777778 -0.30303030303 0 -1.6 1e-06 
0.833333333333 -0.30303030303 0 -1.6 1e-06 
0.888888888889 -0.30303030303 0 -1.6 1e-06 
0.944444444444 -0.30303030303 0 -1.6 1e-06 
1.0 -0.30303030303 0 -1.6 1e-06 
0.5 -0.262626262626 0 -1.6 1e-06 
0.555555555556 -0.262626262626 0 -1.6 1e-06 
0.611111111111 -0.262626262626 0 -1.6 1e-06 
0.666666666667 -0.262626262626 0 -1.6 1e-06 
0.722222222222 -0.262626262626 0 -1.6 1e-06 
0.777777777778 -0.262626262626 0 -1.6 1e-06 
0.833333333333 -0.262626262626 0 -1.6 1e-06 
0.888888888889 -0.262626262626 0 -1.6 1e-06 
0.944444444444 -0.262626262626 0 -1.6 1e-06 
1.0 -0.262626262626 0 -1.6 1e-06 
0.5 -0.222222222222 0 -1.6 1e-06 
0.555555555556 -0.222222222222 0 -1.6 1e-06 
0.611111111111 -0.222222222222 0 -1.6 1e-06 
0.666666666667 -0.222222222222 0 -1.6 1e-06 
0.722222222222 -0.222222222222 0 -1.6 1e-06 
0.777777777778 -0.222222222222 0 -1.6 1e-06 
0.833333333333 -0.222222222222 0 -1.6 1e-06 
0.888888888889 -0.222222222222 0 -1.6 1e-06 
0.944444444444 -0.222222222222 0 -1.6 1e-06 
1.0 -0.222222222222 0 -1.6 1e-06 
0.5 -0.181818181818 0 -1.6 1e-06 
0.555555555556 -0.181818181818 0 -1.6 1e-06 
0.611111111111 -0.181818181818 0 -1.6 1e-06 
0.666666666667 -0.181818181818 0 -1.6 1e-06 
0.722222222222 -0.181818181818 0 -1.6 1e-06 
0.777777777778 -0.181818181818 0 -1.6 1e-06 
0.833333333333 -0.181818181818 0 -1.6 1e-06 
0.888888888889 -0.181818181818 0 -1.6 1e-06 
0.944444444444 -0.181818181818 0 -1.6 1e-06 
1.0 -0.181818181818 0 -1.6 1e-06 
0.5 -0.141414141414 0 -1.6 1e-06 
0.555555555556 -0.141414141414 0 -1.6 1e-06 
0.611111111111 -0.141414141414 0 -1.6 1e-06 
0.666666666667 -0.141414141414 0 -1.6 1e-06 
0.722222222222 -0.141414141414 0 -1.6 1e-06 
0.777777777778 -0.141414141414 0 -1.6 1e-06 
0.833333333333 -0.141414141414 0 -1.6 1e-06 
0.888888888889 -0.141414141414 0 -1.6 1e-06 
0.944444444444 -0.141414141414 0 -1.6 1e-06 
1.0 -0.141414141414 0 -1.6 1e-06 
0.5 -0.10101010101 0 -1.6 1e-06 
0.555555555556 -0.10101010101 0 -1.6 1e-06 
0.611111111111 -0.10101010101 0 -1.6 1e-06 
0.666666666667 -0.10101010101 0 -1.6 1e-06 
0.722222222222 -0.10101010101 0 -1.6 1e-06 
0.777777777778 -0.10101010101 0 -1.6 1e-06 
0.833333333333 -0.10101010101 0 -1.6 1e-06 
0.888888888889 -0.10101010101 0 -1.6 1e-06 
0.944444444444 -0.10101010101 0 -1.6 1e-06 
1.0 -0.10101010101 0 -1.6 1e-06 
0.5 -0.0606060606061 0 -1.6 1e-06 
0.555555555556 -0.0606060606061 0 -1.6 1e-06 
0.611111111111 -0.0606060606061 0 -1.6 1e-06 
0.666666666667 -0.0606060606061 0 -1.6 1e-06 
0.722222222222 -0.0606060606061 0 -1.6 1e-06 
0.777777777778 -0.0606060606061 0 -1.6 1e-06 
0.833333333333 -0.0606060606061 0 -1.6 1e-06 
0.888888888889 -0.0606060606061 0 -1.6 1e-06 
0.944444444444 -0.0606060606061 0 -1.6 1e-06 
1.0 -0.0606060606061 0 -1.6 1e-06 
0.5 -0.020202020202 0 -1.6 1e-06 
0.555555555556 -0.020202020202 0 -1.6 1e-06 
0.611111111111 -0.020202020202 0 -1.6 1e-06 
0.666666666667 -0.020202020202 0 -1.6 1e-06 
0.722222222222 -0.020202020202 0 -1.6 1e-06 
0.777777777778 -0.020202020202 0 -1.6 1e-06 
0.833333333333 -0.020202020202 0 -1.6 1e-06 
0.888888888889 -0.020202020202 0 -1.6 1e-06 
0.944444444444 -0.020202020202 0 -1.6 1e-06 
1.0 -0.020202020202 0 -1.6 1e-06 
0.5 0.020202020202 0 -1.6 1e-06 
0.555555555556 0.020202020202 0 -1.6 1e-06 
0.611111111111 0.020202020202 0 -1.6 1e-06 
0.666666666667 0.020202020202 0 -1.6 1e-06 
0.722222222222 0.020202020202 0 -1.6 1e-06 
0.777777777778 0.020202020202 0 -1.6 1e-06 
0.833333333333 0.020202020202 0 -1.6 1e-06 
0.888888888889 0.020202020202 0 -1.6 1e-06 
0.944444444444 0.020202020202 0 -1.6 1e-06 
1.0 0.020202020202 0 -1.6 1e-06 
0.5 0.0606060606061 0 -1.6 1e-06 
0.555555555556 0.0606060606061 0 -1.6 1e-06 
0.611111111111 0.0606060606061 0 -1.6 1e-06 
0.666666666667 0.0606060606061 0 -1.6 1e-06 
0.722222222222 0.0606060606061 0 -1.6 1e-06 
0.777777777778 0.0606060606061 0 -1.6 1e-06 
0.833333333333 0.0606060606061 0 -1.6 1e-06 
0.888888888889 0.0606060606061 0 -1.6 1e-06 
0.944444444444 0.0606060606061 0 -1.6 1e-06 
1.0 0.0606060606061 0 -1.6 1e-06 
0.5 0.10101010101 0 -1.6 1e-06 
0.555555555556 0.10101010101 0 -1.6 1e-06 
0.611111111111 0.10101010101 0 -1.6 1e-06 
0.666666666667 0.10101010101 0 -1.6 1e-06 
0.722222222222 0.10101010101 0 -1.6 1e-06 
0.777777777778 0.10101010101 0 -1.6 1e-06 
0.833333333333 0.10101010101 0 -1.6 1e-06 
0.888888888889 0.10101010101 0 -1.6 1e-06 
0.944444444444 0.10101010101 0 -1.6 1e-06 
1.0 0.10101010101 0 -1.6 1e-06 
0.5 0.141414141414 0 -1.6 1e-06 
0.555555555556 0.141414141414 0 -1.6 1e-06 
0.611111111111 0.141414141414 0 -1.6 1e-06 
0.666666666667 0.141414141414 0 -1.6 1e-06 
0.722222222222 0.141414141414 0 -1.6 1e-06 
0.777777777778 0.141414141414 0 -1.6 1e-06 
0.833333333333 0.141414141414 0 -1.6 1e-06 
0.888888888889 0.141414141414 0 -1.6 1e-06 
0.944444444444 0.141414141414 0 -1.6 1e-06 
1.0 0.141414141414 0 -1.6 1e-06 
0.5 0.181818181818 0 -1.6 1e-06 
0.555555555556 0.181818181818 0 -1.6 1e-06 
0.611111111111 0.181818181818 0 -1.6 1e-06 
0.666666666667 0.181818181818 0 -1.6 1e-06 
0.722222222222 0.181818181818 0 -1.6 1e-06 
0.777777777778 0.181818181818 0 -1.6 1e-06 
0.833333333333 0.181818181818 0 -1.6 1e-06 
0.888888888889 0.181818181818 0 -1.6 1e-06 
0.944444444444 0.181818181818 0 -1.6 1e-06 
1.0 0.181818181818 0 -1.6 1e-06 
0.5 0.222222222222 0 -1.6 1e-06 
0.555555555556 0.222222222222 0 -1.6 1e-06 
0.611111111111 0.222222222222 0 -1.6 1e-06 
0.666666666667 0.222222222222 0 -1.6 1e-06 
0.722222222222 0.222222222222 0 -1.6 1e-06 
0.777777777778 0.222222222222 0 -1.6 1e-06 
0.833333333333 0.222222222222 0 -1.6 1e-06 
0.888888888889 0.222222222222 0 -1.6 1e-06 
0.944444444444 0.222222222222 0 -1.6 1e-06 
1.0 0.222222222222 0 -1.6 1e-06 
0.5 0.262626262626 0 -1.6 1e-06 
0.555555555556 0.262626262626 0 -1.6 1e-06 
0.611111111111 0.262626262626 0 -1.6 1e-06 
0.666666666667 0.262626262626 0 -1.6 1e-06 
0.722222222222 0.262626262626 0 -1.6 1e-06 
0.777777777778 0.262626262626 0 -1.6 1e-06 
0.833333333333 0.262626262626 0 -1.6 1e-06 
0.888888888889 0.262626262626 0 -1.6 1e-06 
0.944444444444 0.262626262626 0 -1.6 1e-06 
1.0 0.262626262626 0 -1.6 1e-06 
0.5 0.30303030303 0 -1.6 1e-06 
0.555555555556 0.30303030303 0 -1.6 1e-06 
0.611111111111 0.30303030303 0 -1.6 1e-06 
0.666666666667 0.30303030303 0 -1.6 1e-06 
0.722222222222 0.30303030303 0 -1.6 1e-06 
0.777777777778 0.30303030303 0 -1.6 1e-06 
0.833333333333 0.30303030303 0 -1.6 1e-06 
0.888888888889 0.30303030303 0 -1.6 1e-06 
0.944444444444 0.30303030303 0 -1.6 1e-06 
1.0 0.30303030303 0 -1.6 1e-06 
0.5 0.343434343434 0 -1.6 1e-06 
0.555555555556 0.343434343434 0 -1.6 1e-06 
0.611111111111 0.343434343434 0 -1.6 1e-06 
0.666666666667 0.343434343434 0 -1.6 1e-06 
0.722222222222 0.343434343434 0 -1.6 1e-06 
0.777777777778 0.343434343434 0 -1.6 1e-06 
0.833333333333 0.343434343434 0 -1.6 1e-06 
0.888888888889 0.343434343434 0 -1.6 1e-06 
0.944444444444 0.343434343434 0 -1.6 1e-06 
1.0 0.343434343434 0 -1.6 1e-06 
0.5 0.383838383838 0 -1.6 1e-06 
0.555555555556 0.383838383838 0 -1.6 1e-06 
0.611111111111 0.383838383838 0 -1.6 1e-06 
0.666666666667 0.383838383838 0 -1.6 1e-06 
0.722222222222 0.383838383838 0 -1.6 1e-06 
0.777777777778 0.383838383838 0 -1.6 1e-06 
0.833333333333 0.383838383838 0 -1.6 1e-06 
0.888888888889 0.383838383838 0 -1.6 1e-06 
0.944444444444 0.383838383838 0 -1.6 1e-06 
1.0 0.383838383838 0 -1.6 1e-06 
0.5 0.424242424242 0 -1.6 1e-06 
0.555555555556 0.424242424242 0 -1.6 1e-06 
0.611111111111 0.424242424242 0 -1.6 1e-06 
0.666666666667 0.424242424242 0 -1.6 1e-06 
0.722222222222 0.424242424242 0 -1.6 1e-06 
0.777777777778 0.424242424242 0 -1.6 1e-06 
0.833333333333 0.424242424242 0 -1.6 1e-06 
0.888888888889 0.424242424242 0 -1.6 1e-06 
0.944444444444 0.424242424242 0 -1.6 1e-06 
1.0 0.424242424242 0 -1.6 1e-06 
0.5 0.464646464646 0 -1.6 1e-06 
0.555555555556 0.464646464646 0 -1.6 1e-06 
0.611111111111 0.464646464646 0 -1.6 1e-06 
0.666666666667 0.464646464646 0 -1.6 1e-06 
0.722222222222 0.464646464646 0 -1.6 1e-06 
0.777777777778 0.464646464646 0 -1.6 1e-06 
0.833333333333 0.464646464646 0 -1.6 1e-06 
0.888888888889 0.464646464646 0 -1.6 1e-06 
0.944444444444 0.464646464646 0 -1.6 1e-06 
1.0 0.464646464646 0 -1.6 1e-06 
0.5 0.505050505051 0 -1.6 1e-06 
0.555555555556 0.505050505051 0 -1.6 1e-06 
0.611111111111 0.505050505051 0 -1.6 1e-06 
0.666666666667 0.505050505051 0 -1.6 1e-06 
0.722222222222 0.505050505051 0 -1.6 1e-06 
0.777777777778 0.505050505051 0 -1.6 1e-06 
0.833333333333 0.505050505051 0 -1.6 1e-06 
0.888888888889 0.505050505051 0 -1.6 1e-06 
0.944444444444 0.505050505051 0 -1.6 1e-06 
1.0 0.505050505051 0 -1.6 1e-06 
0.5 0.545454545455 0 -1.6 1e-06 
0.555555555556 0.545454545455 0 -1.6 1e-06 
0.611111111111 0.545454545455 0 -1.6 1e-06 
0.666666666667 0.545454545455 0 -1.6 1e-06 
0.722222222222 0.545454545455 0 -1.6 1e-06 
0.777777777778 0.545454545455 0 -1.6 1e-06 
0.833333333333 0.545454545455 0 -1.6 1e-06 
0.888888888889 0.545454545455 0 -1.6 1e-06 
0.944444444444 0.545454545455 0 -1.6 1e-06 
1.0 0.545454545455 0 -1.6 1e-06 
0.5 0.585858585859 0 -1.6 1e-06 
0.555555555556 0.585858585859 0 -1.6 1e-06 
0.611111111111 0.585858585859 0 -1.6 1e-06 
0.666666666667 0.585858585859 0 -1.6 1e-06 
0.722222222222 0.585858585859 0 -1.6 1e-06 
0.777777777778 0.585858585859 0 -1.6 1e-06 
0.833333333333 0.585858585859 0 -1.6 1e-06 
0.888888888889 0.585858585859 0 -1.6 1e-06 
0.944444444444 0.585858585859 0 -1.6 1e-06 
1.0 0.585858585859 0 -1.6 1e-06 
0.5 0.626262626263 0 -1.6 1e-06 
0.555555555556 0.626262626263 0 -1.6 1e-06 
0.611111111111 0.626262626263 0 -1.6 1e-06 
0.666666666667 0.626262626263 0 -1.6 1e-06 
0.722222222222 0.626262626263 0 -1.6 1e-06 
0.777777777778 0.626262626263 0 -1.6 1e-06 
0.833333333333 0.626262626263 0 -1.6 1e-06 
0.888888888889 0.626262626263 0 -1.6 1e-06 
0.944444444444 0.626262626263 0 -1.6 1e-06 
1.0 0.626262626263 0 -1.6 1e-06 
0.5 0.666666666667 0 -1.6 1e-06 
0.555555555556 0.666666666667 0 -1.6 1e-06 
0.611111111111 0.666666666667 0 -1.6 1e-06 
0.666666666667 0.666666666667 0 -1.6 1e-06 
0.722222222222 0.666666666667 0 -1.6 1e-06 
0.777777777778 0.666666666667 0 -1.6 1e-06 
0.833333333333 0.666666666667 0 -1.6 1e-06 
0.888888888889 0.666666666667 0 -1.6 1e-06 
0.944444444444 0.666666666667 0 -1.6 1e-06 
1.0 0.666666666667 0 -1.6 1e-06 
0.5 0.707070707071 0 -1.6 1e-06 
0.555555555556 0.707070707071 0 -1.6 1e-06 
0.611111111111 0.707070707071 0 -1.6 1e-06 
0.666666666667 0.707070707071 0 -1.6 1e-06 
0.722222222222 0.707070707071 0 -1.6 1e-06 
0.777777777778 0.707070707071 0 -1.6 1e-06 
0.833333333333 0.707070707071 0 -1.6 1e-06 
0.888888888889 0.707070707071 0 -1.6 1e-06 
0.944444444444 0.707070707071 0 -1.6 1e-06 
1.0 0.707070707071 0 -1.6 1e-06 
0.5 0.747474747475 0 -1.6 1e-06 
0.555555555556 0.747474747475 0 -1.6 1e-06 
0.611111111111 0.747474747475 0 -1.6 1e-06 
0.666666666667 0.747474747475 0 -1.6 1e-06 
0.722222222222 0.747474747475 0 -1.6 1e-06 
0.777777777778 0.747474747475 0 -1.6 1e-06 
0.833333333333 0.747474747475 0 -1.6 1e-06 
0.888888888889 0.747474747475 0 -1.6 1e-06 
0.944444444444 0.747474747475 0 -1.6 1e-06 
1.0 0.747474747475 0 -1.6 1e-06 
0.5 0.787878787879 0 -1.6 1e-06 
0.555555555556 0.787878787879 0 -1.6 1e-06 
0.611111111111 0.787878787879 0 -1.6 1e-06 
0.666666666667 0.787878787879 0 -1.6 1e-06 
0.722222222222 0.787878787879 0 -1.6 1e-06 
0.777777777778 0.787878787879 0 -1.6 1e-06 
0.833333333333 0.787878787879 0 -1.6 1e-06 
0.888888888889 0.787878787879 0 -1.6 1e-06 
0.944444444444 0.787878787879 0 -1.6 1e-06 
1.0 0.787878787879 0 -1.6 1e-06 
0.5 0.828282828283 0 -1.6 1e-06 
0.555555555556 0.828282828283 0 -1.6 1e-06 
0.611111111111 0.828282828283 0 -1.6 1e-06 
0.666666666667 0.828282828283 0 -1.6 1e-06 
0.722222222222 0.828282828283 0 -1.6 1e-06 
0.777777777778 0.828282828283 0 -1.6 1e-06 
0.833333333333 0.828282828283 0 -1.6 1e-06 
0.888888888889 0.828282828283 0 -1.6 1e-06 
0.944444444444 0.828282828283 0 -1.6 1e-06 
1.0 0.828282828283 0 -1.6 1e-06 
0.5 0.868686868687 0 -1.6 1e-06 
0.555555555556 0.868686868687 0 -1.6 1e-06 
0.611111111111 0.868686868687 0 -1.6 1e-06 
0.666666666667 0.868686868687 0 -1.6 1e-06 
0.722222222222 0.868686868687 0 -1.6 1e-06 
0.777777777778 0.868686868687 0 -1.6 1e-06 
0.833333333333 0.868686868687 0 -1.6 1e-06 
0.888888888889 0.868686868687 0 -1.6 1e-06 
0.944444444444 0.868686868687 0 -1.6 1e-06 
1.0 0.868686868687 0 -1.6 1e-06 
0.5 0.909090909091 0 -1.6 1e-06 
0.555555555556 0.909090909091 0 -1.6 1e-06 
0.611111111111 0.909090909091 0 -1.6 1e-06 
0.666666666667 0.909090909091 0 -1.6 1e-06 
0.722222222222 0.909090909091 0 -1.6 1e-06 
0.777777777778 0.909090909091 0 -1.6 1e-06 
0.833333333333 0.909090909091 0 -1.6 1e-06 
0.888888888889 0.909090909091 0 -1.6 1e-06 
0.944444444444 0.909090909091 0 -1.6 1e-06 
1.0 0.909090909091 0 -1.6 1e-06 
0.5 0.949494949495 0 -1.6 1e-06 
0.555555555556 0.949494949495 0 -1.6 1e-06 
0.611111111111 0.949494949495 0 -1.6 1e-06 
0.666666666667 0.949494949495 0 -1.6 1e-06 
0.722222222222 0.949494949495 0 -1.6 1e-06 
0.777777777778 0.949494949495 0 -1.6 1e-06 
0.833333333333 0.949494949495 0 -1.6 1e-06 
0.888888888889 0.949494949495 0 -1.6 1e-06 
0.944444444444 0.949494949495 0 -1.6 1e-06 
1.0 0.949494949495 0 -1.6 1e-06 
0.5 0.989898989899 0 -1.6 1e-06 
0.555555555556 0.989898989899 0 -1.6 1e-06 
0.611111111111 0.989898989899 0 -1.6 1e-06 
0.666666666667 0.989898989899 0 -1.6 1e-06 
0.722222222222 0.989898989899 0 -1.6 1e-06 
0.777777777778 0.989898989899 0 -1.6 1e-06 
0.833333333333 0.989898989899 0 -1.6 1e-06 
0.888888888889 0.989898989899 0 -1.6 1e-06 
0.944444444444 0.989898989899 0 -1.6 1e-06 
1.0 0.989898989899 0 -1.6 1e-06 
0.5 1.0303030303 0 -1.6 1e-06 
0.555555555556 1.0303030303 0 -1.6 1e-06 
0.611111111111 1.0303030303 0 -1.6 1e-06 
0.666666666667 1.0303030303 0 -1.6 1e-06 
0.722222222222 1.0303030303 0 -1.6 1e-06 
0.777777777778 1.0303030303 0 -1.6 1e-06 
0.833333333333 1.0303030303 0 -1.6 1e-06 
0.888888888889 1.0303030303 0 -1.6 1e-06 
0.944444444444 1.0303030303 0 -1.6 1e-06 
1.0 1.0303030303 0 -1.6 1e-06 
0.5 1.07070707071 0 -1.6 1e-06 
0.555555555556 1.07070707071 0 -1.6 1e-06 
0.611111111111 1.07070707071 0 -1.6 1e-06 
0.666666666667 1.07070707071 0 -1.6 1e-06 
0.722222222222 1.07070707071 0 -1.6 1e-06 
0.777777777778 1.07070707071 0 -1.6 1e-06 
0.833333333333 1.07070707071 0 -1.6 1e-06 
0.888888888889 1.07070707071 0 -1.6 1e-06 
0.944444444444 1.07070707071 0 -1.6 1e-06 
1.0 1.07070707071 0 -1.6 1e-06 
0.5 1.11111111111 0 -1.6 1e-06 
0.555555555556 1.11111111111 0 -1.6 1e-06 
0.611111111111 1.11111111111 0 -1.6 1e-06 
0.666666666667 1.11111111111 0 -1.6 1e-06 
0.722222222222 1.11111111111 0 -1.6 1e-06 
0.777777777778 1.11111111111 0 -1.6 1e-06 
0.833333333333 1.11111111111 0 -1.6 1e-06 
0.888888888889 1.11111111111 0 -1.6 1e-06 
0.944444444444 1.11111111111 0 -1.6 1e-06 
1.0 1.11111111111 0 -1.6 1e-06 
0.5 1.15151515152 0 -1.6 1e-06 
0.555555555556 1.15151515152 0 -1.6 1e-06 
0.611111111111 1.15151515152 0 -1.6 1e-06 
0.666666666667 1.15151515152 0 -1.6 1e-06 
0.722222222222 1.15151515152 0 -1.6 1e-06 
0.777777777778 1.15151515152 0 -1.6 1e-06 
0.833333333333 1.15151515152 0 -1.6 1e-06 
0.888888888889 1.15151515152 0 -1.6 1e-06 
0.944444444444 1.15151515152 0 -1.6 1e-06 
1.0 1.15151515152 0 -1.6 1e-06 
0.5 1.19191919192 0 -1.6 1e-06 
0.555555555556 1.19191919192 0 -1.6 1e-06 
0.611111111111 1.19191919192 0 -1.6 1e-06 
0.666666666667 1.19191919192 0 -1.6 1e-06 
0.722222222222 1.19191919192 0 -1.6 1e-06 
0.777777777778 1.19191919192 0 -1.6 1e-06 
0.833333333333 1.19191919192 0 -1.6 1e-06 
0.888888888889 1.19191919192 0 -1.6 1e-06 
0.944444444444 1.19191919192 0 -1.6 1e-06 
1.0 1.19191919192 0 -1.6 1e-06 
0.5 1.23232323232 0 -1.6 1e-06 
0.555555555556 1.23232323232 0 -1.6 1e-06 
0.611111111111 1.23232323232 0 -1.6 1e-06 
0.666666666667 1.23232323232 0 -1.6 1e-06 
0.722222222222 1.23232323232 0 -1.6 1e-06 
0.777777777778 1.23232323232 0 -1.6 1e-06 
0.833333333333 1.23232323232 0 -1.6 1e-06 
0.888888888889 1.23232323232 0 -1.6 1e-06 
0.944444444444 1.23232323232 0 -1.6 1e-06 
1.0 1.23232323232 0 -1.6 1e-06 
0.5 1.27272727273 0 -1.6 1e-06 
0.555555555556 1.27272727273 0 -1.6 1e-06 
0.611111111111 1.27272727273 0 -1.6 1e-06 
0.666666666667 1.27272727273 0 -1.6 1e-06 
0.722222222222 1.27272727273 0 -1.6 1e-06 
0.777777777778 1.27272727273 0 -1.6 1e-06 
0.833333333333 1.27272727273 0 -1.6 1e-06 
0.888888888889 1.27272727273 0 -1.6 1e-06 
0.944444444444 1.27272727273 0 -1.6 1e-06 
1.0 1.27272727273 0 -1.6 1e-06 
0.5 1.31313131313 0 -1.6 1e-06 
0.555555555556 1.31313131313 0 -1.6 1e-06 
0.611111111111 1.31313131313 0 -1.6 1e-06 
0.666666666667 1.31313131313 0 -1.6 1e-06 
0.722222222222 1.31313131313 0 -1.6 1e-06 
0.777777777778 1.31313131313 0 -1.6 1e-06 
0.833333333333 1.31313131313 0 -1.6 1e-06 
0.888888888889 1.31313131313 0 -1.6 1e-06 
0.944444444444 1.31313131313 0 -1.6 1e-06 
1.0 1.31313131313 0 -1.6 1e-06 
0.5 1.35353535354 0 -1.6 1e-06 
0.555555555556 1.35353535354 0 -1.6 1e-06 
0.611111111111 1.35353535354 0 -1.6 1e-06 
0.666666666667 1.35353535354 0 -1.6 1e-06 
0.722222222222 1.35353535354 0 -1.6 1e-06 
0.777777777778 1.35353535354 0 -1.6 1e-06 
0.833333333333 1.35353535354 0 -1.6 1e-06 
0.888888888889 1.35353535354 0 -1.6 1e-06 
0.944444444444 1.35353535354 0 -1.6 1e-06 
1.0 1.35353535354 0 -1.6 1e-06 
0.5 1.39393939394 0 -1.6 1e-06 
0.555555555556 1.39393939394 0 -1.6 1e-06 
0.611111111111 1.39393939394 0 -1.6 1e-06 
0.666666666667 1.39393939394 0 -1.6 1e-06 
0.722222222222 1.39393939394 0 -1.6 1e-06 
0.777777777778 1.39393939394 0 -1.6 1e-06 
0.833333333333 1.39393939394 0 -1.6 1e-06 
0.888888888889 1.39393939394 0 -1.6 1e-06 
0.944444444444 1.39393939394 0 -1.6 1e-06 
1.0 1.39393939394 0 -1.6 1e-06 
0.5 1.43434343434 0 -1.6 1e-06 
0.555555555556 1.43434343434 0 -1.6 1e-06 
0.611111111111 1.43434343434 0 -1.6 1e-06 
0.666666666667 1.43434343434 0 -1.6 1e-06 
0.722222222222 1.43434343434 0 -1.6 1e-06 
0.777777777778 1.43434343434 0 -1.6 1e-06 
0.833333333333 1.43434343434 0 -1.6 1e-06 
0.888888888889 1.43434343434 0 -1.6 1e-06 
0.944444444444 1.43434343434 0 -1.6 1e-06 
1.0 1.43434343434 0 -1.6 1e-06 
0.5 1.47474747475 0 -1.6 1e-06 
0.555555555556 1.47474747475 0 -1.6 1e-06 
0.611111111111 1.47474747475 0 -1.6 1e-06 
0.666666666667 1.47474747475 0 -1.6 1e-06 
0.722222222222 1.47474747475 0 -1.6 1e-06 
0.777777777778 1.47474747475 0 -1.6 1e-06 
0.833333333333 1.47474747475 0 -1.6 1e-06 
0.888888888889 1.47474747475 0 -1.6 1e-06 
0.944444444444 1.47474747475 0 -1.6 1e-06 
1.0 1.47474747475 0 -1.6 1e-06 
0.5 1.51515151515 0 -1.6 1e-06 
0.555555555556 1.51515151515 0 -1.6 1e-06 
0.611111111111 1.51515151515 0 -1.6 1e-06 
0.666666666667 1.51515151515 0 -1.6 1e-06 
0.722222222222 1.51515151515 0 -1.6 1e-06 
0.777777777778 1.51515151515 0 -1.6 1e-06 
0.833333333333 1.51515151515 0 -1.6 1e-06 
0.888888888889 1.51515151515 0 -1.6 1e-06 
0.944444444444 1.51515151515 0 -1.6 1e-06 
1.0 1.51515151515 0 -1.6 1e-06 
0.5 1.55555555556 0 -1.6 1e-06 
0.555555555556 1.55555555556 0 -1.6 1e-06 
0.611111111111 1.55555555556 0 -1.6 1e-06 
0.666666666667 1.55555555556 0 -1.6 1e-06 
0.722222222222 1.55555555556 0 -1.6 1e-06 
0.777777777778 1.55555555556 0 -1.6 1e-06 
0.833333333333 1.55555555556 0 -1.6 1e-06 
0.888888888889 1.55555555556 0 -1.6 1e-06 
0.944444444444 1.55555555556 0 -1.6 1e-06 
1.0 1.55555555556 0 -1.6 1e-06 
0.5 1.59595959596 0 -1.6 1e-06 
0.555555555556 1.59595959596 0 -1.6 1e-06 
0.611111111111 1.59595959596 0 -1.6 1e-06 
0.666666666667 1.59595959596 0 -1.6 1e-06 
0.722222222222 1.59595959596 0 -1.6 1e-06 
0.777777777778 1.59595959596 0 -1.6 1e-06 
0.833333333333 1.59595959596 0 -1.6 1e-06 
0.888888888889 1.59595959596 0 -1.6 1e-06 
0.944444444444 1.59595959596 0 -1.6 1e-06 
1.0 1.59595959596 0 -1.6 1e-06 
0.5 1.63636363636 0 -1.6 1e-06 
0.555555555556 1.63636363636 0 -1.6 1e-06 
0.611111111111 1.63636363636 0 -1.6 1e-06 
0.666666666667 1.63636363636 0 -1.6 1e-06 
0.722222222222 1.63636363636 0 -1.6 1e-06 
0.777777777778 1.63636363636 0 -1.6 1e-06 
0.833333333333 1.63636363636 0 -1.6 1e-06 
0.888888888889 1.63636363636 0 -1.6 1e-06 
0.944444444444 1.63636363636 0 -1.6 1e-06 
1.0 1.63636363636 0 -1.6 1e-06 
0.5 1.67676767677 0 -1.6 1e-06 
0.555555555556 1.67676767677 0 -1.6 1e-06 
0.611111111111 1.67676767677 0 -1.6 1e-06 
0.666666666667 1.67676767677 0 -1.6 1e-06 
0.722222222222 1.67676767677 0 -1.6 1e-06 
0.777777777778 1.67676767677 0 -1.6 1e-06 
0.833333333333 1.67676767677 0 -1.6 1e-06 
0.888888888889 1.67676767677 0 -1.6 1e-06 
0.944444444444 1.67676767677 0 -1.6 1e-06 
1.0 1.67676767677 0 -1.6 1e-06 
0.5 1.71717171717 0 -1.6 1e-06 
0.555555555556 1.71717171717 0 -1.6 1e-06 
0.611111111111 1.71717171717 0 -1.6 1e-06 
0.666666666667 1.71717171717 0 -1.6 1e-06 
0.722222222222 1.71717171717 0 -1.6 1e-06 
0.777777777778 1.71717171717 0 -1.6 1e-06 
0.833333333333 1.71717171717 0 -1.6 1e-06 
0.888888888889 1.71717171717 0 -1.6 1e-06 
0.944444444444 1.71717171717 0 -1.6 1e-06 
1.0 1.71717171717 0 -1.6 1e-06 
0.5 1.75757575758 0 -1.6 1e-06 
0.555555555556 1.75757575758 0 -1.6 1e-06 
0.611111111111 1.75757575758 0 -1.6 1e-06 
0.666666666667 1.75757575758 0 -1.6 1e-06 
0.722222222222 1.75757575758 0 -1.6 1e-06 
0.777777777778 1.75757575758 0 -1.6 1e-06 
0.833333333333 1.75757575758 0 -1.6 1e-06 
0.888888888889 1.75757575758 0 -1.6 1e-06 
0.944444444444 1.75757575758 0 -1.6 1e-06 
1.0 1.75757575758 0 -1.6 1e-06 
0.5 1.79797979798 0 -1.6 1e-06 
0.555555555556 1.79797979798 0 -1.6 1e-06 
0.611111111111 1.79797979798 0 -1.6 1e-06 
0.666666666667 1.79797979798 0 -1.6 1e-06 
0.722222222222 1.79797979798 0 -1.6 1e-06 
0.777777777778 1.79797979798 0 -1.6 1e-06 
0.833333333333 1.79797979798 0 -1.6 1e-06 
0.888888888889 1.79797979798 0 -1.6 1e-06 
0.944444444444 1.79797979798 0 -1.6 1e-06 
1.0 1.79797979798 0 -1.6 1e-06 
0.5 1.83838383838 0 -1.6 1e-06 
0.555555555556 1.83838383838 0 -1.6 1e-06 
0.611111111111 1.83838383838 0 -1.6 1e-06 
0.666666666667 1.83838383838 0 -1.6 1e-06 
0.722222222222 1.83838383838 0 -1.6 1e-06 
0.777777777778 1.83838383838 0 -1.6 1e-06 
0.833333333333 1.83838383838 0 -1.6 1e-06 
0.888888888889 1.83838383838 0 -1.6 1e-06 
0.944444444444 1.83838383838 0 -1.6 1e-06 
1.0 1.83838383838 0 -1.6 1e-06 
0.5 1.87878787879 0 -1.6 1e-06 
0.555555555556 1.87878787879 0 -1.6 1e-06 
0.611111111111 1.87878787879 0 -1.6 1e-06 
0.666666666667 1.87878787879 0 -1.6 1e-06 
0.722222222222 1.87878787879 0 -1.6 1e-06 
0.777777777778 1.87878787879 0 -1.6 1e-06 
0.833333333333 1.87878787879 0 -1.6 1e-06 
0.888888888889 1.87878787879 0 -1.6 1e-06 
0.944444444444 1.87878787879 0 -1.6 1e-06 
1.0 1.87878787879 0 -1.6 1e-06 
0.5 1.91919191919 0 -1.6 1e-06 
0.555555555556 1.91919191919 0 -1.6 1e-06 
0.611111111111 1.91919191919 0 -1.6 1e-06 
0.666666666667 1.91919191919 0 -1.6 1e-06 
0.722222222222 1.91919191919 0 -1.6 1e-06 
0.777777777778 1.91919191919 0 -1.6 1e-06 
0.833333333333 1.91919191919 0 -1.6 1e-06 
0.888888888889 1.91919191919 0 -1.6 1e-06 
0.944444444444 1.91919191919 0 -1.6 1e-06 
1.0 1.91919191919 0 -1.6 1e-06 
0.5 1.9595959596 0 -1.6 1e-06 
0.555555555556 1.9595959596 0 -1.6 1e-06 
0.611111111111 1.9595959596 0 -1.6 1e-06 
0.666666666667 1.9595959596 0 -1.6 1e-06 
0.722222222222 1.9595959596 0 -1.6 1e-06 
0.777777777778 1.9595959596 0 -1.6 1e-06 
0.833333333333 1.9595959596 0 -1.6 1e-06 
0.888888888889 1.9595959596 0 -1.6 1e-06 
0.944444444444 1.9595959596 0 -1.6 1e-06 
1.0 1.9595959596 0 -1.6 1e-06 
0.5 2.0 0 -1.6 1e-06 
0.555555555556 2.0 0 -1.6 1e-06 
0.611111111111 2.0 0 -1.6 1e-06 
0.666666666667 2.0 0 -1.6 1e-06 
0.722222222222 2.0 0 -1.6 1e-06 
0.777777777778 2.0 0 -1.6 1e-06 
0.833333333333 2.0 0 -1.6 1e-06 
0.888888888889 2.0 0 -1.6 1e-06 
0.944444444444 2.0 0 -1.6 1e-06 
1.0 2.0 0 -1.6 1e-06 
0.5 -2.0 0 -1.2 1e-06 
0.555555555556 -2.0 0 -1.2 1e-06 
0.611111111111 -2.0 0 -1.2 1e-06 
0.666666666667 -2.0 0 -1.2 1e-06 
0.722222222222 -2.0 0 -1.2 1e-06 
0.777777777778 -2.0 0 -1.2 1e-06 
0.833333333333 -2.0 0 -1.2 1e-06 
0.888888888889 -2.0 0 -1.2 1e-06 
0.944444444444 -2.0 0 -1.2 1e-06 
1.0 -2.0 0 -1.2 1e-06 
0.5 -1.9595959596 0 -1.2 1e-06 
0.555555555556 -1.9595959596 0 -1.2 1e-06 
0.611111111111 -1.9595959596 0 -1.2 1e-06 
0.666666666667 -1.9595959596 0 -1.2 1e-06 
0.722222222222 -1.9595959596 0 -1.2 1e-06 
0.777777777778 -1.9595959596 0 -1.2 1e-06 
0.833333333333 -1.9595959596 0 -1.2 1e-06 
0.888888888889 -1.9595959596 0 -1.2 1e-06 
0.944444444444 -1.9595959596 0 -1.2 1e-06 
1.0 -1.9595959596 0 -1.2 1e-06 
0.5 -1.91919191919 0 -1.2 1e-06 
0.555555555556 -1.91919191919 0 -1.2 1e-06 
0.611111111111 -1.91919191919 0 -1.2 1e-06 
0.666666666667 -1.91919191919 0 -1.2 1e-06 
0.722222222222 -1.91919191919 0 -1.2 1e-06 
0.777777777778 -1.91919191919 0 -1.2 1e-06 
0.833333333333 -1.91919191919 0 -1.2 1e-06 
0.888888888889 -1.91919191919 0 -1.2 1e-06 
0.944444444444 -1.91919191919 0 -1.2 1e-06 
1.0 -1.91919191919 0 -1.2 1e-06 
0.5 -1.87878787879 0 -1.2 1e-06 
0.555555555556 -1.87878787879 0 -1.2 1e-06 
0.611111111111 -1.87878787879 0 -1.2 1e-06 
0.666666666667 -1.87878787879 0 -1.2 1e-06 
0.722222222222 -1.87878787879 0 -1.2 1e-06 
0.777777777778 -1.87878787879 0 -1.2 1e-06 
0.833333333333 -1.87878787879 0 -1.2 1e-06 
0.888888888889 -1.87878787879 0 -1.2 1e-06 
0.944444444444 -1.87878787879 0 -1.2 1e-06 
1.0 -1.87878787879 0 -1.2 1e-06 
0.5 -1.83838383838 0 -1.2 1e-06 
0.555555555556 -1.83838383838 0 -1.2 1e-06 
0.611111111111 -1.83838383838 0 -1.2 1e-06 
0.666666666667 -1.83838383838 0 -1.2 1e-06 
0.722222222222 -1.83838383838 0 -1.2 1e-06 
0.777777777778 -1.83838383838 0 -1.2 1e-06 
0.833333333333 -1.83838383838 0 -1.2 1e-06 
0.888888888889 -1.83838383838 0 -1.2 1e-06 
0.944444444444 -1.83838383838 0 -1.2 1e-06 
1.0 -1.83838383838 0 -1.2 1e-06 
0.5 -1.79797979798 0 -1.2 1e-06 
0.555555555556 -1.79797979798 0 -1.2 1e-06 
0.611111111111 -1.79797979798 0 -1.2 1e-06 
0.666666666667 -1.79797979798 0 -1.2 1e-06 
0.722222222222 -1.79797979798 0 -1.2 1e-06 
0.777777777778 -1.79797979798 0 -1.2 1e-06 
0.833333333333 -1.79797979798 0 -1.2 1e-06 
0.888888888889 -1.79797979798 0 -1.2 1e-06 
0.944444444444 -1.79797979798 0 -1.2 1e-06 
1.0 -1.79797979798 0 -1.2 1e-06 
0.5 -1.75757575758 0 -1.2 1e-06 
0.555555555556 -1.75757575758 0 -1.2 1e-06 
0.611111111111 -1.75757575758 0 -1.2 1e-06 
0.666666666667 -1.75757575758 0 -1.2 1e-06 
0.722222222222 -1.75757575758 0 -1.2 1e-06 
0.777777777778 -1.75757575758 0 -1.2 1e-06 
0.833333333333 -1.75757575758 0 -1.2 1e-06 
0.888888888889 -1.75757575758 0 -1.2 1e-06 
0.944444444444 -1.75757575758 0 -1.2 1e-06 
1.0 -1.75757575758 0 -1.2 1e-06 
0.5 -1.71717171717 0 -1.2 1e-06 
0.555555555556 -1.71717171717 0 -1.2 1e-06 
0.611111111111 -1.71717171717 0 -1.2 1e-06 
0.666666666667 -1.71717171717 0 -1.2 1e-06 
0.722222222222 -1.71717171717 0 -1.2 1e-06 
0.777777777778 -1.71717171717 0 -1.2 1e-06 
0.833333333333 -1.71717171717 0 -1.2 1e-06 
0.888888888889 -1.71717171717 0 -1.2 1e-06 
0.944444444444 -1.71717171717 0 -1.2 1e-06 
1.0 -1.71717171717 0 -1.2 1e-06 
0.5 -1.67676767677 0 -1.2 1e-06 
0.555555555556 -1.67676767677 0 -1.2 1e-06 
0.611111111111 -1.67676767677 0 -1.2 1e-06 
0.666666666667 -1.67676767677 0 -1.2 1e-06 
0.722222222222 -1.67676767677 0 -1.2 1e-06 
0.777777777778 -1.67676767677 0 -1.2 1e-06 
0.833333333333 -1.67676767677 0 -1.2 1e-06 
0.888888888889 -1.67676767677 0 -1.2 1e-06 
0.944444444444 -1.67676767677 0 -1.2 1e-06 
1.0 -1.67676767677 0 -1.2 1e-06 
0.5 -1.63636363636 0 -1.2 1e-06 
0.555555555556 -1.63636363636 0 -1.2 1e-06 
0.611111111111 -1.63636363636 0 -1.2 1e-06 
0.666666666667 -1.63636363636 0 -1.2 1e-06 
0.722222222222 -1.63636363636 0 -1.2 1e-06 
0.777777777778 -1.63636363636 0 -1.2 1e-06 
0.833333333333 -1.63636363636 0 -1.2 1e-06 
0.888888888889 -1.63636363636 0 -1.2 1e-06 
0.944444444444 -1.63636363636 0 -1.2 1e-06 
1.0 -1.63636363636 0 -1.2 1e-06 
0.5 -1.59595959596 0 -1.2 1e-06 
0.555555555556 -1.59595959596 0 -1.2 1e-06 
0.611111111111 -1.59595959596 0 -1.2 1e-06 
0.666666666667 -1.59595959596 0 -1.2 1e-06 
0.722222222222 -1.59595959596 0 -1.2 1e-06 
0.777777777778 -1.59595959596 0 -1.2 1e-06 
0.833333333333 -1.59595959596 0 -1.2 1e-06 
0.888888888889 -1.59595959596 0 -1.2 1e-06 
0.944444444444 -1.59595959596 0 -1.2 1e-06 
1.0 -1.59595959596 0 -1.2 1e-06 
0.5 -1.55555555556 0 -1.2 1e-06 
0.555555555556 -1.55555555556 0 -1.2 1e-06 
0.611111111111 -1.55555555556 0 -1.2 1e-06 
0.666666666667 -1.55555555556 0 -1.2 1e-06 
0.722222222222 -1.55555555556 0 -1.2 1e-06 
0.777777777778 -1.55555555556 0 -1.2 1e-06 
0.833333333333 -1.55555555556 0 -1.2 1e-06 
0.888888888889 -1.55555555556 0 -1.2 1e-06 
0.944444444444 -1.55555555556 0 -1.2 1e-06 
1.0 -1.55555555556 0 -1.2 1e-06 
0.5 -1.51515151515 0 -1.2 1e-06 
0.555555555556 -1.51515151515 0 -1.2 1e-06 
0.611111111111 -1.51515151515 0 -1.2 1e-06 
0.666666666667 -1.51515151515 0 -1.2 1e-06 
0.722222222222 -1.51515151515 0 -1.2 1e-06 
0.777777777778 -1.51515151515 0 -1.2 1e-06 
0.833333333333 -1.51515151515 0 -1.2 1e-06 
0.888888888889 -1.51515151515 0 -1.2 1e-06 
0.944444444444 -1.51515151515 0 -1.2 1e-06 
1.0 -1.51515151515 0 -1.2 1e-06 
0.5 -1.47474747475 0 -1.2 1e-06 
0.555555555556 -1.47474747475 0 -1.2 1e-06 
0.611111111111 -1.47474747475 0 -1.2 1e-06 
0.666666666667 -1.47474747475 0 -1.2 1e-06 
0.722222222222 -1.47474747475 0 -1.2 1e-06 
0.777777777778 -1.47474747475 0 -1.2 1e-06 
0.833333333333 -1.47474747475 0 -1.2 1e-06 
0.888888888889 -1.47474747475 0 -1.2 1e-06 
0.944444444444 -1.47474747475 0 -1.2 1e-06 
1.0 -1.47474747475 0 -1.2 1e-06 
0.5 -1.43434343434 0 -1.2 1e-06 
0.555555555556 -1.43434343434 0 -1.2 1e-06 
0.611111111111 -1.43434343434 0 -1.2 1e-06 
0.666666666667 -1.43434343434 0 -1.2 1e-06 
0.722222222222 -1.43434343434 0 -1.2 1e-06 
0.777777777778 -1.43434343434 0 -1.2 1e-06 
0.833333333333 -1.43434343434 0 -1.2 1e-06 
0.888888888889 -1.43434343434 0 -1.2 1e-06 
0.944444444444 -1.43434343434 0 -1.2 1e-06 
1.0 -1.43434343434 0 -1.2 1e-06 
0.5 -1.39393939394 0 -1.2 1e-06 
0.555555555556 -1.39393939394 0 -1.2 1e-06 
0.611111111111 -1.39393939394 0 -1.2 1e-06 
0.666666666667 -1.39393939394 0 -1.2 1e-06 
0.722222222222 -1.39393939394 0 -1.2 1e-06 
0.777777777778 -1.39393939394 0 -1.2 1e-06 
0.833333333333 -1.39393939394 0 -1.2 1e-06 
0.888888888889 -1.39393939394 0 -1.2 1e-06 
0.944444444444 -1.39393939394 0 -1.2 1e-06 
1.0 -1.39393939394 0 -1.2 1e-06 
0.5 -1.35353535354 0 -1.2 1e-06 
0.555555555556 -1.35353535354 0 -1.2 1e-06 
0.611111111111 -1.35353535354 0 -1.2 1e-06 
0.666666666667 -1.35353535354 0 -1.2 1e-06 
0.722222222222 -1.35353535354 0 -1.2 1e-06 
0.777777777778 -1.35353535354 0 -1.2 1e-06 
0.833333333333 -1.35353535354 0 -1.2 1e-06 
0.888888888889 -1.35353535354 0 -1.2 1e-06 
0.944444444444 -1.35353535354 0 -1.2 1e-06 
1.0 -1.35353535354 0 -1.2 1e-06 
0.5 -1.31313131313 0 -1.2 1e-06 
0.555555555556 -1.31313131313 0 -1.2 1e-06 
0.611111111111 -1.31313131313 0 -1.2 1e-06 
0.666666666667 -1.31313131313 0 -1.2 1e-06 
0.722222222222 -1.31313131313 0 -1.2 1e-06 
0.777777777778 -1.31313131313 0 -1.2 1e-06 
0.833333333333 -1.31313131313 0 -1.2 1e-06 
0.888888888889 -1.31313131313 0 -1.2 1e-06 
0.944444444444 -1.31313131313 0 -1.2 1e-06 
1.0 -1.31313131313 0 -1.2 1e-06 
0.5 -1.27272727273 0 -1.2 1e-06 
0.555555555556 -1.27272727273 0 -1.2 1e-06 
0.611111111111 -1.27272727273 0 -1.2 1e-06 
0.666666666667 -1.27272727273 0 -1.2 1e-06 
0.722222222222 -1.27272727273 0 -1.2 1e-06 
0.777777777778 -1.27272727273 0 -1.2 1e-06 
0.833333333333 -1.27272727273 0 -1.2 1e-06 
0.888888888889 -1.27272727273 0 -1.2 1e-06 
0.944444444444 -1.27272727273 0 -1.2 1e-06 
1.0 -1.27272727273 0 -1.2 1e-06 
0.5 -1.23232323232 0 -1.2 1e-06 
0.555555555556 -1.23232323232 0 -1.2 1e-06 
0.611111111111 -1.23232323232 0 -1.2 1e-06 
0.666666666667 -1.23232323232 0 -1.2 1e-06 
0.722222222222 -1.23232323232 0 -1.2 1e-06 
0.777777777778 -1.23232323232 0 -1.2 1e-06 
0.833333333333 -1.23232323232 0 -1.2 1e-06 
0.888888888889 -1.23232323232 0 -1.2 1e-06 
0.944444444444 -1.23232323232 0 -1.2 1e-06 
1.0 -1.23232323232 0 -1.2 1e-06 
0.5 -1.19191919192 0 -1.2 1e-06 
0.555555555556 -1.19191919192 0 -1.2 1e-06 
0.611111111111 -1.19191919192 0 -1.2 1e-06 
0.666666666667 -1.19191919192 0 -1.2 1e-06 
0.722222222222 -1.19191919192 0 -1.2 1e-06 
0.777777777778 -1.19191919192 0 -1.2 1e-06 
0.833333333333 -1.19191919192 0 -1.2 1e-06 
0.888888888889 -1.19191919192 0 -1.2 1e-06 
0.944444444444 -1.19191919192 0 -1.2 1e-06 
1.0 -1.19191919192 0 -1.2 1e-06 
0.5 -1.15151515152 0 -1.2 1e-06 
0.555555555556 -1.15151515152 0 -1.2 1e-06 
0.611111111111 -1.15151515152 0 -1.2 1e-06 
0.666666666667 -1.15151515152 0 -1.2 1e-06 
0.722222222222 -1.15151515152 0 -1.2 1e-06 
0.777777777778 -1.15151515152 0 -1.2 1e-06 
0.833333333333 -1.15151515152 0 -1.2 1e-06 
0.888888888889 -1.15151515152 0 -1.2 1e-06 
0.944444444444 -1.15151515152 0 -1.2 1e-06 
1.0 -1.15151515152 0 -1.2 1e-06 
0.5 -1.11111111111 0 -1.2 1e-06 
0.555555555556 -1.11111111111 0 -1.2 1e-06 
0.611111111111 -1.11111111111 0 -1.2 1e-06 
0.666666666667 -1.11111111111 0 -1.2 1e-06 
0.722222222222 -1.11111111111 0 -1.2 1e-06 
0.777777777778 -1.11111111111 0 -1.2 1e-06 
0.833333333333 -1.11111111111 0 -1.2 1e-06 
0.888888888889 -1.11111111111 0 -1.2 1e-06 
0.944444444444 -1.11111111111 0 -1.2 1e-06 
1.0 -1.11111111111 0 -1.2 1e-06 
0.5 -1.07070707071 0 -1.2 1e-06 
0.555555555556 -1.07070707071 0 -1.2 1e-06 
0.611111111111 -1.07070707071 0 -1.2 1e-06 
0.666666666667 -1.07070707071 0 -1.2 1e-06 
0.722222222222 -1.07070707071 0 -1.2 1e-06 
0.777777777778 -1.07070707071 0 -1.2 1e-06 
0.833333333333 -1.07070707071 0 -1.2 1e-06 
0.888888888889 -1.07070707071 0 -1.2 1e-06 
0.944444444444 -1.07070707071 0 -1.2 1e-06 
1.0 -1.07070707071 0 -1.2 1e-06 
0.5 -1.0303030303 0 -1.2 1e-06 
0.555555555556 -1.0303030303 0 -1.2 1e-06 
0.611111111111 -1.0303030303 0 -1.2 1e-06 
0.666666666667 -1.0303030303 0 -1.2 1e-06 
0.722222222222 -1.0303030303 0 -1.2 1e-06 
0.777777777778 -1.0303030303 0 -1.2 1e-06 
0.833333333333 -1.0303030303 0 -1.2 1e-06 
0.888888888889 -1.0303030303 0 -1.2 1e-06 
0.944444444444 -1.0303030303 0 -1.2 1e-06 
1.0 -1.0303030303 0 -1.2 1e-06 
0.5 -0.989898989899 0 -1.2 1e-06 
0.555555555556 -0.989898989899 0 -1.2 1e-06 
0.611111111111 -0.989898989899 0 -1.2 1e-06 
0.666666666667 -0.989898989899 0 -1.2 1e-06 
0.722222222222 -0.989898989899 0 -1.2 1e-06 
0.777777777778 -0.989898989899 0 -1.2 1e-06 
0.833333333333 -0.989898989899 0 -1.2 1e-06 
0.888888888889 -0.989898989899 0 -1.2 1e-06 
0.944444444444 -0.989898989899 0 -1.2 1e-06 
1.0 -0.989898989899 0 -1.2 1e-06 
0.5 -0.949494949495 0 -1.2 1e-06 
0.555555555556 -0.949494949495 0 -1.2 1e-06 
0.611111111111 -0.949494949495 0 -1.2 1e-06 
0.666666666667 -0.949494949495 0 -1.2 1e-06 
0.722222222222 -0.949494949495 0 -1.2 1e-06 
0.777777777778 -0.949494949495 0 -1.2 1e-06 
0.833333333333 -0.949494949495 0 -1.2 1e-06 
0.888888888889 -0.949494949495 0 -1.2 1e-06 
0.944444444444 -0.949494949495 0 -1.2 1e-06 
1.0 -0.949494949495 0 -1.2 1e-06 
0.5 -0.909090909091 0 -1.2 1e-06 
0.555555555556 -0.909090909091 0 -1.2 1e-06 
0.611111111111 -0.909090909091 0 -1.2 1e-06 
0.666666666667 -0.909090909091 0 -1.2 1e-06 
0.722222222222 -0.909090909091 0 -1.2 1e-06 
0.777777777778 -0.909090909091 0 -1.2 1e-06 
0.833333333333 -0.909090909091 0 -1.2 1e-06 
0.888888888889 -0.909090909091 0 -1.2 1e-06 
0.944444444444 -0.909090909091 0 -1.2 1e-06 
1.0 -0.909090909091 0 -1.2 1e-06 
0.5 -0.868686868687 0 -1.2 1e-06 
0.555555555556 -0.868686868687 0 -1.2 1e-06 
0.611111111111 -0.868686868687 0 -1.2 1e-06 
0.666666666667 -0.868686868687 0 -1.2 1e-06 
0.722222222222 -0.868686868687 0 -1.2 1e-06 
0.777777777778 -0.868686868687 0 -1.2 1e-06 
0.833333333333 -0.868686868687 0 -1.2 1e-06 
0.888888888889 -0.868686868687 0 -1.2 1e-06 
0.944444444444 -0.868686868687 0 -1.2 1e-06 
1.0 -0.868686868687 0 -1.2 1e-06 
0.5 -0.828282828283 0 -1.2 1e-06 
0.555555555556 -0.828282828283 0 -1.2 1e-06 
0.611111111111 -0.828282828283 0 -1.2 1e-06 
0.666666666667 -0.828282828283 0 -1.2 1e-06 
0.722222222222 -0.828282828283 0 -1.2 1e-06 
0.777777777778 -0.828282828283 0 -1.2 1e-06 
0.833333333333 -0.828282828283 0 -1.2 1e-06 
0.888888888889 -0.828282828283 0 -1.2 1e-06 
0.944444444444 -0.828282828283 0 -1.2 1e-06 
1.0 -0.828282828283 0 -1.2 1e-06 
0.5 -0.787878787879 0 -1.2 1e-06 
0.555555555556 -0.787878787879 0 -1.2 1e-06 
0.611111111111 -0.787878787879 0 -1.2 1e-06 
0.666666666667 -0.787878787879 0 -1.2 1e-06 
0.722222222222 -0.787878787879 0 -1.2 1e-06 
0.777777777778 -0.787878787879 0 -1.2 1e-06 
0.833333333333 -0.787878787879 0 -1.2 1e-06 
0.888888888889 -0.787878787879 0 -1.2 1e-06 
0.944444444444 -0.787878787879 0 -1.2 1e-06 
1.0 -0.787878787879 0 -1.2 1e-06 
0.5 -0.747474747475 0 -1.2 1e-06 
0.555555555556 -0.747474747475 0 -1.2 1e-06 
0.611111111111 -0.747474747475 0 -1.2 1e-06 
0.666666666667 -0.747474747475 0 -1.2 1e-06 
0.722222222222 -0.747474747475 0 -1.2 1e-06 
0.777777777778 -0.747474747475 0 -1.2 1e-06 
0.833333333333 -0.747474747475 0 -1.2 1e-06 
0.888888888889 -0.747474747475 0 -1.2 1e-06 
0.944444444444 -0.747474747475 0 -1.2 1e-06 
1.0 -0.747474747475 0 -1.2 1e-06 
0.5 -0.707070707071 0 -1.2 1e-06 
0.555555555556 -0.707070707071 0 -1.2 1e-06 
0.611111111111 -0.707070707071 0 -1.2 1e-06 
0.666666666667 -0.707070707071 0 -1.2 1e-06 
0.722222222222 -0.707070707071 0 -1.2 1e-06 
0.777777777778 -0.707070707071 0 -1.2 1e-06 
0.833333333333 -0.707070707071 0 -1.2 1e-06 
0.888888888889 -0.707070707071 0 -1.2 1e-06 
0.944444444444 -0.707070707071 0 -1.2 1e-06 
1.0 -0.707070707071 0 -1.2 1e-06 
0.5 -0.666666666667 0 -1.2 1e-06 
0.555555555556 -0.666666666667 0 -1.2 1e-06 
0.611111111111 -0.666666666667 0 -1.2 1e-06 
0.666666666667 -0.666666666667 0 -1.2 1e-06 
0.722222222222 -0.666666666667 0 -1.2 1e-06 
0.777777777778 -0.666666666667 0 -1.2 1e-06 
0.833333333333 -0.666666666667 0 -1.2 1e-06 
0.888888888889 -0.666666666667 0 -1.2 1e-06 
0.944444444444 -0.666666666667 0 -1.2 1e-06 
1.0 -0.666666666667 0 -1.2 1e-06 
0.5 -0.626262626263 0 -1.2 1e-06 
0.555555555556 -0.626262626263 0 -1.2 1e-06 
0.611111111111 -0.626262626263 0 -1.2 1e-06 
0.666666666667 -0.626262626263 0 -1.2 1e-06 
0.722222222222 -0.626262626263 0 -1.2 1e-06 
0.777777777778 -0.626262626263 0 -1.2 1e-06 
0.833333333333 -0.626262626263 0 -1.2 1e-06 
0.888888888889 -0.626262626263 0 -1.2 1e-06 
0.944444444444 -0.626262626263 0 -1.2 1e-06 
1.0 -0.626262626263 0 -1.2 1e-06 
0.5 -0.585858585859 0 -1.2 1e-06 
0.555555555556 -0.585858585859 0 -1.2 1e-06 
0.611111111111 -0.585858585859 0 -1.2 1e-06 
0.666666666667 -0.585858585859 0 -1.2 1e-06 
0.722222222222 -0.585858585859 0 -1.2 1e-06 
0.777777777778 -0.585858585859 0 -1.2 1e-06 
0.833333333333 -0.585858585859 0 -1.2 1e-06 
0.888888888889 -0.585858585859 0 -1.2 1e-06 
0.944444444444 -0.585858585859 0 -1.2 1e-06 
1.0 -0.585858585859 0 -1.2 1e-06 
0.5 -0.545454545455 0 -1.2 1e-06 
0.555555555556 -0.545454545455 0 -1.2 1e-06 
0.611111111111 -0.545454545455 0 -1.2 1e-06 
0.666666666667 -0.545454545455 0 -1.2 1e-06 
0.722222222222 -0.545454545455 0 -1.2 1e-06 
0.777777777778 -0.545454545455 0 -1.2 1e-06 
0.833333333333 -0.545454545455 0 -1.2 1e-06 
0.888888888889 -0.545454545455 0 -1.2 1e-06 
0.944444444444 -0.545454545455 0 -1.2 1e-06 
1.0 -0.545454545455 0 -1.2 1e-06 
0.5 -0.505050505051 0 -1.2 1e-06 
0.555555555556 -0.505050505051 0 -1.2 1e-06 
0.611111111111 -0.505050505051 0 -1.2 1e-06 
0.666666666667 -0.505050505051 0 -1.2 1e-06 
0.722222222222 -0.505050505051 0 -1.2 1e-06 
0.777777777778 -0.505050505051 0 -1.2 1e-06 
0.833333333333 -0.505050505051 0 -1.2 1e-06 
0.888888888889 -0.505050505051 0 -1.2 1e-06 
0.944444444444 -0.505050505051 0 -1.2 1e-06 
1.0 -0.505050505051 0 -1.2 1e-06 
0.5 -0.464646464646 0 -1.2 1e-06 
0.555555555556 -0.464646464646 0 -1.2 1e-06 
0.611111111111 -0.464646464646 0 -1.2 1e-06 
0.666666666667 -0.464646464646 0 -1.2 1e-06 
0.722222222222 -0.464646464646 0 -1.2 1e-06 
0.777777777778 -0.464646464646 0 -1.2 1e-06 
0.833333333333 -0.464646464646 0 -1.2 1e-06 
0.888888888889 -0.464646464646 0 -1.2 1e-06 
0.944444444444 -0.464646464646 0 -1.2 1e-06 
1.0 -0.464646464646 0 -1.2 1e-06 
0.5 -0.424242424242 0 -1.2 1e-06 
0.555555555556 -0.424242424242 0 -1.2 1e-06 
0.611111111111 -0.424242424242 0 -1.2 1e-06 
0.666666666667 -0.424242424242 0 -1.2 1e-06 
0.722222222222 -0.424242424242 0 -1.2 1e-06 
0.777777777778 -0.424242424242 0 -1.2 1e-06 
0.833333333333 -0.424242424242 0 -1.2 1e-06 
0.888888888889 -0.424242424242 0 -1.2 1e-06 
0.944444444444 -0.424242424242 0 -1.2 1e-06 
1.0 -0.424242424242 0 -1.2 1e-06 
0.5 -0.383838383838 0 -1.2 1e-06 
0.555555555556 -0.383838383838 0 -1.2 1e-06 
0.611111111111 -0.383838383838 0 -1.2 1e-06 
0.666666666667 -0.383838383838 0 -1.2 1e-06 
0.722222222222 -0.383838383838 0 -1.2 1e-06 
0.777777777778 -0.383838383838 0 -1.2 1e-06 
0.833333333333 -0.383838383838 0 -1.2 1e-06 
0.888888888889 -0.383838383838 0 -1.2 1e-06 
0.944444444444 -0.383838383838 0 -1.2 1e-06 
1.0 -0.383838383838 0 -1.2 1e-06 
0.5 -0.343434343434 0 -1.2 1e-06 
0.555555555556 -0.343434343434 0 -1.2 1e-06 
0.611111111111 -0.343434343434 0 -1.2 1e-06 
0.666666666667 -0.343434343434 0 -1.2 1e-06 
0.722222222222 -0.343434343434 0 -1.2 1e-06 
0.777777777778 -0.343434343434 0 -1.2 1e-06 
0.833333333333 -0.343434343434 0 -1.2 1e-06 
0.888888888889 -0.343434343434 0 -1.2 1e-06 
0.944444444444 -0.343434343434 0 -1.2 1e-06 
1.0 -0.343434343434 0 -1.2 1e-06 
0.5 -0.30303030303 0 -1.2 1e-06 
0.555555555556 -0.30303030303 0 -1.2 1e-06 
0.611111111111 -0.30303030303 0 -1.2 1e-06 
0.666666666667 -0.30303030303 0 -1.2 1e-06 
0.722222222222 -0.30303030303 0 -1.2 1e-06 
0.777777777778 -0.30303030303 0 -1.2 1e-06 
0.833333333333 -0.30303030303 0 -1.2 1e-06 
0.888888888889 -0.30303030303 0 -1.2 1e-06 
0.944444444444 -0.30303030303 0 -1.2 1e-06 
1.0 -0.30303030303 0 -1.2 1e-06 
0.5 -0.262626262626 0 -1.2 1e-06 
0.555555555556 -0.262626262626 0 -1.2 1e-06 
0.611111111111 -0.262626262626 0 -1.2 1e-06 
0.666666666667 -0.262626262626 0 -1.2 1e-06 
0.722222222222 -0.262626262626 0 -1.2 1e-06 
0.777777777778 -0.262626262626 0 -1.2 1e-06 
0.833333333333 -0.262626262626 0 -1.2 1e-06 
0.888888888889 -0.262626262626 0 -1.2 1e-06 
0.944444444444 -0.262626262626 0 -1.2 1e-06 
1.0 -0.262626262626 0 -1.2 1e-06 
0.5 -0.222222222222 0 -1.2 1e-06 
0.555555555556 -0.222222222222 0 -1.2 1e-06 
0.611111111111 -0.222222222222 0 -1.2 1e-06 
0.666666666667 -0.222222222222 0 -1.2 1e-06 
0.722222222222 -0.222222222222 0 -1.2 1e-06 
0.777777777778 -0.222222222222 0 -1.2 1e-06 
0.833333333333 -0.222222222222 0 -1.2 1e-06 
0.888888888889 -0.222222222222 0 -1.2 1e-06 
0.944444444444 -0.222222222222 0 -1.2 1e-06 
1.0 -0.222222222222 0 -1.2 1e-06 
0.5 -0.181818181818 0 -1.2 1e-06 
0.555555555556 -0.181818181818 0 -1.2 1e-06 
0.611111111111 -0.181818181818 0 -1.2 1e-06 
0.666666666667 -0.181818181818 0 -1.2 1e-06 
0.722222222222 -0.181818181818 0 -1.2 1e-06 
0.777777777778 -0.181818181818 0 -1.2 1e-06 
0.833333333333 -0.181818181818 0 -1.2 1e-06 
0.888888888889 -0.181818181818 0 -1.2 1e-06 
0.944444444444 -0.181818181818 0 -1.2 1e-06 
1.0 -0.181818181818 0 -1.2 1e-06 
0.5 -0.141414141414 0 -1.2 1e-06 
0.555555555556 -0.141414141414 0 -1.2 1e-06 
0.611111111111 -0.141414141414 0 -1.2 1e-06 
0.666666666667 -0.141414141414 0 -1.2 1e-06 
0.722222222222 -0.141414141414 0 -1.2 1e-06 
0.777777777778 -0.141414141414 0 -1.2 1e-06 
0.833333333333 -0.141414141414 0 -1.2 1e-06 
0.888888888889 -0.141414141414 0 -1.2 1e-06 
0.944444444444 -0.141414141414 0 -1.2 1e-06 
1.0 -0.141414141414 0 -1.2 1e-06 
0.5 -0.10101010101 0 -1.2 1e-06 
0.555555555556 -0.10101010101 0 -1.2 1e-06 
0.611111111111 -0.10101010101 0 -1.2 1e-06 
0.666666666667 -0.10101010101 0 -1.2 1e-06 
0.722222222222 -0.10101010101 0 -1.2 1e-06 
0.777777777778 -0.10101010101 0 -1.2 1e-06 
0.833333333333 -0.10101010101 0 -1.2 1e-06 
0.888888888889 -0.10101010101 0 -1.2 1e-06 
0.944444444444 -0.10101010101 0 -1.2 1e-06 
1.0 -0.10101010101 0 -1.2 1e-06 
0.5 -0.0606060606061 0 -1.2 1e-06 
0.555555555556 -0.0606060606061 0 -1.2 1e-06 
0.611111111111 -0.0606060606061 0 -1.2 1e-06 
0.666666666667 -0.0606060606061 0 -1.2 1e-06 
0.722222222222 -0.0606060606061 0 -1.2 1e-06 
0.777777777778 -0.0606060606061 0 -1.2 1e-06 
0.833333333333 -0.0606060606061 0 -1.2 1e-06 
0.888888888889 -0.0606060606061 0 -1.2 1e-06 
0.944444444444 -0.0606060606061 0 -1.2 1e-06 
1.0 -0.0606060606061 0 -1.2 1e-06 
0.5 -0.020202020202 0 -1.2 1e-06 
0.555555555556 -0.020202020202 0 -1.2 1e-06 
0.611111111111 -0.020202020202 0 -1.2 1e-06 
0.666666666667 -0.020202020202 0 -1.2 1e-06 
0.722222222222 -0.020202020202 0 -1.2 1e-06 
0.777777777778 -0.020202020202 0 -1.2 1e-06 
0.833333333333 -0.020202020202 0 -1.2 1e-06 
0.888888888889 -0.020202020202 0 -1.2 1e-06 
0.944444444444 -0.020202020202 0 -1.2 1e-06 
1.0 -0.020202020202 0 -1.2 1e-06 
0.5 0.020202020202 0 -1.2 1e-06 
0.555555555556 0.020202020202 0 -1.2 1e-06 
0.611111111111 0.020202020202 0 -1.2 1e-06 
0.666666666667 0.020202020202 0 -1.2 1e-06 
0.722222222222 0.020202020202 0 -1.2 1e-06 
0.777777777778 0.020202020202 0 -1.2 1e-06 
0.833333333333 0.020202020202 0 -1.2 1e-06 
0.888888888889 0.020202020202 0 -1.2 1e-06 
0.944444444444 0.020202020202 0 -1.2 1e-06 
1.0 0.020202020202 0 -1.2 1e-06 
0.5 0.0606060606061 0 -1.2 1e-06 
0.555555555556 0.0606060606061 0 -1.2 1e-06 
0.611111111111 0.0606060606061 0 -1.2 1e-06 
0.666666666667 0.0606060606061 0 -1.2 1e-06 
0.722222222222 0.0606060606061 0 -1.2 1e-06 
0.777777777778 0.0606060606061 0 -1.2 1e-06 
0.833333333333 0.0606060606061 0 -1.2 1e-06 
0.888888888889 0.0606060606061 0 -1.2 1e-06 
0.944444444444 0.0606060606061 0 -1.2 1e-06 
1.0 0.0606060606061 0 -1.2 1e-06 
0.5 0.10101010101 0 -1.2 1e-06 
0.555555555556 0.10101010101 0 -1.2 1e-06 
0.611111111111 0.10101010101 0 -1.2 1e-06 
0.666666666667 0.10101010101 0 -1.2 1e-06 
0.722222222222 0.10101010101 0 -1.2 1e-06 
0.777777777778 0.10101010101 0 -1.2 1e-06 
0.833333333333 0.10101010101 0 -1.2 1e-06 
0.888888888889 0.10101010101 0 -1.2 1e-06 
0.944444444444 0.10101010101 0 -1.2 1e-06 
1.0 0.10101010101 0 -1.2 1e-06 
0.5 0.141414141414 0 -1.2 1e-06 
0.555555555556 0.141414141414 0 -1.2 1e-06 
0.611111111111 0.141414141414 0 -1.2 1e-06 
0.666666666667 0.141414141414 0 -1.2 1e-06 
0.722222222222 0.141414141414 0 -1.2 1e-06 
0.777777777778 0.141414141414 0 -1.2 1e-06 
0.833333333333 0.141414141414 0 -1.2 1e-06 
0.888888888889 0.141414141414 0 -1.2 1e-06 
0.944444444444 0.141414141414 0 -1.2 1e-06 
1.0 0.141414141414 0 -1.2 1e-06 
0.5 0.181818181818 0 -1.2 1e-06 
0.555555555556 0.181818181818 0 -1.2 1e-06 
0.611111111111 0.181818181818 0 -1.2 1e-06 
0.666666666667 0.181818181818 0 -1.2 1e-06 
0.722222222222 0.181818181818 0 -1.2 1e-06 
0.777777777778 0.181818181818 0 -1.2 1e-06 
0.833333333333 0.181818181818 0 -1.2 1e-06 
0.888888888889 0.181818181818 0 -1.2 1e-06 
0.944444444444 0.181818181818 0 -1.2 1e-06 
1.0 0.181818181818 0 -1.2 1e-06 
0.5 0.222222222222 0 -1.2 1e-06 
0.555555555556 0.222222222222 0 -1.2 1e-06 
0.611111111111 0.222222222222 0 -1.2 1e-06 
0.666666666667 0.222222222222 0 -1.2 1e-06 
0.722222222222 0.222222222222 0 -1.2 1e-06 
0.777777777778 0.222222222222 0 -1.2 1e-06 
0.833333333333 0.222222222222 0 -1.2 1e-06 
0.888888888889 0.222222222222 0 -1.2 1e-06 
0.944444444444 0.222222222222 0 -1.2 1e-06 
1.0 0.222222222222 0 -1.2 1e-06 
0.5 0.262626262626 0 -1.2 1e-06 
0.555555555556 0.262626262626 0 -1.2 1e-06 
0.611111111111 0.262626262626 0 -1.2 1e-06 
0.666666666667 0.262626262626 0 -1.2 1e-06 
0.722222222222 0.262626262626 0 -1.2 1e-06 
0.777777777778 0.262626262626 0 -1.2 1e-06 
0.833333333333 0.262626262626 0 -1.2 1e-06 
0.888888888889 0.262626262626 0 -1.2 1e-06 
0.944444444444 0.262626262626 0 -1.2 1e-06 
1.0 0.262626262626 0 -1.2 1e-06 
0.5 0.30303030303 0 -1.2 1e-06 
0.555555555556 0.30303030303 0 -1.2 1e-06 
0.611111111111 0.30303030303 0 -1.2 1e-06 
0.666666666667 0.30303030303 0 -1.2 1e-06 
0.722222222222 0.30303030303 0 -1.2 1e-06 
0.777777777778 0.30303030303 0 -1.2 1e-06 
0.833333333333 0.30303030303 0 -1.2 1e-06 
0.888888888889 0.30303030303 0 -1.2 1e-06 
0.944444444444 0.30303030303 0 -1.2 1e-06 
1.0 0.30303030303 0 -1.2 1e-06 
0.5 0.343434343434 0 -1.2 1e-06 
0.555555555556 0.343434343434 0 -1.2 1e-06 
0.611111111111 0.343434343434 0 -1.2 1e-06 
0.666666666667 0.343434343434 0 -1.2 1e-06 
0.722222222222 0.343434343434 0 -1.2 1e-06 
0.777777777778 0.343434343434 0 -1.2 1e-06 
0.833333333333 0.343434343434 0 -1.2 1e-06 
0.888888888889 0.343434343434 0 -1.2 1e-06 
0.944444444444 0.343434343434 0 -1.2 1e-06 
1.0 0.343434343434 0 -1.2 1e-06 
0.5 0.383838383838 0 -1.2 1e-06 
0.555555555556 0.383838383838 0 -1.2 1e-06 
0.611111111111 0.383838383838 0 -1.2 1e-06 
0.666666666667 0.383838383838 0 -1.2 1e-06 
0.722222222222 0.383838383838 0 -1.2 1e-06 
0.777777777778 0.383838383838 0 -1.2 1e-06 
0.833333333333 0.383838383838 0 -1.2 1e-06 
0.888888888889 0.383838383838 0 -1.2 1e-06 
0.944444444444 0.383838383838 0 -1.2 1e-06 
1.0 0.383838383838 0 -1.2 1e-06 
0.5 0.424242424242 0 -1.2 1e-06 
0.555555555556 0.424242424242 0 -1.2 1e-06 
0.611111111111 0.424242424242 0 -1.2 1e-06 
0.666666666667 0.424242424242 0 -1.2 1e-06 
0.722222222222 0.424242424242 0 -1.2 1e-06 
0.777777777778 0.424242424242 0 -1.2 1e-06 
0.833333333333 0.424242424242 0 -1.2 1e-06 
0.888888888889 0.424242424242 0 -1.2 1e-06 
0.944444444444 0.424242424242 0 -1.2 1e-06 
1.0 0.424242424242 0 -1.2 1e-06 
0.5 0.464646464646 0 -1.2 1e-06 
0.555555555556 0.464646464646 0 -1.2 1e-06 
0.611111111111 0.464646464646 0 -1.2 1e-06 
0.666666666667 0.464646464646 0 -1.2 1e-06 
0.722222222222 0.464646464646 0 -1.2 1e-06 
0.777777777778 0.464646464646 0 -1.2 1e-06 
0.833333333333 0.464646464646 0 -1.2 1e-06 
0.888888888889 0.464646464646 0 -1.2 1e-06 
0.944444444444 0.464646464646 0 -1.2 1e-06 
1.0 0.464646464646 0 -1.2 1e-06 
0.5 0.505050505051 0 -1.2 1e-06 
0.555555555556 0.505050505051 0 -1.2 1e-06 
0.611111111111 0.505050505051 0 -1.2 1e-06 
0.666666666667 0.505050505051 0 -1.2 1e-06 
0.722222222222 0.505050505051 0 -1.2 1e-06 
0.777777777778 0.505050505051 0 -1.2 1e-06 
0.833333333333 0.505050505051 0 -1.2 1e-06 
0.888888888889 0.505050505051 0 -1.2 1e-06 
0.944444444444 0.505050505051 0 -1.2 1e-06 
1.0 0.505050505051 0 -1.2 1e-06 
0.5 0.545454545455 0 -1.2 1e-06 
0.555555555556 0.545454545455 0 -1.2 1e-06 
0.611111111111 0.545454545455 0 -1.2 1e-06 
0.666666666667 0.545454545455 0 -1.2 1e-06 
0.722222222222 0.545454545455 0 -1.2 1e-06 
0.777777777778 0.545454545455 0 -1.2 1e-06 
0.833333333333 0.545454545455 0 -1.2 1e-06 
0.888888888889 0.545454545455 0 -1.2 1e-06 
0.944444444444 0.545454545455 0 -1.2 1e-06 
1.0 0.545454545455 0 -1.2 1e-06 
0.5 0.585858585859 0 -1.2 1e-06 
0.555555555556 0.585858585859 0 -1.2 1e-06 
0.611111111111 0.585858585859 0 -1.2 1e-06 
0.666666666667 0.585858585859 0 -1.2 1e-06 
0.722222222222 0.585858585859 0 -1.2 1e-06 
0.777777777778 0.585858585859 0 -1.2 1e-06 
0.833333333333 0.585858585859 0 -1.2 1e-06 
0.888888888889 0.585858585859 0 -1.2 1e-06 
0.944444444444 0.585858585859 0 -1.2 1e-06 
1.0 0.585858585859 0 -1.2 1e-06 
0.5 0.626262626263 0 -1.2 1e-06 
0.555555555556 0.626262626263 0 -1.2 1e-06 
0.611111111111 0.626262626263 0 -1.2 1e-06 
0.666666666667 0.626262626263 0 -1.2 1e-06 
0.722222222222 0.626262626263 0 -1.2 1e-06 
0.777777777778 0.626262626263 0 -1.2 1e-06 
0.833333333333 0.626262626263 0 -1.2 1e-06 
0.888888888889 0.626262626263 0 -1.2 1e-06 
0.944444444444 0.626262626263 0 -1.2 1e-06 
1.0 0.626262626263 0 -1.2 1e-06 
0.5 0.666666666667 0 -1.2 1e-06 
0.555555555556 0.666666666667 0 -1.2 1e-06 
0.611111111111 0.666666666667 0 -1.2 1e-06 
0.666666666667 0.666666666667 0 -1.2 1e-06 
0.722222222222 0.666666666667 0 -1.2 1e-06 
0.777777777778 0.666666666667 0 -1.2 1e-06 
0.833333333333 0.666666666667 0 -1.2 1e-06 
0.888888888889 0.666666666667 0 -1.2 1e-06 
0.944444444444 0.666666666667 0 -1.2 1e-06 
1.0 0.666666666667 0 -1.2 1e-06 
0.5 0.707070707071 0 -1.2 1e-06 
0.555555555556 0.707070707071 0 -1.2 1e-06 
0.611111111111 0.707070707071 0 -1.2 1e-06 
0.666666666667 0.707070707071 0 -1.2 1e-06 
0.722222222222 0.707070707071 0 -1.2 1e-06 
0.777777777778 0.707070707071 0 -1.2 1e-06 
0.833333333333 0.707070707071 0 -1.2 1e-06 
0.888888888889 0.707070707071 0 -1.2 1e-06 
0.944444444444 0.707070707071 0 -1.2 1e-06 
1.0 0.707070707071 0 -1.2 1e-06 
0.5 0.747474747475 0 -1.2 1e-06 
0.555555555556 0.747474747475 0 -1.2 1e-06 
0.611111111111 0.747474747475 0 -1.2 1e-06 
0.666666666667 0.747474747475 0 -1.2 1e-06 
0.722222222222 0.747474747475 0 -1.2 1e-06 
0.777777777778 0.747474747475 0 -1.2 1e-06 
0.833333333333 0.747474747475 0 -1.2 1e-06 
0.888888888889 0.747474747475 0 -1.2 1e-06 
0.944444444444 0.747474747475 0 -1.2 1e-06 
1.0 0.747474747475 0 -1.2 1e-06 
0.5 0.787878787879 0 -1.2 1e-06 
0.555555555556 0.787878787879 0 -1.2 1e-06 
0.611111111111 0.787878787879 0 -1.2 1e-06 
0.666666666667 0.787878787879 0 -1.2 1e-06 
0.722222222222 0.787878787879 0 -1.2 1e-06 
0.777777777778 0.787878787879 0 -1.2 1e-06 
0.833333333333 0.787878787879 0 -1.2 1e-06 
0.888888888889 0.787878787879 0 -1.2 1e-06 
0.944444444444 0.787878787879 0 -1.2 1e-06 
1.0 0.787878787879 0 -1.2 1e-06 
0.5 0.828282828283 0 -1.2 1e-06 
0.555555555556 0.828282828283 0 -1.2 1e-06 
0.611111111111 0.828282828283 0 -1.2 1e-06 
0.666666666667 0.828282828283 0 -1.2 1e-06 
0.722222222222 0.828282828283 0 -1.2 1e-06 
0.777777777778 0.828282828283 0 -1.2 1e-06 
0.833333333333 0.828282828283 0 -1.2 1e-06 
0.888888888889 0.828282828283 0 -1.2 1e-06 
0.944444444444 0.828282828283 0 -1.2 1e-06 
1.0 0.828282828283 0 -1.2 1e-06 
0.5 0.868686868687 0 -1.2 1e-06 
0.555555555556 0.868686868687 0 -1.2 1e-06 
0.611111111111 0.868686868687 0 -1.2 1e-06 
0.666666666667 0.868686868687 0 -1.2 1e-06 
0.722222222222 0.868686868687 0 -1.2 1e-06 
0.777777777778 0.868686868687 0 -1.2 1e-06 
0.833333333333 0.868686868687 0 -1.2 1e-06 
0.888888888889 0.868686868687 0 -1.2 1e-06 
0.944444444444 0.868686868687 0 -1.2 1e-06 
1.0 0.868686868687 0 -1.2 1e-06 
0.5 0.909090909091 0 -1.2 1e-06 
0.555555555556 0.909090909091 0 -1.2 1e-06 
0.611111111111 0.909090909091 0 -1.2 1e-06 
0.666666666667 0.909090909091 0 -1.2 1e-06 
0.722222222222 0.909090909091 0 -1.2 1e-06 
0.777777777778 0.909090909091 0 -1.2 1e-06 
0.833333333333 0.909090909091 0 -1.2 1e-06 
0.888888888889 0.909090909091 0 -1.2 1e-06 
0.944444444444 0.909090909091 0 -1.2 1e-06 
1.0 0.909090909091 0 -1.2 1e-06 
0.5 0.949494949495 0 -1.2 1e-06 
0.555555555556 0.949494949495 0 -1.2 1e-06 
0.611111111111 0.949494949495 0 -1.2 1e-06 
0.666666666667 0.949494949495 0 -1.2 1e-06 
0.722222222222 0.949494949495 0 -1.2 1e-06 
0.777777777778 0.949494949495 0 -1.2 1e-06 
0.833333333333 0.949494949495 0 -1.2 1e-06 
0.888888888889 0.949494949495 0 -1.2 1e-06 
0.944444444444 0.949494949495 0 -1.2 1e-06 
1.0 0.949494949495 0 -1.2 1e-06 
0.5 0.989898989899 0 -1.2 1e-06 
0.555555555556 0.989898989899 0 -1.2 1e-06 
0.611111111111 0.989898989899 0 -1.2 1e-06 
0.666666666667 0.989898989899 0 -1.2 1e-06 
0.722222222222 0.989898989899 0 -1.2 1e-06 
0.777777777778 0.989898989899 0 -1.2 1e-06 
0.833333333333 0.989898989899 0 -1.2 1e-06 
0.888888888889 0.989898989899 0 -1.2 1e-06 
0.944444444444 0.989898989899 0 -1.2 1e-06 
1.0 0.989898989899 0 -1.2 1e-06 
0.5 1.0303030303 0 -1.2 1e-06 
0.555555555556 1.0303030303 0 -1.2 1e-06 
0.611111111111 1.0303030303 0 -1.2 1e-06 
0.666666666667 1.0303030303 0 -1.2 1e-06 
0.722222222222 1.0303030303 0 -1.2 1e-06 
0.777777777778 1.0303030303 0 -1.2 1e-06 
0.833333333333 1.0303030303 0 -1.2 1e-06 
0.888888888889 1.0303030303 0 -1.2 1e-06 
0.944444444444 1.0303030303 0 -1.2 1e-06 
1.0 1.0303030303 0 -1.2 1e-06 
0.5 1.07070707071 0 -1.2 1e-06 
0.555555555556 1.07070707071 0 -1.2 1e-06 
0.611111111111 1.07070707071 0 -1.2 1e-06 
0.666666666667 1.07070707071 0 -1.2 1e-06 
0.722222222222 1.07070707071 0 -1.2 1e-06 
0.777777777778 1.07070707071 0 -1.2 1e-06 
0.833333333333 1.07070707071 0 -1.2 1e-06 
0.888888888889 1.07070707071 0 -1.2 1e-06 
0.944444444444 1.07070707071 0 -1.2 1e-06 
1.0 1.07070707071 0 -1.2 1e-06 
0.5 1.11111111111 0 -1.2 1e-06 
0.555555555556 1.11111111111 0 -1.2 1e-06 
0.611111111111 1.11111111111 0 -1.2 1e-06 
0.666666666667 1.11111111111 0 -1.2 1e-06 
0.722222222222 1.11111111111 0 -1.2 1e-06 
0.777777777778 1.11111111111 0 -1.2 1e-06 
0.833333333333 1.11111111111 0 -1.2 1e-06 
0.888888888889 1.11111111111 0 -1.2 1e-06 
0.944444444444 1.11111111111 0 -1.2 1e-06 
1.0 1.11111111111 0 -1.2 1e-06 
0.5 1.15151515152 0 -1.2 1e-06 
0.555555555556 1.15151515152 0 -1.2 1e-06 
0.611111111111 1.15151515152 0 -1.2 1e-06 
0.666666666667 1.15151515152 0 -1.2 1e-06 
0.722222222222 1.15151515152 0 -1.2 1e-06 
0.777777777778 1.15151515152 0 -1.2 1e-06 
0.833333333333 1.15151515152 0 -1.2 1e-06 
0.888888888889 1.15151515152 0 -1.2 1e-06 
0.944444444444 1.15151515152 0 -1.2 1e-06 
1.0 1.15151515152 0 -1.2 1e-06 
0.5 1.19191919192 0 -1.2 1e-06 
0.555555555556 1.19191919192 0 -1.2 1e-06 
0.611111111111 1.19191919192 0 -1.2 1e-06 
0.666666666667 1.19191919192 0 -1.2 1e-06 
0.722222222222 1.19191919192 0 -1.2 1e-06 
0.777777777778 1.19191919192 0 -1.2 1e-06 
0.833333333333 1.19191919192 0 -1.2 1e-06 
0.888888888889 1.19191919192 0 -1.2 1e-06 
0.944444444444 1.19191919192 0 -1.2 1e-06 
1.0 1.19191919192 0 -1.2 1e-06 
0.5 1.23232323232 0 -1.2 1e-06 
0.555555555556 1.23232323232 0 -1.2 1e-06 
0.611111111111 1.23232323232 0 -1.2 1e-06 
0.666666666667 1.23232323232 0 -1.2 1e-06 
0.722222222222 1.23232323232 0 -1.2 1e-06 
0.777777777778 1.23232323232 0 -1.2 1e-06 
0.833333333333 1.23232323232 0 -1.2 1e-06 
0.888888888889 1.23232323232 0 -1.2 1e-06 
0.944444444444 1.23232323232 0 -1.2 1e-06 
1.0 1.23232323232 0 -1.2 1e-06 
0.5 1.27272727273 0 -1.2 1e-06 
0.555555555556 1.27272727273 0 -1.2 1e-06 
0.611111111111 1.27272727273 0 -1.2 1e-06 
0.666666666667 1.27272727273 0 -1.2 1e-06 
0.722222222222 1.27272727273 0 -1.2 1e-06 
0.777777777778 1.27272727273 0 -1.2 1e-06 
0.833333333333 1.27272727273 0 -1.2 1e-06 
0.888888888889 1.27272727273 0 -1.2 1e-06 
0.944444444444 1.27272727273 0 -1.2 1e-06 
1.0 1.27272727273 0 -1.2 1e-06 
0.5 1.31313131313 0 -1.2 1e-06 
0.555555555556 1.31313131313 0 -1.2 1e-06 
0.611111111111 1.31313131313 0 -1.2 1e-06 
0.666666666667 1.31313131313 0 -1.2 1e-06 
0.722222222222 1.31313131313 0 -1.2 1e-06 
0.777777777778 1.31313131313 0 -1.2 1e-06 
0.833333333333 1.31313131313 0 -1.2 1e-06 
0.888888888889 1.31313131313 0 -1.2 1e-06 
0.944444444444 1.31313131313 0 -1.2 1e-06 
1.0 1.31313131313 0 -1.2 1e-06 
0.5 1.35353535354 0 -1.2 1e-06 
0.555555555556 1.35353535354 0 -1.2 1e-06 
0.611111111111 1.35353535354 0 -1.2 1e-06 
0.666666666667 1.35353535354 0 -1.2 1e-06 
0.722222222222 1.35353535354 0 -1.2 1e-06 
0.777777777778 1.35353535354 0 -1.2 1e-06 
0.833333333333 1.35353535354 0 -1.2 1e-06 
0.888888888889 1.35353535354 0 -1.2 1e-06 
0.944444444444 1.35353535354 0 -1.2 1e-06 
1.0 1.35353535354 0 -1.2 1e-06 
0.5 1.39393939394 0 -1.2 1e-06 
0.555555555556 1.39393939394 0 -1.2 1e-06 
0.611111111111 1.39393939394 0 -1.2 1e-06 
0.666666666667 1.39393939394 0 -1.2 1e-06 
0.722222222222 1.39393939394 0 -1.2 1e-06 
0.777777777778 1.39393939394 0 -1.2 1e-06 
0.833333333333 1.39393939394 0 -1.2 1e-06 
0.888888888889 1.39393939394 0 -1.2 1e-06 
0.944444444444 1.39393939394 0 -1.2 1e-06 
1.0 1.39393939394 0 -1.2 1e-06 
0.5 1.43434343434 0 -1.2 1e-06 
0.555555555556 1.43434343434 0 -1.2 1e-06 
0.611111111111 1.43434343434 0 -1.2 1e-06 
0.666666666667 1.43434343434 0 -1.2 1e-06 
0.722222222222 1.43434343434 0 -1.2 1e-06 
0.777777777778 1.43434343434 0 -1.2 1e-06 
0.833333333333 1.43434343434 0 -1.2 1e-06 
0.888888888889 1.43434343434 0 -1.2 1e-06 
0.944444444444 1.43434343434 0 -1.2 1e-06 
1.0 1.43434343434 0 -1.2 1e-06 
0.5 1.47474747475 0 -1.2 1e-06 
0.555555555556 1.47474747475 0 -1.2 1e-06 
0.611111111111 1.47474747475 0 -1.2 1e-06 
0.666666666667 1.47474747475 0 -1.2 1e-06 
0.722222222222 1.47474747475 0 -1.2 1e-06 
0.777777777778 1.47474747475 0 -1.2 1e-06 
0.833333333333 1.47474747475 0 -1.2 1e-06 
0.888888888889 1.47474747475 0 -1.2 1e-06 
0.944444444444 1.47474747475 0 -1.2 1e-06 
1.0 1.47474747475 0 -1.2 1e-06 
0.5 1.51515151515 0 -1.2 1e-06 
0.555555555556 1.51515151515 0 -1.2 1e-06 
0.611111111111 1.51515151515 0 -1.2 1e-06 
0.666666666667 1.51515151515 0 -1.2 1e-06 
0.722222222222 1.51515151515 0 -1.2 1e-06 
0.777777777778 1.51515151515 0 -1.2 1e-06 
0.833333333333 1.51515151515 0 -1.2 1e-06 
0.888888888889 1.51515151515 0 -1.2 1e-06 
0.944444444444 1.51515151515 0 -1.2 1e-06 
1.0 1.51515151515 0 -1.2 1e-06 
0.5 1.55555555556 0 -1.2 1e-06 
0.555555555556 1.55555555556 0 -1.2 1e-06 
0.611111111111 1.55555555556 0 -1.2 1e-06 
0.666666666667 1.55555555556 0 -1.2 1e-06 
0.722222222222 1.55555555556 0 -1.2 1e-06 
0.777777777778 1.55555555556 0 -1.2 1e-06 
0.833333333333 1.55555555556 0 -1.2 1e-06 
0.888888888889 1.55555555556 0 -1.2 1e-06 
0.944444444444 1.55555555556 0 -1.2 1e-06 
1.0 1.55555555556 0 -1.2 1e-06 
0.5 1.59595959596 0 -1.2 1e-06 
0.555555555556 1.59595959596 0 -1.2 1e-06 
0.611111111111 1.59595959596 0 -1.2 1e-06 
0.666666666667 1.59595959596 0 -1.2 1e-06 
0.722222222222 1.59595959596 0 -1.2 1e-06 
0.777777777778 1.59595959596 0 -1.2 1e-06 
0.833333333333 1.59595959596 0 -1.2 1e-06 
0.888888888889 1.59595959596 0 -1.2 1e-06 
0.944444444444 1.59595959596 0 -1.2 1e-06 
1.0 1.59595959596 0 -1.2 1e-06 
0.5 1.63636363636 0 -1.2 1e-06 
0.555555555556 1.63636363636 0 -1.2 1e-06 
0.611111111111 1.63636363636 0 -1.2 1e-06 
0.666666666667 1.63636363636 0 -1.2 1e-06 
0.722222222222 1.63636363636 0 -1.2 1e-06 
0.777777777778 1.63636363636 0 -1.2 1e-06 
0.833333333333 1.63636363636 0 -1.2 1e-06 
0.888888888889 1.63636363636 0 -1.2 1e-06 
0.944444444444 1.63636363636 0 -1.2 1e-06 
1.0 1.63636363636 0 -1.2 1e-06 
0.5 1.67676767677 0 -1.2 1e-06 
0.555555555556 1.67676767677 0 -1.2 1e-06 
0.611111111111 1.67676767677 0 -1.2 1e-06 
0.666666666667 1.67676767677 0 -1.2 1e-06 
0.722222222222 1.67676767677 0 -1.2 1e-06 
0.777777777778 1.67676767677 0 -1.2 1e-06 
0.833333333333 1.67676767677 0 -1.2 1e-06 
0.888888888889 1.67676767677 0 -1.2 1e-06 
0.944444444444 1.67676767677 0 -1.2 1e-06 
1.0 1.67676767677 0 -1.2 1e-06 
0.5 1.71717171717 0 -1.2 1e-06 
0.555555555556 1.71717171717 0 -1.2 1e-06 
0.611111111111 1.71717171717 0 -1.2 1e-06 
0.666666666667 1.71717171717 0 -1.2 1e-06 
0.722222222222 1.71717171717 0 -1.2 1e-06 
0.777777777778 1.71717171717 0 -1.2 1e-06 
0.833333333333 1.71717171717 0 -1.2 1e-06 
0.888888888889 1.71717171717 0 -1.2 1e-06 
0.944444444444 1.71717171717 0 -1.2 1e-06 
1.0 1.71717171717 0 -1.2 1e-06 
0.5 1.75757575758 0 -1.2 1e-06 
0.555555555556 1.75757575758 0 -1.2 1e-06 
0.611111111111 1.75757575758 0 -1.2 1e-06 
0.666666666667 1.75757575758 0 -1.2 1e-06 
0.722222222222 1.75757575758 0 -1.2 1e-06 
0.777777777778 1.75757575758 0 -1.2 1e-06 
0.833333333333 1.75757575758 0 -1.2 1e-06 
0.888888888889 1.75757575758 0 -1.2 1e-06 
0.944444444444 1.75757575758 0 -1.2 1e-06 
1.0 1.75757575758 0 -1.2 1e-06 
0.5 1.79797979798 0 -1.2 1e-06 
0.555555555556 1.79797979798 0 -1.2 1e-06 
0.611111111111 1.79797979798 0 -1.2 1e-06 
0.666666666667 1.79797979798 0 -1.2 1e-06 
0.722222222222 1.79797979798 0 -1.2 1e-06 
0.777777777778 1.79797979798 0 -1.2 1e-06 
0.833333333333 1.79797979798 0 -1.2 1e-06 
0.888888888889 1.79797979798 0 -1.2 1e-06 
0.944444444444 1.79797979798 0 -1.2 1e-06 
1.0 1.79797979798 0 -1.2 1e-06 
0.5 1.83838383838 0 -1.2 1e-06 
0.555555555556 1.83838383838 0 -1.2 1e-06 
0.611111111111 1.83838383838 0 -1.2 1e-06 
0.666666666667 1.83838383838 0 -1.2 1e-06 
0.722222222222 1.83838383838 0 -1.2 1e-06 
0.777777777778 1.83838383838 0 -1.2 1e-06 
0.833333333333 1.83838383838 0 -1.2 1e-06 
0.888888888889 1.83838383838 0 -1.2 1e-06 
0.944444444444 1.83838383838 0 -1.2 1e-06 
1.0 1.83838383838 0 -1.2 1e-06 
0.5 1.87878787879 0 -1.2 1e-06 
0.555555555556 1.87878787879 0 -1.2 1e-06 
0.611111111111 1.87878787879 0 -1.2 1e-06 
0.666666666667 1.87878787879 0 -1.2 1e-06 
0.722222222222 1.87878787879 0 -1.2 1e-06 
0.777777777778 1.87878787879 0 -1.2 1e-06 
0.833333333333 1.87878787879 0 -1.2 1e-06 
0.888888888889 1.87878787879 0 -1.2 1e-06 
0.944444444444 1.87878787879 0 -1.2 1e-06 
1.0 1.87878787879 0 -1.2 1e-06 
0.5 1.91919191919 0 -1.2 1e-06 
0.555555555556 1.91919191919 0 -1.2 1e-06 
0.611111111111 1.91919191919 0 -1.2 1e-06 
0.666666666667 1.91919191919 0 -1.2 1e-06 
0.722222222222 1.91919191919 0 -1.2 1e-06 
0.777777777778 1.91919191919 0 -1.2 1e-06 
0.833333333333 1.91919191919 0 -1.2 1e-06 
0.888888888889 1.91919191919 0 -1.2 1e-06 
0.944444444444 1.91919191919 0 -1.2 1e-06 
1.0 1.91919191919 0 -1.2 1e-06 
0.5 1.9595959596 0 -1.2 1e-06 
0.555555555556 1.9595959596 0 -1.2 1e-06 
0.611111111111 1.9595959596 0 -1.2 1e-06 
0.666666666667 1.9595959596 0 -1.2 1e-06 
0.722222222222 1.9595959596 0 -1.2 1e-06 
0.777777777778 1.9595959596 0 -1.2 1e-06 
0.833333333333 1.9595959596 0 -1.2 1e-06 
0.888888888889 1.9595959596 0 -1.2 1e-06 
0.944444444444 1.9595959596 0 -1.2 1e-06 
1.0 1.9595959596 0 -1.2 1e-06 
0.5 2.0 0 -1.2 1e-06 
0.555555555556 2.0 0 -1.2 1e-06 
0.611111111111 2.0 0 -1.2 1e-06 
0.666666666667 2.0 0 -1.2 1e-06 
0.722222222222 2.0 0 -1.2 1e-06 
0.777777777778 2.0 0 -1.2 1e-06 
0.833333333333 2.0 0 -1.2 1e-06 
0.888888888889 2.0 0 -1.2 1e-06 
0.944444444444 2.0 0 -1.2 1e-06 
1.0 2.0 0 -1.2 1e-06 
0.5 -2.0 0 -0.8 1e-06 
0.555555555556 -2.0 0 -0.8 1e-06 
0.611111111111 -2.0 0 -0.8 1e-06 
0.666666666667 -2.0 0 -0.8 1e-06 
0.722222222222 -2.0 0 -0.8 1e-06 
0.777777777778 -2.0 0 -0.8 1e-06 
0.833333333333 -2.0 0 -0.8 1e-06 
0.888888888889 -2.0 0 -0.8 1e-06 
0.944444444444 -2.0 0 -0.8 1e-06 
1.0 -2.0 0 -0.8 1e-06 
0.5 -1.9595959596 0 -0.8 1e-06 
0.555555555556 -1.9595959596 0 -0.8 1e-06 
0.611111111111 -1.9595959596 0 -0.8 1e-06 
0.666666666667 -1.9595959596 0 -0.8 1e-06 
0.722222222222 -1.9595959596 0 -0.8 1e-06 
0.777777777778 -1.9595959596 0 -0.8 1e-06 
0.833333333333 -1.9595959596 0 -0.8 1e-06 
0.888888888889 -1.9595959596 0 -0.8 1e-06 
0.944444444444 -1.9595959596 0 -0.8 1e-06 
1.0 -1.9595959596 0 -0.8 1e-06 
0.5 -1.91919191919 0 -0.8 1e-06 
0.555555555556 -1.91919191919 0 -0.8 1e-06 
0.611111111111 -1.91919191919 0 -0.8 1e-06 
0.666666666667 -1.91919191919 0 -0.8 1e-06 
0.722222222222 -1.91919191919 0 -0.8 1e-06 
0.777777777778 -1.91919191919 0 -0.8 1e-06 
0.833333333333 -1.91919191919 0 -0.8 1e-06 
0.888888888889 -1.91919191919 0 -0.8 1e-06 
0.944444444444 -1.91919191919 0 -0.8 1e-06 
1.0 -1.91919191919 0 -0.8 1e-06 
0.5 -1.87878787879 0 -0.8 1e-06 
0.555555555556 -1.87878787879 0 -0.8 1e-06 
0.611111111111 -1.87878787879 0 -0.8 1e-06 
0.666666666667 -1.87878787879 0 -0.8 1e-06 
0.722222222222 -1.87878787879 0 -0.8 1e-06 
0.777777777778 -1.87878787879 0 -0.8 1e-06 
0.833333333333 -1.87878787879 0 -0.8 1e-06 
0.888888888889 -1.87878787879 0 -0.8 1e-06 
0.944444444444 -1.87878787879 0 -0.8 1e-06 
1.0 -1.87878787879 0 -0.8 1e-06 
0.5 -1.83838383838 0 -0.8 1e-06 
0.555555555556 -1.83838383838 0 -0.8 1e-06 
0.611111111111 -1.83838383838 0 -0.8 1e-06 
0.666666666667 -1.83838383838 0 -0.8 1e-06 
0.722222222222 -1.83838383838 0 -0.8 1e-06 
0.777777777778 -1.83838383838 0 -0.8 1e-06 
0.833333333333 -1.83838383838 0 -0.8 1e-06 
0.888888888889 -1.83838383838 0 -0.8 1e-06 
0.944444444444 -1.83838383838 0 -0.8 1e-06 
1.0 -1.83838383838 0 -0.8 1e-06 
0.5 -1.79797979798 0 -0.8 1e-06 
0.555555555556 -1.79797979798 0 -0.8 1e-06 
0.611111111111 -1.79797979798 0 -0.8 1e-06 
0.666666666667 -1.79797979798 0 -0.8 1e-06 
0.722222222222 -1.79797979798 0 -0.8 1e-06 
0.777777777778 -1.79797979798 0 -0.8 1e-06 
0.833333333333 -1.79797979798 0 -0.8 1e-06 
0.888888888889 -1.79797979798 0 -0.8 1e-06 
0.944444444444 -1.79797979798 0 -0.8 1e-06 
1.0 -1.79797979798 0 -0.8 1e-06 
0.5 -1.75757575758 0 -0.8 1e-06 
0.555555555556 -1.75757575758 0 -0.8 1e-06 
0.611111111111 -1.75757575758 0 -0.8 1e-06 
0.666666666667 -1.75757575758 0 -0.8 1e-06 
0.722222222222 -1.75757575758 0 -0.8 1e-06 
0.777777777778 -1.75757575758 0 -0.8 1e-06 
0.833333333333 -1.75757575758 0 -0.8 1e-06 
0.888888888889 -1.75757575758 0 -0.8 1e-06 
0.944444444444 -1.75757575758 0 -0.8 1e-06 
1.0 -1.75757575758 0 -0.8 1e-06 
0.5 -1.71717171717 0 -0.8 1e-06 
0.555555555556 -1.71717171717 0 -0.8 1e-06 
0.611111111111 -1.71717171717 0 -0.8 1e-06 
0.666666666667 -1.71717171717 0 -0.8 1e-06 
0.722222222222 -1.71717171717 0 -0.8 1e-06 
0.777777777778 -1.71717171717 0 -0.8 1e-06 
0.833333333333 -1.71717171717 0 -0.8 1e-06 
0.888888888889 -1.71717171717 0 -0.8 1e-06 
0.944444444444 -1.71717171717 0 -0.8 1e-06 
1.0 -1.71717171717 0 -0.8 1e-06 
0.5 -1.67676767677 0 -0.8 1e-06 
0.555555555556 -1.67676767677 0 -0.8 1e-06 
0.611111111111 -1.67676767677 0 -0.8 1e-06 
0.666666666667 -1.67676767677 0 -0.8 1e-06 
0.722222222222 -1.67676767677 0 -0.8 1e-06 
0.777777777778 -1.67676767677 0 -0.8 1e-06 
0.833333333333 -1.67676767677 0 -0.8 1e-06 
0.888888888889 -1.67676767677 0 -0.8 1e-06 
0.944444444444 -1.67676767677 0 -0.8 1e-06 
1.0 -1.67676767677 0 -0.8 1e-06 
0.5 -1.63636363636 0 -0.8 1e-06 
0.555555555556 -1.63636363636 0 -0.8 1e-06 
0.611111111111 -1.63636363636 0 -0.8 1e-06 
0.666666666667 -1.63636363636 0 -0.8 1e-06 
0.722222222222 -1.63636363636 0 -0.8 1e-06 
0.777777777778 -1.63636363636 0 -0.8 1e-06 
0.833333333333 -1.63636363636 0 -0.8 1e-06 
0.888888888889 -1.63636363636 0 -0.8 1e-06 
0.944444444444 -1.63636363636 0 -0.8 1e-06 
1.0 -1.63636363636 0 -0.8 1e-06 
0.5 -1.59595959596 0 -0.8 1e-06 
0.555555555556 -1.59595959596 0 -0.8 1e-06 
0.611111111111 -1.59595959596 0 -0.8 1e-06 
0.666666666667 -1.59595959596 0 -0.8 1e-06 
0.722222222222 -1.59595959596 0 -0.8 1e-06 
0.777777777778 -1.59595959596 0 -0.8 1e-06 
0.833333333333 -1.59595959596 0 -0.8 1e-06 
0.888888888889 -1.59595959596 0 -0.8 1e-06 
0.944444444444 -1.59595959596 0 -0.8 1e-06 
1.0 -1.59595959596 0 -0.8 1e-06 
0.5 -1.55555555556 0 -0.8 1e-06 
0.555555555556 -1.55555555556 0 -0.8 1e-06 
0.611111111111 -1.55555555556 0 -0.8 1e-06 
0.666666666667 -1.55555555556 0 -0.8 1e-06 
0.722222222222 -1.55555555556 0 -0.8 1e-06 
0.777777777778 -1.55555555556 0 -0.8 1e-06 
0.833333333333 -1.55555555556 0 -0.8 1e-06 
0.888888888889 -1.55555555556 0 -0.8 1e-06 
0.944444444444 -1.55555555556 0 -0.8 1e-06 
1.0 -1.55555555556 0 -0.8 1e-06 
0.5 -1.51515151515 0 -0.8 1e-06 
0.555555555556 -1.51515151515 0 -0.8 1e-06 
0.611111111111 -1.51515151515 0 -0.8 1e-06 
0.666666666667 -1.51515151515 0 -0.8 1e-06 
0.722222222222 -1.51515151515 0 -0.8 1e-06 
0.777777777778 -1.51515151515 0 -0.8 1e-06 
0.833333333333 -1.51515151515 0 -0.8 1e-06 
0.888888888889 -1.51515151515 0 -0.8 1e-06 
0.944444444444 -1.51515151515 0 -0.8 1e-06 
1.0 -1.51515151515 0 -0.8 1e-06 
0.5 -1.47474747475 0 -0.8 1e-06 
0.555555555556 -1.47474747475 0 -0.8 1e-06 
0.611111111111 -1.47474747475 0 -0.8 1e-06 
0.666666666667 -1.47474747475 0 -0.8 1e-06 
0.722222222222 -1.47474747475 0 -0.8 1e-06 
0.777777777778 -1.47474747475 0 -0.8 1e-06 
0.833333333333 -1.47474747475 0 -0.8 1e-06 
0.888888888889 -1.47474747475 0 -0.8 1e-06 
0.944444444444 -1.47474747475 0 -0.8 1e-06 
1.0 -1.47474747475 0 -0.8 1e-06 
0.5 -1.43434343434 0 -0.8 1e-06 
0.555555555556 -1.43434343434 0 -0.8 1e-06 
0.611111111111 -1.43434343434 0 -0.8 1e-06 
0.666666666667 -1.43434343434 0 -0.8 1e-06 
0.722222222222 -1.43434343434 0 -0.8 1e-06 
0.777777777778 -1.43434343434 0 -0.8 1e-06 
0.833333333333 -1.43434343434 0 -0.8 1e-06 
0.888888888889 -1.43434343434 0 -0.8 1e-06 
0.944444444444 -1.43434343434 0 -0.8 1e-06 
1.0 -1.43434343434 0 -0.8 1e-06 
0.5 -1.39393939394 0 -0.8 1e-06 
0.555555555556 -1.39393939394 0 -0.8 1e-06 
0.611111111111 -1.39393939394 0 -0.8 1e-06 
0.666666666667 -1.39393939394 0 -0.8 1e-06 
0.722222222222 -1.39393939394 0 -0.8 1e-06 
0.777777777778 -1.39393939394 0 -0.8 1e-06 
0.833333333333 -1.39393939394 0 -0.8 1e-06 
0.888888888889 -1.39393939394 0 -0.8 1e-06 
0.944444444444 -1.39393939394 0 -0.8 1e-06 
1.0 -1.39393939394 0 -0.8 1e-06 
0.5 -1.35353535354 0 -0.8 1e-06 
0.555555555556 -1.35353535354 0 -0.8 1e-06 
0.611111111111 -1.35353535354 0 -0.8 1e-06 
0.666666666667 -1.35353535354 0 -0.8 1e-06 
0.722222222222 -1.35353535354 0 -0.8 1e-06 
0.777777777778 -1.35353535354 0 -0.8 1e-06 
0.833333333333 -1.35353535354 0 -0.8 1e-06 
0.888888888889 -1.35353535354 0 -0.8 1e-06 
0.944444444444 -1.35353535354 0 -0.8 1e-06 
1.0 -1.35353535354 0 -0.8 1e-06 
0.5 -1.31313131313 0 -0.8 1e-06 
0.555555555556 -1.31313131313 0 -0.8 1e-06 
0.611111111111 -1.31313131313 0 -0.8 1e-06 
0.666666666667 -1.31313131313 0 -0.8 1e-06 
0.722222222222 -1.31313131313 0 -0.8 1e-06 
0.777777777778 -1.31313131313 0 -0.8 1e-06 
0.833333333333 -1.31313131313 0 -0.8 1e-06 
0.888888888889 -1.31313131313 0 -0.8 1e-06 
0.944444444444 -1.31313131313 0 -0.8 1e-06 
1.0 -1.31313131313 0 -0.8 1e-06 
0.5 -1.27272727273 0 -0.8 1e-06 
0.555555555556 -1.27272727273 0 -0.8 1e-06 
0.611111111111 -1.27272727273 0 -0.8 1e-06 
0.666666666667 -1.27272727273 0 -0.8 1e-06 
0.722222222222 -1.27272727273 0 -0.8 1e-06 
0.777777777778 -1.27272727273 0 -0.8 1e-06 
0.833333333333 -1.27272727273 0 -0.8 1e-06 
0.888888888889 -1.27272727273 0 -0.8 1e-06 
0.944444444444 -1.27272727273 0 -0.8 1e-06 
1.0 -1.27272727273 0 -0.8 1e-06 
0.5 -1.23232323232 0 -0.8 1e-06 
0.555555555556 -1.23232323232 0 -0.8 1e-06 
0.611111111111 -1.23232323232 0 -0.8 1e-06 
0.666666666667 -1.23232323232 0 -0.8 1e-06 
0.722222222222 -1.23232323232 0 -0.8 1e-06 
0.777777777778 -1.23232323232 0 -0.8 1e-06 
0.833333333333 -1.23232323232 0 -0.8 1e-06 
0.888888888889 -1.23232323232 0 -0.8 1e-06 
0.944444444444 -1.23232323232 0 -0.8 1e-06 
1.0 -1.23232323232 0 -0.8 1e-06 
0.5 -1.19191919192 0 -0.8 1e-06 
0.555555555556 -1.19191919192 0 -0.8 1e-06 
0.611111111111 -1.19191919192 0 -0.8 1e-06 
0.666666666667 -1.19191919192 0 -0.8 1e-06 
0.722222222222 -1.19191919192 0 -0.8 1e-06 
0.777777777778 -1.19191919192 0 -0.8 1e-06 
0.833333333333 -1.19191919192 0 -0.8 1e-06 
0.888888888889 -1.19191919192 0 -0.8 1e-06 
0.944444444444 -1.19191919192 0 -0.8 1e-06 
1.0 -1.19191919192 0 -0.8 1e-06 
0.5 -1.15151515152 0 -0.8 1e-06 
0.555555555556 -1.15151515152 0 -0.8 1e-06 
0.611111111111 -1.15151515152 0 -0.8 1e-06 
0.666666666667 -1.15151515152 0 -0.8 1e-06 
0.722222222222 -1.15151515152 0 -0.8 1e-06 
0.777777777778 -1.15151515152 0 -0.8 1e-06 
0.833333333333 -1.15151515152 0 -0.8 1e-06 
0.888888888889 -1.15151515152 0 -0.8 1e-06 
0.944444444444 -1.15151515152 0 -0.8 1e-06 
1.0 -1.15151515152 0 -0.8 1e-06 
0.5 -1.11111111111 0 -0.8 1e-06 
0.555555555556 -1.11111111111 0 -0.8 1e-06 
0.611111111111 -1.11111111111 0 -0.8 1e-06 
0.666666666667 -1.11111111111 0 -0.8 1e-06 
0.722222222222 -1.11111111111 0 -0.8 1e-06 
0.777777777778 -1.11111111111 0 -0.8 1e-06 
0.833333333333 -1.11111111111 0 -0.8 1e-06 
0.888888888889 -1.11111111111 0 -0.8 1e-06 
0.944444444444 -1.11111111111 0 -0.8 1e-06 
1.0 -1.11111111111 0 -0.8 1e-06 
0.5 -1.07070707071 0 -0.8 1e-06 
0.555555555556 -1.07070707071 0 -0.8 1e-06 
0.611111111111 -1.07070707071 0 -0.8 1e-06 
0.666666666667 -1.07070707071 0 -0.8 1e-06 
0.722222222222 -1.07070707071 0 -0.8 1e-06 
0.777777777778 -1.07070707071 0 -0.8 1e-06 
0.833333333333 -1.07070707071 0 -0.8 1e-06 
0.888888888889 -1.07070707071 0 -0.8 1e-06 
0.944444444444 -1.07070707071 0 -0.8 1e-06 
1.0 -1.07070707071 0 -0.8 1e-06 
0.5 -1.0303030303 0 -0.8 1e-06 
0.555555555556 -1.0303030303 0 -0.8 1e-06 
0.611111111111 -1.0303030303 0 -0.8 1e-06 
0.666666666667 -1.0303030303 0 -0.8 1e-06 
0.722222222222 -1.0303030303 0 -0.8 1e-06 
0.777777777778 -1.0303030303 0 -0.8 1e-06 
0.833333333333 -1.0303030303 0 -0.8 1e-06 
0.888888888889 -1.0303030303 0 -0.8 1e-06 
0.944444444444 -1.0303030303 0 -0.8 1e-06 
1.0 -1.0303030303 0 -0.8 1e-06 
0.5 -0.989898989899 0 -0.8 1e-06 
0.555555555556 -0.989898989899 0 -0.8 1e-06 
0.611111111111 -0.989898989899 0 -0.8 1e-06 
0.666666666667 -0.989898989899 0 -0.8 1e-06 
0.722222222222 -0.989898989899 0 -0.8 1e-06 
0.777777777778 -0.989898989899 0 -0.8 1e-06 
0.833333333333 -0.989898989899 0 -0.8 1e-06 
0.888888888889 -0.989898989899 0 -0.8 1e-06 
0.944444444444 -0.989898989899 0 -0.8 1e-06 
1.0 -0.989898989899 0 -0.8 1e-06 
0.5 -0.949494949495 0 -0.8 1e-06 
0.555555555556 -0.949494949495 0 -0.8 1e-06 
0.611111111111 -0.949494949495 0 -0.8 1e-06 
0.666666666667 -0.949494949495 0 -0.8 1e-06 
0.722222222222 -0.949494949495 0 -0.8 1e-06 
0.777777777778 -0.949494949495 0 -0.8 1e-06 
0.833333333333 -0.949494949495 0 -0.8 1e-06 
0.888888888889 -0.949494949495 0 -0.8 1e-06 
0.944444444444 -0.949494949495 0 -0.8 1e-06 
1.0 -0.949494949495 0 -0.8 1e-06 
0.5 -0.909090909091 0 -0.8 1e-06 
0.555555555556 -0.909090909091 0 -0.8 1e-06 
0.611111111111 -0.909090909091 0 -0.8 1e-06 
0.666666666667 -0.909090909091 0 -0.8 1e-06 
0.722222222222 -0.909090909091 0 -0.8 1e-06 
0.777777777778 -0.909090909091 0 -0.8 1e-06 
0.833333333333 -0.909090909091 0 -0.8 1e-06 
0.888888888889 -0.909090909091 0 -0.8 1e-06 
0.944444444444 -0.909090909091 0 -0.8 1e-06 
1.0 -0.909090909091 0 -0.8 1e-06 
0.5 -0.868686868687 0 -0.8 1e-06 
0.555555555556 -0.868686868687 0 -0.8 1e-06 
0.611111111111 -0.868686868687 0 -0.8 1e-06 
0.666666666667 -0.868686868687 0 -0.8 1e-06 
0.722222222222 -0.868686868687 0 -0.8 1e-06 
0.777777777778 -0.868686868687 0 -0.8 1e-06 
0.833333333333 -0.868686868687 0 -0.8 1e-06 
0.888888888889 -0.868686868687 0 -0.8 1e-06 
0.944444444444 -0.868686868687 0 -0.8 1e-06 
1.0 -0.868686868687 0 -0.8 1e-06 
0.5 -0.828282828283 0 -0.8 1e-06 
0.555555555556 -0.828282828283 0 -0.8 1e-06 
0.611111111111 -0.828282828283 0 -0.8 1e-06 
0.666666666667 -0.828282828283 0 -0.8 1e-06 
0.722222222222 -0.828282828283 0 -0.8 1e-06 
0.777777777778 -0.828282828283 0 -0.8 1e-06 
0.833333333333 -0.828282828283 0 -0.8 1e-06 
0.888888888889 -0.828282828283 0 -0.8 1e-06 
0.944444444444 -0.828282828283 0 -0.8 1e-06 
1.0 -0.828282828283 0 -0.8 1e-06 
0.5 -0.787878787879 0 -0.8 1e-06 
0.555555555556 -0.787878787879 0 -0.8 1e-06 
0.611111111111 -0.787878787879 0 -0.8 1e-06 
0.666666666667 -0.787878787879 0 -0.8 1e-06 
0.722222222222 -0.787878787879 0 -0.8 1e-06 
0.777777777778 -0.787878787879 0 -0.8 1e-06 
0.833333333333 -0.787878787879 0 -0.8 1e-06 
0.888888888889 -0.787878787879 0 -0.8 1e-06 
0.944444444444 -0.787878787879 0 -0.8 1e-06 
1.0 -0.787878787879 0 -0.8 1e-06 
0.5 -0.747474747475 0 -0.8 1e-06 
0.555555555556 -0.747474747475 0 -0.8 1e-06 
0.611111111111 -0.747474747475 0 -0.8 1e-06 
0.666666666667 -0.747474747475 0 -0.8 1e-06 
0.722222222222 -0.747474747475 0 -0.8 1e-06 
0.777777777778 -0.747474747475 0 -0.8 1e-06 
0.833333333333 -0.747474747475 0 -0.8 1e-06 
0.888888888889 -0.747474747475 0 -0.8 1e-06 
0.944444444444 -0.747474747475 0 -0.8 1e-06 
1.0 -0.747474747475 0 -0.8 1e-06 
0.5 -0.707070707071 0 -0.8 1e-06 
0.555555555556 -0.707070707071 0 -0.8 1e-06 
0.611111111111 -0.707070707071 0 -0.8 1e-06 
0.666666666667 -0.707070707071 0 -0.8 1e-06 
0.722222222222 -0.707070707071 0 -0.8 1e-06 
0.777777777778 -0.707070707071 0 -0.8 1e-06 
0.833333333333 -0.707070707071 0 -0.8 1e-06 
0.888888888889 -0.707070707071 0 -0.8 1e-06 
0.944444444444 -0.707070707071 0 -0.8 1e-06 
1.0 -0.707070707071 0 -0.8 1e-06 
0.5 -0.666666666667 0 -0.8 1e-06 
0.555555555556 -0.666666666667 0 -0.8 1e-06 
0.611111111111 -0.666666666667 0 -0.8 1e-06 
0.666666666667 -0.666666666667 0 -0.8 1e-06 
0.722222222222 -0.666666666667 0 -0.8 1e-06 
0.777777777778 -0.666666666667 0 -0.8 1e-06 
0.833333333333 -0.666666666667 0 -0.8 1e-06 
0.888888888889 -0.666666666667 0 -0.8 1e-06 
0.944444444444 -0.666666666667 0 -0.8 1e-06 
1.0 -0.666666666667 0 -0.8 1e-06 
0.5 -0.626262626263 0 -0.8 1e-06 
0.555555555556 -0.626262626263 0 -0.8 1e-06 
0.611111111111 -0.626262626263 0 -0.8 1e-06 
0.666666666667 -0.626262626263 0 -0.8 1e-06 
0.722222222222 -0.626262626263 0 -0.8 1e-06 
0.777777777778 -0.626262626263 0 -0.8 1e-06 
0.833333333333 -0.626262626263 0 -0.8 1e-06 
0.888888888889 -0.626262626263 0 -0.8 1e-06 
0.944444444444 -0.626262626263 0 -0.8 1e-06 
1.0 -0.626262626263 0 -0.8 1e-06 
0.5 -0.585858585859 0 -0.8 1e-06 
0.555555555556 -0.585858585859 0 -0.8 1e-06 
0.611111111111 -0.585858585859 0 -0.8 1e-06 
0.666666666667 -0.585858585859 0 -0.8 1e-06 
0.722222222222 -0.585858585859 0 -0.8 1e-06 
0.777777777778 -0.585858585859 0 -0.8 1e-06 
0.833333333333 -0.585858585859 0 -0.8 1e-06 
0.888888888889 -0.585858585859 0 -0.8 1e-06 
0.944444444444 -0.585858585859 0 -0.8 1e-06 
1.0 -0.585858585859 0 -0.8 1e-06 
0.5 -0.545454545455 0 -0.8 1e-06 
0.555555555556 -0.545454545455 0 -0.8 1e-06 
0.611111111111 -0.545454545455 0 -0.8 1e-06 
0.666666666667 -0.545454545455 0 -0.8 1e-06 
0.722222222222 -0.545454545455 0 -0.8 1e-06 
0.777777777778 -0.545454545455 0 -0.8 1e-06 
0.833333333333 -0.545454545455 0 -0.8 1e-06 
0.888888888889 -0.545454545455 0 -0.8 1e-06 
0.944444444444 -0.545454545455 0 -0.8 1e-06 
1.0 -0.545454545455 0 -0.8 1e-06 
0.5 -0.505050505051 0 -0.8 1e-06 
0.555555555556 -0.505050505051 0 -0.8 1e-06 
0.611111111111 -0.505050505051 0 -0.8 1e-06 
0.666666666667 -0.505050505051 0 -0.8 1e-06 
0.722222222222 -0.505050505051 0 -0.8 1e-06 
0.777777777778 -0.505050505051 0 -0.8 1e-06 
0.833333333333 -0.505050505051 0 -0.8 1e-06 
0.888888888889 -0.505050505051 0 -0.8 1e-06 
0.944444444444 -0.505050505051 0 -0.8 1e-06 
1.0 -0.505050505051 0 -0.8 1e-06 
0.5 -0.464646464646 0 -0.8 1e-06 
0.555555555556 -0.464646464646 0 -0.8 1e-06 
0.611111111111 -0.464646464646 0 -0.8 1e-06 
0.666666666667 -0.464646464646 0 -0.8 1e-06 
0.722222222222 -0.464646464646 0 -0.8 1e-06 
0.777777777778 -0.464646464646 0 -0.8 1e-06 
0.833333333333 -0.464646464646 0 -0.8 1e-06 
0.888888888889 -0.464646464646 0 -0.8 1e-06 
0.944444444444 -0.464646464646 0 -0.8 1e-06 
1.0 -0.464646464646 0 -0.8 1e-06 
0.5 -0.424242424242 0 -0.8 1e-06 
0.555555555556 -0.424242424242 0 -0.8 1e-06 
0.611111111111 -0.424242424242 0 -0.8 1e-06 
0.666666666667 -0.424242424242 0 -0.8 1e-06 
0.722222222222 -0.424242424242 0 -0.8 1e-06 
0.777777777778 -0.424242424242 0 -0.8 1e-06 
0.833333333333 -0.424242424242 0 -0.8 1e-06 
0.888888888889 -0.424242424242 0 -0.8 1e-06 
0.944444444444 -0.424242424242 0 -0.8 1e-06 
1.0 -0.424242424242 0 -0.8 1e-06 
0.5 -0.383838383838 0 -0.8 1e-06 
0.555555555556 -0.383838383838 0 -0.8 1e-06 
0.611111111111 -0.383838383838 0 -0.8 1e-06 
0.666666666667 -0.383838383838 0 -0.8 1e-06 
0.722222222222 -0.383838383838 0 -0.8 1e-06 
0.777777777778 -0.383838383838 0 -0.8 1e-06 
0.833333333333 -0.383838383838 0 -0.8 1e-06 
0.888888888889 -0.383838383838 0 -0.8 1e-06 
0.944444444444 -0.383838383838 0 -0.8 1e-06 
1.0 -0.383838383838 0 -0.8 1e-06 
0.5 -0.343434343434 0 -0.8 1e-06 
0.555555555556 -0.343434343434 0 -0.8 1e-06 
0.611111111111 -0.343434343434 0 -0.8 1e-06 
0.666666666667 -0.343434343434 0 -0.8 1e-06 
0.722222222222 -0.343434343434 0 -0.8 1e-06 
0.777777777778 -0.343434343434 0 -0.8 1e-06 
0.833333333333 -0.343434343434 0 -0.8 1e-06 
0.888888888889 -0.343434343434 0 -0.8 1e-06 
0.944444444444 -0.343434343434 0 -0.8 1e-06 
1.0 -0.343434343434 0 -0.8 1e-06 
0.5 -0.30303030303 0 -0.8 1e-06 
0.555555555556 -0.30303030303 0 -0.8 1e-06 
0.611111111111 -0.30303030303 0 -0.8 1e-06 
0.666666666667 -0.30303030303 0 -0.8 1e-06 
0.722222222222 -0.30303030303 0 -0.8 1e-06 
0.777777777778 -0.30303030303 0 -0.8 1e-06 
0.833333333333 -0.30303030303 0 -0.8 1e-06 
0.888888888889 -0.30303030303 0 -0.8 1e-06 
0.944444444444 -0.30303030303 0 -0.8 1e-06 
1.0 -0.30303030303 0 -0.8 1e-06 
0.5 -0.262626262626 0 -0.8 1e-06 
0.555555555556 -0.262626262626 0 -0.8 1e-06 
0.611111111111 -0.262626262626 0 -0.8 1e-06 
0.666666666667 -0.262626262626 0 -0.8 1e-06 
0.722222222222 -0.262626262626 0 -0.8 1e-06 
0.777777777778 -0.262626262626 0 -0.8 1e-06 
0.833333333333 -0.262626262626 0 -0.8 1e-06 
0.888888888889 -0.262626262626 0 -0.8 1e-06 
0.944444444444 -0.262626262626 0 -0.8 1e-06 
1.0 -0.262626262626 0 -0.8 1e-06 
0.5 -0.222222222222 0 -0.8 1e-06 
0.555555555556 -0.222222222222 0 -0.8 1e-06 
0.611111111111 -0.222222222222 0 -0.8 1e-06 
0.666666666667 -0.222222222222 0 -0.8 1e-06 
0.722222222222 -0.222222222222 0 -0.8 1e-06 
0.777777777778 -0.222222222222 0 -0.8 1e-06 
0.833333333333 -0.222222222222 0 -0.8 1e-06 
0.888888888889 -0.222222222222 0 -0.8 1e-06 
0.944444444444 -0.222222222222 0 -0.8 1e-06 
1.0 -0.222222222222 0 -0.8 1e-06 
0.5 -0.181818181818 0 -0.8 1e-06 
0.555555555556 -0.181818181818 0 -0.8 1e-06 
0.611111111111 -0.181818181818 0 -0.8 1e-06 
0.666666666667 -0.181818181818 0 -0.8 1e-06 
0.722222222222 -0.181818181818 0 -0.8 1e-06 
0.777777777778 -0.181818181818 0 -0.8 1e-06 
0.833333333333 -0.181818181818 0 -0.8 1e-06 
0.888888888889 -0.181818181818 0 -0.8 1e-06 
0.944444444444 -0.181818181818 0 -0.8 1e-06 
1.0 -0.181818181818 0 -0.8 1e-06 
0.5 -0.141414141414 0 -0.8 1e-06 
0.555555555556 -0.141414141414 0 -0.8 1e-06 
0.611111111111 -0.141414141414 0 -0.8 1e-06 
0.666666666667 -0.141414141414 0 -0.8 1e-06 
0.722222222222 -0.141414141414 0 -0.8 1e-06 
0.777777777778 -0.141414141414 0 -0.8 1e-06 
0.833333333333 -0.141414141414 0 -0.8 1e-06 
0.888888888889 -0.141414141414 0 -0.8 1e-06 
0.944444444444 -0.141414141414 0 -0.8 1e-06 
1.0 -0.141414141414 0 -0.8 1e-06 
0.5 -0.10101010101 0 -0.8 1e-06 
0.555555555556 -0.10101010101 0 -0.8 1e-06 
0.611111111111 -0.10101010101 0 -0.8 1e-06 
0.666666666667 -0.10101010101 0 -0.8 1e-06 
0.722222222222 -0.10101010101 0 -0.8 1e-06 
0.777777777778 -0.10101010101 0 -0.8 1e-06 
0.833333333333 -0.10101010101 0 -0.8 1e-06 
0.888888888889 -0.10101010101 0 -0.8 1e-06 
0.944444444444 -0.10101010101 0 -0.8 1e-06 
1.0 -0.10101010101 0 -0.8 1e-06 
0.5 -0.0606060606061 0 -0.8 1e-06 
0.555555555556 -0.0606060606061 0 -0.8 1e-06 
0.611111111111 -0.0606060606061 0 -0.8 1e-06 
0.666666666667 -0.0606060606061 0 -0.8 1e-06 
0.722222222222 -0.0606060606061 0 -0.8 1e-06 
0.777777777778 -0.0606060606061 0 -0.8 1e-06 
0.833333333333 -0.0606060606061 0 -0.8 1e-06 
0.888888888889 -0.0606060606061 0 -0.8 1e-06 
0.944444444444 -0.0606060606061 0 -0.8 1e-06 
1.0 -0.0606060606061 0 -0.8 1e-06 
0.5 -0.020202020202 0 -0.8 1e-06 
0.555555555556 -0.020202020202 0 -0.8 1e-06 
0.611111111111 -0.020202020202 0 -0.8 1e-06 
0.666666666667 -0.020202020202 0 -0.8 1e-06 
0.722222222222 -0.020202020202 0 -0.8 1e-06 
0.777777777778 -0.020202020202 0 -0.8 1e-06 
0.833333333333 -0.020202020202 0 -0.8 1e-06 
0.888888888889 -0.020202020202 0 -0.8 1e-06 
0.944444444444 -0.020202020202 0 -0.8 1e-06 
1.0 -0.020202020202 0 -0.8 1e-06 
0.5 0.020202020202 0 -0.8 1e-06 
0.555555555556 0.020202020202 0 -0.8 1e-06 
0.611111111111 0.020202020202 0 -0.8 1e-06 
0.666666666667 0.020202020202 0 -0.8 1e-06 
0.722222222222 0.020202020202 0 -0.8 1e-06 
0.777777777778 0.020202020202 0 -0.8 1e-06 
0.833333333333 0.020202020202 0 -0.8 1e-06 
0.888888888889 0.020202020202 0 -0.8 1e-06 
0.944444444444 0.020202020202 0 -0.8 1e-06 
1.0 0.020202020202 0 -0.8 1e-06 
0.5 0.0606060606061 0 -0.8 1e-06 
0.555555555556 0.0606060606061 0 -0.8 1e-06 
0.611111111111 0.0606060606061 0 -0.8 1e-06 
0.666666666667 0.0606060606061 0 -0.8 1e-06 
0.722222222222 0.0606060606061 0 -0.8 1e-06 
0.777777777778 0.0606060606061 0 -0.8 1e-06 
0.833333333333 0.0606060606061 0 -0.8 1e-06 
0.888888888889 0.0606060606061 0 -0.8 1e-06 
0.944444444444 0.0606060606061 0 -0.8 1e-06 
1.0 0.0606060606061 0 -0.8 1e-06 
0.5 0.10101010101 0 -0.8 1e-06 
0.555555555556 0.10101010101 0 -0.8 1e-06 
0.611111111111 0.10101010101 0 -0.8 1e-06 
0.666666666667 0.10101010101 0 -0.8 1e-06 
0.722222222222 0.10101010101 0 -0.8 1e-06 
0.777777777778 0.10101010101 0 -0.8 1e-06 
0.833333333333 0.10101010101 0 -0.8 1e-06 
0.888888888889 0.10101010101 0 -0.8 1e-06 
0.944444444444 0.10101010101 0 -0.8 1e-06 
1.0 0.10101010101 0 -0.8 1e-06 
0.5 0.141414141414 0 -0.8 1e-06 
0.555555555556 0.141414141414 0 -0.8 1e-06 
0.611111111111 0.141414141414 0 -0.8 1e-06 
0.666666666667 0.141414141414 0 -0.8 1e-06 
0.722222222222 0.141414141414 0 -0.8 1e-06 
0.777777777778 0.141414141414 0 -0.8 1e-06 
0.833333333333 0.141414141414 0 -0.8 1e-06 
0.888888888889 0.141414141414 0 -0.8 1e-06 
0.944444444444 0.141414141414 0 -0.8 1e-06 
1.0 0.141414141414 0 -0.8 1e-06 
0.5 0.181818181818 0 -0.8 1e-06 
0.555555555556 0.181818181818 0 -0.8 1e-06 
0.611111111111 0.181818181818 0 -0.8 1e-06 
0.666666666667 0.181818181818 0 -0.8 1e-06 
0.722222222222 0.181818181818 0 -0.8 1e-06 
0.777777777778 0.181818181818 0 -0.8 1e-06 
0.833333333333 0.181818181818 0 -0.8 1e-06 
0.888888888889 0.181818181818 0 -0.8 1e-06 
0.944444444444 0.181818181818 0 -0.8 1e-06 
1.0 0.181818181818 0 -0.8 1e-06 
0.5 0.222222222222 0 -0.8 1e-06 
0.555555555556 0.222222222222 0 -0.8 1e-06 
0.611111111111 0.222222222222 0 -0.8 1e-06 
0.666666666667 0.222222222222 0 -0.8 1e-06 
0.722222222222 0.222222222222 0 -0.8 1e-06 
0.777777777778 0.222222222222 0 -0.8 1e-06 
0.833333333333 0.222222222222 0 -0.8 1e-06 
0.888888888889 0.222222222222 0 -0.8 1e-06 
0.944444444444 0.222222222222 0 -0.8 1e-06 
1.0 0.222222222222 0 -0.8 1e-06 
0.5 0.262626262626 0 -0.8 1e-06 
0.555555555556 0.262626262626 0 -0.8 1e-06 
0.611111111111 0.262626262626 0 -0.8 1e-06 
0.666666666667 0.262626262626 0 -0.8 1e-06 
0.722222222222 0.262626262626 0 -0.8 1e-06 
0.777777777778 0.262626262626 0 -0.8 1e-06 
0.833333333333 0.262626262626 0 -0.8 1e-06 
0.888888888889 0.262626262626 0 -0.8 1e-06 
0.944444444444 0.262626262626 0 -0.8 1e-06 
1.0 0.262626262626 0 -0.8 1e-06 
0.5 0.30303030303 0 -0.8 1e-06 
0.555555555556 0.30303030303 0 -0.8 1e-06 
0.611111111111 0.30303030303 0 -0.8 1e-06 
0.666666666667 0.30303030303 0 -0.8 1e-06 
0.722222222222 0.30303030303 0 -0.8 1e-06 
0.777777777778 0.30303030303 0 -0.8 1e-06 
0.833333333333 0.30303030303 0 -0.8 1e-06 
0.888888888889 0.30303030303 0 -0.8 1e-06 
0.944444444444 0.30303030303 0 -0.8 1e-06 
1.0 0.30303030303 0 -0.8 1e-06 
0.5 0.343434343434 0 -0.8 1e-06 
0.555555555556 0.343434343434 0 -0.8 1e-06 
0.611111111111 0.343434343434 0 -0.8 1e-06 
0.666666666667 0.343434343434 0 -0.8 1e-06 
0.722222222222 0.343434343434 0 -0.8 1e-06 
0.777777777778 0.343434343434 0 -0.8 1e-06 
0.833333333333 0.343434343434 0 -0.8 1e-06 
0.888888888889 0.343434343434 0 -0.8 1e-06 
0.944444444444 0.343434343434 0 -0.8 1e-06 
1.0 0.343434343434 0 -0.8 1e-06 
0.5 0.383838383838 0 -0.8 1e-06 
0.555555555556 0.383838383838 0 -0.8 1e-06 
0.611111111111 0.383838383838 0 -0.8 1e-06 
0.666666666667 0.383838383838 0 -0.8 1e-06 
0.722222222222 0.383838383838 0 -0.8 1e-06 
0.777777777778 0.383838383838 0 -0.8 1e-06 
0.833333333333 0.383838383838 0 -0.8 1e-06 
0.888888888889 0.383838383838 0 -0.8 1e-06 
0.944444444444 0.383838383838 0 -0.8 1e-06 
1.0 0.383838383838 0 -0.8 1e-06 
0.5 0.424242424242 0 -0.8 1e-06 
0.555555555556 0.424242424242 0 -0.8 1e-06 
0.611111111111 0.424242424242 0 -0.8 1e-06 
0.666666666667 0.424242424242 0 -0.8 1e-06 
0.722222222222 0.424242424242 0 -0.8 1e-06 
0.777777777778 0.424242424242 0 -0.8 1e-06 
0.833333333333 0.424242424242 0 -0.8 1e-06 
0.888888888889 0.424242424242 0 -0.8 1e-06 
0.944444444444 0.424242424242 0 -0.8 1e-06 
1.0 0.424242424242 0 -0.8 1e-06 
0.5 0.464646464646 0 -0.8 1e-06 
0.555555555556 0.464646464646 0 -0.8 1e-06 
0.611111111111 0.464646464646 0 -0.8 1e-06 
0.666666666667 0.464646464646 0 -0.8 1e-06 
0.722222222222 0.464646464646 0 -0.8 1e-06 
0.777777777778 0.464646464646 0 -0.8 1e-06 
0.833333333333 0.464646464646 0 -0.8 1e-06 
0.888888888889 0.464646464646 0 -0.8 1e-06 
0.944444444444 0.464646464646 0 -0.8 1e-06 
1.0 0.464646464646 0 -0.8 1e-06 
0.5 0.505050505051 0 -0.8 1e-06 
0.555555555556 0.505050505051 0 -0.8 1e-06 
0.611111111111 0.505050505051 0 -0.8 1e-06 
0.666666666667 0.505050505051 0 -0.8 1e-06 
0.722222222222 0.505050505051 0 -0.8 1e-06 
0.777777777778 0.505050505051 0 -0.8 1e-06 
0.833333333333 0.505050505051 0 -0.8 1e-06 
0.888888888889 0.505050505051 0 -0.8 1e-06 
0.944444444444 0.505050505051 0 -0.8 1e-06 
1.0 0.505050505051 0 -0.8 1e-06 
0.5 0.545454545455 0 -0.8 1e-06 
0.555555555556 0.545454545455 0 -0.8 1e-06 
0.611111111111 0.545454545455 0 -0.8 1e-06 
0.666666666667 0.545454545455 0 -0.8 1e-06 
0.722222222222 0.545454545455 0 -0.8 1e-06 
0.777777777778 0.545454545455 0 -0.8 1e-06 
0.833333333333 0.545454545455 0 -0.8 1e-06 
0.888888888889 0.545454545455 0 -0.8 1e-06 
0.944444444444 0.545454545455 0 -0.8 1e-06 
1.0 0.545454545455 0 -0.8 1e-06 
0.5 0.585858585859 0 -0.8 1e-06 
0.555555555556 0.585858585859 0 -0.8 1e-06 
0.611111111111 0.585858585859 0 -0.8 1e-06 
0.666666666667 0.585858585859 0 -0.8 1e-06 
0.722222222222 0.585858585859 0 -0.8 1e-06 
0.777777777778 0.585858585859 0 -0.8 1e-06 
0.833333333333 0.585858585859 0 -0.8 1e-06 
0.888888888889 0.585858585859 0 -0.8 1e-06 
0.944444444444 0.585858585859 0 -0.8 1e-06 
1.0 0.585858585859 0 -0.8 1e-06 
0.5 0.626262626263 0 -0.8 1e-06 
0.555555555556 0.626262626263 0 -0.8 1e-06 
0.611111111111 0.626262626263 0 -0.8 1e-06 
0.666666666667 0.626262626263 0 -0.8 1e-06 
0.722222222222 0.626262626263 0 -0.8 1e-06 
0.777777777778 0.626262626263 0 -0.8 1e-06 
0.833333333333 0.626262626263 0 -0.8 1e-06 
0.888888888889 0.626262626263 0 -0.8 1e-06 
0.944444444444 0.626262626263 0 -0.8 1e-06 
1.0 0.626262626263 0 -0.8 1e-06 
0.5 0.666666666667 0 -0.8 1e-06 
0.555555555556 0.666666666667 0 -0.8 1e-06 
0.611111111111 0.666666666667 0 -0.8 1e-06 
0.666666666667 0.666666666667 0 -0.8 1e-06 
0.722222222222 0.666666666667 0 -0.8 1e-06 
0.777777777778 0.666666666667 0 -0.8 1e-06 
0.833333333333 0.666666666667 0 -0.8 1e-06 
0.888888888889 0.666666666667 0 -0.8 1e-06 
0.944444444444 0.666666666667 0 -0.8 1e-06 
1.0 0.666666666667 0 -0.8 1e-06 
0.5 0.707070707071 0 -0.8 1e-06 
0.555555555556 0.707070707071 0 -0.8 1e-06 
0.611111111111 0.707070707071 0 -0.8 1e-06 
0.666666666667 0.707070707071 0 -0.8 1e-06 
0.722222222222 0.707070707071 0 -0.8 1e-06 
0.777777777778 0.707070707071 0 -0.8 1e-06 
0.833333333333 0.707070707071 0 -0.8 1e-06 
0.888888888889 0.707070707071 0 -0.8 1e-06 
0.944444444444 0.707070707071 0 -0.8 1e-06 
1.0 0.707070707071 0 -0.8 1e-06 
0.5 0.747474747475 0 -0.8 1e-06 
0.555555555556 0.747474747475 0 -0.8 1e-06 
0.611111111111 0.747474747475 0 -0.8 1e-06 
0.666666666667 0.747474747475 0 -0.8 1e-06 
0.722222222222 0.747474747475 0 -0.8 1e-06 
0.777777777778 0.747474747475 0 -0.8 1e-06 
0.833333333333 0.747474747475 0 -0.8 1e-06 
0.888888888889 0.747474747475 0 -0.8 1e-06 
0.944444444444 0.747474747475 0 -0.8 1e-06 
1.0 0.747474747475 0 -0.8 1e-06 
0.5 0.787878787879 0 -0.8 1e-06 
0.555555555556 0.787878787879 0 -0.8 1e-06 
0.611111111111 0.787878787879 0 -0.8 1e-06 
0.666666666667 0.787878787879 0 -0.8 1e-06 
0.722222222222 0.787878787879 0 -0.8 1e-06 
0.777777777778 0.787878787879 0 -0.8 1e-06 
0.833333333333 0.787878787879 0 -0.8 1e-06 
0.888888888889 0.787878787879 0 -0.8 1e-06 
0.944444444444 0.787878787879 0 -0.8 1e-06 
1.0 0.787878787879 0 -0.8 1e-06 
0.5 0.828282828283 0 -0.8 1e-06 
0.555555555556 0.828282828283 0 -0.8 1e-06 
0.611111111111 0.828282828283 0 -0.8 1e-06 
0.666666666667 0.828282828283 0 -0.8 1e-06 
0.722222222222 0.828282828283 0 -0.8 1e-06 
0.777777777778 0.828282828283 0 -0.8 1e-06 
0.833333333333 0.828282828283 0 -0.8 1e-06 
0.888888888889 0.828282828283 0 -0.8 1e-06 
0.944444444444 0.828282828283 0 -0.8 1e-06 
1.0 0.828282828283 0 -0.8 1e-06 
0.5 0.868686868687 0 -0.8 1e-06 
0.555555555556 0.868686868687 0 -0.8 1e-06 
0.611111111111 0.868686868687 0 -0.8 1e-06 
0.666666666667 0.868686868687 0 -0.8 1e-06 
0.722222222222 0.868686868687 0 -0.8 1e-06 
0.777777777778 0.868686868687 0 -0.8 1e-06 
0.833333333333 0.868686868687 0 -0.8 1e-06 
0.888888888889 0.868686868687 0 -0.8 1e-06 
0.944444444444 0.868686868687 0 -0.8 1e-06 
1.0 0.868686868687 0 -0.8 1e-06 
0.5 0.909090909091 0 -0.8 1e-06 
0.555555555556 0.909090909091 0 -0.8 1e-06 
0.611111111111 0.909090909091 0 -0.8 1e-06 
0.666666666667 0.909090909091 0 -0.8 1e-06 
0.722222222222 0.909090909091 0 -0.8 1e-06 
0.777777777778 0.909090909091 0 -0.8 1e-06 
0.833333333333 0.909090909091 0 -0.8 1e-06 
0.888888888889 0.909090909091 0 -0.8 1e-06 
0.944444444444 0.909090909091 0 -0.8 1e-06 
1.0 0.909090909091 0 -0.8 1e-06 
0.5 0.949494949495 0 -0.8 1e-06 
0.555555555556 0.949494949495 0 -0.8 1e-06 
0.611111111111 0.949494949495 0 -0.8 1e-06 
0.666666666667 0.949494949495 0 -0.8 1e-06 
0.722222222222 0.949494949495 0 -0.8 1e-06 
0.777777777778 0.949494949495 0 -0.8 1e-06 
0.833333333333 0.949494949495 0 -0.8 1e-06 
0.888888888889 0.949494949495 0 -0.8 1e-06 
0.944444444444 0.949494949495 0 -0.8 1e-06 
1.0 0.949494949495 0 -0.8 1e-06 
0.5 0.989898989899 0 -0.8 1e-06 
0.555555555556 0.989898989899 0 -0.8 1e-06 
0.611111111111 0.989898989899 0 -0.8 1e-06 
0.666666666667 0.989898989899 0 -0.8 1e-06 
0.722222222222 0.989898989899 0 -0.8 1e-06 
0.777777777778 0.989898989899 0 -0.8 1e-06 
0.833333333333 0.989898989899 0 -0.8 1e-06 
0.888888888889 0.989898989899 0 -0.8 1e-06 
0.944444444444 0.989898989899 0 -0.8 1e-06 
1.0 0.989898989899 0 -0.8 1e-06 
0.5 1.0303030303 0 -0.8 1e-06 
0.555555555556 1.0303030303 0 -0.8 1e-06 
0.611111111111 1.0303030303 0 -0.8 1e-06 
0.666666666667 1.0303030303 0 -0.8 1e-06 
0.722222222222 1.0303030303 0 -0.8 1e-06 
0.777777777778 1.0303030303 0 -0.8 1e-06 
0.833333333333 1.0303030303 0 -0.8 1e-06 
0.888888888889 1.0303030303 0 -0.8 1e-06 
0.944444444444 1.0303030303 0 -0.8 1e-06 
1.0 1.0303030303 0 -0.8 1e-06 
0.5 1.07070707071 0 -0.8 1e-06 
0.555555555556 1.07070707071 0 -0.8 1e-06 
0.611111111111 1.07070707071 0 -0.8 1e-06 
0.666666666667 1.07070707071 0 -0.8 1e-06 
0.722222222222 1.07070707071 0 -0.8 1e-06 
0.777777777778 1.07070707071 0 -0.8 1e-06 
0.833333333333 1.07070707071 0 -0.8 1e-06 
0.888888888889 1.07070707071 0 -0.8 1e-06 
0.944444444444 1.07070707071 0 -0.8 1e-06 
1.0 1.07070707071 0 -0.8 1e-06 
0.5 1.11111111111 0 -0.8 1e-06 
0.555555555556 1.11111111111 0 -0.8 1e-06 
0.611111111111 1.11111111111 0 -0.8 1e-06 
0.666666666667 1.11111111111 0 -0.8 1e-06 
0.722222222222 1.11111111111 0 -0.8 1e-06 
0.777777777778 1.11111111111 0 -0.8 1e-06 
0.833333333333 1.11111111111 0 -0.8 1e-06 
0.888888888889 1.11111111111 0 -0.8 1e-06 
0.944444444444 1.11111111111 0 -0.8 1e-06 
1.0 1.11111111111 0 -0.8 1e-06 
0.5 1.15151515152 0 -0.8 1e-06 
0.555555555556 1.15151515152 0 -0.8 1e-06 
0.611111111111 1.15151515152 0 -0.8 1e-06 
0.666666666667 1.15151515152 0 -0.8 1e-06 
0.722222222222 1.15151515152 0 -0.8 1e-06 
0.777777777778 1.15151515152 0 -0.8 1e-06 
0.833333333333 1.15151515152 0 -0.8 1e-06 
0.888888888889 1.15151515152 0 -0.8 1e-06 
0.944444444444 1.15151515152 0 -0.8 1e-06 
1.0 1.15151515152 0 -0.8 1e-06 
0.5 1.19191919192 0 -0.8 1e-06 
0.555555555556 1.19191919192 0 -0.8 1e-06 
0.611111111111 1.19191919192 0 -0.8 1e-06 
0.666666666667 1.19191919192 0 -0.8 1e-06 
0.722222222222 1.19191919192 0 -0.8 1e-06 
0.777777777778 1.19191919192 0 -0.8 1e-06 
0.833333333333 1.19191919192 0 -0.8 1e-06 
0.888888888889 1.19191919192 0 -0.8 1e-06 
0.944444444444 1.19191919192 0 -0.8 1e-06 
1.0 1.19191919192 0 -0.8 1e-06 
0.5 1.23232323232 0 -0.8 1e-06 
0.555555555556 1.23232323232 0 -0.8 1e-06 
0.611111111111 1.23232323232 0 -0.8 1e-06 
0.666666666667 1.23232323232 0 -0.8 1e-06 
0.722222222222 1.23232323232 0 -0.8 1e-06 
0.777777777778 1.23232323232 0 -0.8 1e-06 
0.833333333333 1.23232323232 0 -0.8 1e-06 
0.888888888889 1.23232323232 0 -0.8 1e-06 
0.944444444444 1.23232323232 0 -0.8 1e-06 
1.0 1.23232323232 0 -0.8 1e-06 
0.5 1.27272727273 0 -0.8 1e-06 
0.555555555556 1.27272727273 0 -0.8 1e-06 
0.611111111111 1.27272727273 0 -0.8 1e-06 
0.666666666667 1.27272727273 0 -0.8 1e-06 
0.722222222222 1.27272727273 0 -0.8 1e-06 
0.777777777778 1.27272727273 0 -0.8 1e-06 
0.833333333333 1.27272727273 0 -0.8 1e-06 
0.888888888889 1.27272727273 0 -0.8 1e-06 
0.944444444444 1.27272727273 0 -0.8 1e-06 
1.0 1.27272727273 0 -0.8 1e-06 
0.5 1.31313131313 0 -0.8 1e-06 
0.555555555556 1.31313131313 0 -0.8 1e-06 
0.611111111111 1.31313131313 0 -0.8 1e-06 
0.666666666667 1.31313131313 0 -0.8 1e-06 
0.722222222222 1.31313131313 0 -0.8 1e-06 
0.777777777778 1.31313131313 0 -0.8 1e-06 
0.833333333333 1.31313131313 0 -0.8 1e-06 
0.888888888889 1.31313131313 0 -0.8 1e-06 
0.944444444444 1.31313131313 0 -0.8 1e-06 
1.0 1.31313131313 0 -0.8 1e-06 
0.5 1.35353535354 0 -0.8 1e-06 
0.555555555556 1.35353535354 0 -0.8 1e-06 
0.611111111111 1.35353535354 0 -0.8 1e-06 
0.666666666667 1.35353535354 0 -0.8 1e-06 
0.722222222222 1.35353535354 0 -0.8 1e-06 
0.777777777778 1.35353535354 0 -0.8 1e-06 
0.833333333333 1.35353535354 0 -0.8 1e-06 
0.888888888889 1.35353535354 0 -0.8 1e-06 
0.944444444444 1.35353535354 0 -0.8 1e-06 
1.0 1.35353535354 0 -0.8 1e-06 
0.5 1.39393939394 0 -0.8 1e-06 
0.555555555556 1.39393939394 0 -0.8 1e-06 
0.611111111111 1.39393939394 0 -0.8 1e-06 
0.666666666667 1.39393939394 0 -0.8 1e-06 
0.722222222222 1.39393939394 0 -0.8 1e-06 
0.777777777778 1.39393939394 0 -0.8 1e-06 
0.833333333333 1.39393939394 0 -0.8 1e-06 
0.888888888889 1.39393939394 0 -0.8 1e-06 
0.944444444444 1.39393939394 0 -0.8 1e-06 
1.0 1.39393939394 0 -0.8 1e-06 
0.5 1.43434343434 0 -0.8 1e-06 
0.555555555556 1.43434343434 0 -0.8 1e-06 
0.611111111111 1.43434343434 0 -0.8 1e-06 
0.666666666667 1.43434343434 0 -0.8 1e-06 
0.722222222222 1.43434343434 0 -0.8 1e-06 
0.777777777778 1.43434343434 0 -0.8 1e-06 
0.833333333333 1.43434343434 0 -0.8 1e-06 
0.888888888889 1.43434343434 0 -0.8 1e-06 
0.944444444444 1.43434343434 0 -0.8 1e-06 
1.0 1.43434343434 0 -0.8 1e-06 
0.5 1.47474747475 0 -0.8 1e-06 
0.555555555556 1.47474747475 0 -0.8 1e-06 
0.611111111111 1.47474747475 0 -0.8 1e-06 
0.666666666667 1.47474747475 0 -0.8 1e-06 
0.722222222222 1.47474747475 0 -0.8 1e-06 
0.777777777778 1.47474747475 0 -0.8 1e-06 
0.833333333333 1.47474747475 0 -0.8 1e-06 
0.888888888889 1.47474747475 0 -0.8 1e-06 
0.944444444444 1.47474747475 0 -0.8 1e-06 
1.0 1.47474747475 0 -0.8 1e-06 
0.5 1.51515151515 0 -0.8 1e-06 
0.555555555556 1.51515151515 0 -0.8 1e-06 
0.611111111111 1.51515151515 0 -0.8 1e-06 
0.666666666667 1.51515151515 0 -0.8 1e-06 
0.722222222222 1.51515151515 0 -0.8 1e-06 
0.777777777778 1.51515151515 0 -0.8 1e-06 
0.833333333333 1.51515151515 0 -0.8 1e-06 
0.888888888889 1.51515151515 0 -0.8 1e-06 
0.944444444444 1.51515151515 0 -0.8 1e-06 
1.0 1.51515151515 0 -0.8 1e-06 
0.5 1.55555555556 0 -0.8 1e-06 
0.555555555556 1.55555555556 0 -0.8 1e-06 
0.611111111111 1.55555555556 0 -0.8 1e-06 
0.666666666667 1.55555555556 0 -0.8 1e-06 
0.722222222222 1.55555555556 0 -0.8 1e-06 
0.777777777778 1.55555555556 0 -0.8 1e-06 
0.833333333333 1.55555555556 0 -0.8 1e-06 
0.888888888889 1.55555555556 0 -0.8 1e-06 
0.944444444444 1.55555555556 0 -0.8 1e-06 
1.0 1.55555555556 0 -0.8 1e-06 
0.5 1.59595959596 0 -0.8 1e-06 
0.555555555556 1.59595959596 0 -0.8 1e-06 
0.611111111111 1.59595959596 0 -0.8 1e-06 
0.666666666667 1.59595959596 0 -0.8 1e-06 
0.722222222222 1.59595959596 0 -0.8 1e-06 
0.777777777778 1.59595959596 0 -0.8 1e-06 
0.833333333333 1.59595959596 0 -0.8 1e-06 
0.888888888889 1.59595959596 0 -0.8 1e-06 
0.944444444444 1.59595959596 0 -0.8 1e-06 
1.0 1.59595959596 0 -0.8 1e-06 
0.5 1.63636363636 0 -0.8 1e-06 
0.555555555556 1.63636363636 0 -0.8 1e-06 
0.611111111111 1.63636363636 0 -0.8 1e-06 
0.666666666667 1.63636363636 0 -0.8 1e-06 
0.722222222222 1.63636363636 0 -0.8 1e-06 
0.777777777778 1.63636363636 0 -0.8 1e-06 
0.833333333333 1.63636363636 0 -0.8 1e-06 
0.888888888889 1.63636363636 0 -0.8 1e-06 
0.944444444444 1.63636363636 0 -0.8 1e-06 
1.0 1.63636363636 0 -0.8 1e-06 
0.5 1.67676767677 0 -0.8 1e-06 
0.555555555556 1.67676767677 0 -0.8 1e-06 
0.611111111111 1.67676767677 0 -0.8 1e-06 
0.666666666667 1.67676767677 0 -0.8 1e-06 
0.722222222222 1.67676767677 0 -0.8 1e-06 
0.777777777778 1.67676767677 0 -0.8 1e-06 
0.833333333333 1.67676767677 0 -0.8 1e-06 
0.888888888889 1.67676767677 0 -0.8 1e-06 
0.944444444444 1.67676767677 0 -0.8 1e-06 
1.0 1.67676767677 0 -0.8 1e-06 
0.5 1.71717171717 0 -0.8 1e-06 
0.555555555556 1.71717171717 0 -0.8 1e-06 
0.611111111111 1.71717171717 0 -0.8 1e-06 
0.666666666667 1.71717171717 0 -0.8 1e-06 
0.722222222222 1.71717171717 0 -0.8 1e-06 
0.777777777778 1.71717171717 0 -0.8 1e-06 
0.833333333333 1.71717171717 0 -0.8 1e-06 
0.888888888889 1.71717171717 0 -0.8 1e-06 
0.944444444444 1.71717171717 0 -0.8 1e-06 
1.0 1.71717171717 0 -0.8 1e-06 
0.5 1.75757575758 0 -0.8 1e-06 
0.555555555556 1.75757575758 0 -0.8 1e-06 
0.611111111111 1.75757575758 0 -0.8 1e-06 
0.666666666667 1.75757575758 0 -0.8 1e-06 
0.722222222222 1.75757575758 0 -0.8 1e-06 
0.777777777778 1.75757575758 0 -0.8 1e-06 
0.833333333333 1.75757575758 0 -0.8 1e-06 
0.888888888889 1.75757575758 0 -0.8 1e-06 
0.944444444444 1.75757575758 0 -0.8 1e-06 
1.0 1.75757575758 0 -0.8 1e-06 
0.5 1.79797979798 0 -0.8 1e-06 
0.555555555556 1.79797979798 0 -0.8 1e-06 
0.611111111111 1.79797979798 0 -0.8 1e-06 
0.666666666667 1.79797979798 0 -0.8 1e-06 
0.722222222222 1.79797979798 0 -0.8 1e-06 
0.777777777778 1.79797979798 0 -0.8 1e-06 
0.833333333333 1.79797979798 0 -0.8 1e-06 
0.888888888889 1.79797979798 0 -0.8 1e-06 
0.944444444444 1.79797979798 0 -0.8 1e-06 
1.0 1.79797979798 0 -0.8 1e-06 
0.5 1.83838383838 0 -0.8 1e-06 
0.555555555556 1.83838383838 0 -0.8 1e-06 
0.611111111111 1.83838383838 0 -0.8 1e-06 
0.666666666667 1.83838383838 0 -0.8 1e-06 
0.722222222222 1.83838383838 0 -0.8 1e-06 
0.777777777778 1.83838383838 0 -0.8 1e-06 
0.833333333333 1.83838383838 0 -0.8 1e-06 
0.888888888889 1.83838383838 0 -0.8 1e-06 
0.944444444444 1.83838383838 0 -0.8 1e-06 
1.0 1.83838383838 0 -0.8 1e-06 
0.5 1.87878787879 0 -0.8 1e-06 
0.555555555556 1.87878787879 0 -0.8 1e-06 
0.611111111111 1.87878787879 0 -0.8 1e-06 
0.666666666667 1.87878787879 0 -0.8 1e-06 
0.722222222222 1.87878787879 0 -0.8 1e-06 
0.777777777778 1.87878787879 0 -0.8 1e-06 
0.833333333333 1.87878787879 0 -0.8 1e-06 
0.888888888889 1.87878787879 0 -0.8 1e-06 
0.944444444444 1.87878787879 0 -0.8 1e-06 
1.0 1.87878787879 0 -0.8 1e-06 
0.5 1.91919191919 0 -0.8 1e-06 
0.555555555556 1.91919191919 0 -0.8 1e-06 
0.611111111111 1.91919191919 0 -0.8 1e-06 
0.666666666667 1.91919191919 0 -0.8 1e-06 
0.722222222222 1.91919191919 0 -0.8 1e-06 
0.777777777778 1.91919191919 0 -0.8 1e-06 
0.833333333333 1.91919191919 0 -0.8 1e-06 
0.888888888889 1.91919191919 0 -0.8 1e-06 
0.944444444444 1.91919191919 0 -0.8 1e-06 
1.0 1.91919191919 0 -0.8 1e-06 
0.5 1.9595959596 0 -0.8 1e-06 
0.555555555556 1.9595959596 0 -0.8 1e-06 
0.611111111111 1.9595959596 0 -0.8 1e-06 
0.666666666667 1.9595959596 0 -0.8 1e-06 
0.722222222222 1.9595959596 0 -0.8 1e-06 
0.777777777778 1.9595959596 0 -0.8 1e-06 
0.833333333333 1.9595959596 0 -0.8 1e-06 
0.888888888889 1.9595959596 0 -0.8 1e-06 
0.944444444444 1.9595959596 0 -0.8 1e-06 
1.0 1.9595959596 0 -0.8 1e-06 
0.5 2.0 0 -0.8 1e-06 
0.555555555556 2.0 0 -0.8 1e-06 
0.611111111111 2.0 0 -0.8 1e-06 
0.666666666667 2.0 0 -0.8 1e-06 
0.722222222222 2.0 0 -0.8 1e-06 
0.777777777778 2.0 0 -0.8 1e-06 
0.833333333333 2.0 0 -0.8 1e-06 
0.888888888889 2.0 0 -0.8 1e-06 
0.944444444444 2.0 0 -0.8 1e-06 
1.0 2.0 0 -0.8 1e-06 
0.5 -2.0 0 -0.4 1e-06 
0.555555555556 -2.0 0 -0.4 1e-06 
0.611111111111 -2.0 0 -0.4 1e-06 
0.666666666667 -2.0 0 -0.4 1e-06 
0.722222222222 -2.0 0 -0.4 1e-06 
0.777777777778 -2.0 0 -0.4 1e-06 
0.833333333333 -2.0 0 -0.4 1e-06 
0.888888888889 -2.0 0 -0.4 1e-06 
0.944444444444 -2.0 0 -0.4 1e-06 
1.0 -2.0 0 -0.4 1e-06 
0.5 -1.9595959596 0 -0.4 1e-06 
0.555555555556 -1.9595959596 0 -0.4 1e-06 
0.611111111111 -1.9595959596 0 -0.4 1e-06 
0.666666666667 -1.9595959596 0 -0.4 1e-06 
0.722222222222 -1.9595959596 0 -0.4 1e-06 
0.777777777778 -1.9595959596 0 -0.4 1e-06 
0.833333333333 -1.9595959596 0 -0.4 1e-06 
0.888888888889 -1.9595959596 0 -0.4 1e-06 
0.944444444444 -1.9595959596 0 -0.4 1e-06 
1.0 -1.9595959596 0 -0.4 1e-06 
0.5 -1.91919191919 0 -0.4 1e-06 
0.555555555556 -1.91919191919 0 -0.4 1e-06 
0.611111111111 -1.91919191919 0 -0.4 1e-06 
0.666666666667 -1.91919191919 0 -0.4 1e-06 
0.722222222222 -1.91919191919 0 -0.4 1e-06 
0.777777777778 -1.91919191919 0 -0.4 1e-06 
0.833333333333 -1.91919191919 0 -0.4 1e-06 
0.888888888889 -1.91919191919 0 -0.4 1e-06 
0.944444444444 -1.91919191919 0 -0.4 1e-06 
1.0 -1.91919191919 0 -0.4 1e-06 
0.5 -1.87878787879 0 -0.4 1e-06 
0.555555555556 -1.87878787879 0 -0.4 1e-06 
0.611111111111 -1.87878787879 0 -0.4 1e-06 
0.666666666667 -1.87878787879 0 -0.4 1e-06 
0.722222222222 -1.87878787879 0 -0.4 1e-06 
0.777777777778 -1.87878787879 0 -0.4 1e-06 
0.833333333333 -1.87878787879 0 -0.4 1e-06 
0.888888888889 -1.87878787879 0 -0.4 1e-06 
0.944444444444 -1.87878787879 0 -0.4 1e-06 
1.0 -1.87878787879 0 -0.4 1e-06 
0.5 -1.83838383838 0 -0.4 1e-06 
0.555555555556 -1.83838383838 0 -0.4 1e-06 
0.611111111111 -1.83838383838 0 -0.4 1e-06 
0.666666666667 -1.83838383838 0 -0.4 1e-06 
0.722222222222 -1.83838383838 0 -0.4 1e-06 
0.777777777778 -1.83838383838 0 -0.4 1e-06 
0.833333333333 -1.83838383838 0 -0.4 1e-06 
0.888888888889 -1.83838383838 0 -0.4 1e-06 
0.944444444444 -1.83838383838 0 -0.4 1e-06 
1.0 -1.83838383838 0 -0.4 1e-06 
0.5 -1.79797979798 0 -0.4 1e-06 
0.555555555556 -1.79797979798 0 -0.4 1e-06 
0.611111111111 -1.79797979798 0 -0.4 1e-06 
0.666666666667 -1.79797979798 0 -0.4 1e-06 
0.722222222222 -1.79797979798 0 -0.4 1e-06 
0.777777777778 -1.79797979798 0 -0.4 1e-06 
0.833333333333 -1.79797979798 0 -0.4 1e-06 
0.888888888889 -1.79797979798 0 -0.4 1e-06 
0.944444444444 -1.79797979798 0 -0.4 1e-06 
1.0 -1.79797979798 0 -0.4 1e-06 
0.5 -1.75757575758 0 -0.4 1e-06 
0.555555555556 -1.75757575758 0 -0.4 1e-06 
0.611111111111 -1.75757575758 0 -0.4 1e-06 
0.666666666667 -1.75757575758 0 -0.4 1e-06 
0.722222222222 -1.75757575758 0 -0.4 1e-06 
0.777777777778 -1.75757575758 0 -0.4 1e-06 
0.833333333333 -1.75757575758 0 -0.4 1e-06 
0.888888888889 -1.75757575758 0 -0.4 1e-06 
0.944444444444 -1.75757575758 0 -0.4 1e-06 
1.0 -1.75757575758 0 -0.4 1e-06 
0.5 -1.71717171717 0 -0.4 1e-06 
0.555555555556 -1.71717171717 0 -0.4 1e-06 
0.611111111111 -1.71717171717 0 -0.4 1e-06 
0.666666666667 -1.71717171717 0 -0.4 1e-06 
0.722222222222 -1.71717171717 0 -0.4 1e-06 
0.777777777778 -1.71717171717 0 -0.4 1e-06 
0.833333333333 -1.71717171717 0 -0.4 1e-06 
0.888888888889 -1.71717171717 0 -0.4 1e-06 
0.944444444444 -1.71717171717 0 -0.4 1e-06 
1.0 -1.71717171717 0 -0.4 1e-06 
0.5 -1.67676767677 0 -0.4 1e-06 
0.555555555556 -1.67676767677 0 -0.4 1e-06 
0.611111111111 -1.67676767677 0 -0.4 1e-06 
0.666666666667 -1.67676767677 0 -0.4 1e-06 
0.722222222222 -1.67676767677 0 -0.4 1e-06 
0.777777777778 -1.67676767677 0 -0.4 1e-06 
0.833333333333 -1.67676767677 0 -0.4 1e-06 
0.888888888889 -1.67676767677 0 -0.4 1e-06 
0.944444444444 -1.67676767677 0 -0.4 1e-06 
1.0 -1.67676767677 0 -0.4 1e-06 
0.5 -1.63636363636 0 -0.4 1e-06 
0.555555555556 -1.63636363636 0 -0.4 1e-06 
0.611111111111 -1.63636363636 0 -0.4 1e-06 
0.666666666667 -1.63636363636 0 -0.4 1e-06 
0.722222222222 -1.63636363636 0 -0.4 1e-06 
0.777777777778 -1.63636363636 0 -0.4 1e-06 
0.833333333333 -1.63636363636 0 -0.4 1e-06 
0.888888888889 -1.63636363636 0 -0.4 1e-06 
0.944444444444 -1.63636363636 0 -0.4 1e-06 
1.0 -1.63636363636 0 -0.4 1e-06 
0.5 -1.59595959596 0 -0.4 1e-06 
0.555555555556 -1.59595959596 0 -0.4 1e-06 
0.611111111111 -1.59595959596 0 -0.4 1e-06 
0.666666666667 -1.59595959596 0 -0.4 1e-06 
0.722222222222 -1.59595959596 0 -0.4 1e-06 
0.777777777778 -1.59595959596 0 -0.4 1e-06 
0.833333333333 -1.59595959596 0 -0.4 1e-06 
0.888888888889 -1.59595959596 0 -0.4 1e-06 
0.944444444444 -1.59595959596 0 -0.4 1e-06 
1.0 -1.59595959596 0 -0.4 1e-06 
0.5 -1.55555555556 0 -0.4 1e-06 
0.555555555556 -1.55555555556 0 -0.4 1e-06 
0.611111111111 -1.55555555556 0 -0.4 1e-06 
0.666666666667 -1.55555555556 0 -0.4 1e-06 
0.722222222222 -1.55555555556 0 -0.4 1e-06 
0.777777777778 -1.55555555556 0 -0.4 1e-06 
0.833333333333 -1.55555555556 0 -0.4 1e-06 
0.888888888889 -1.55555555556 0 -0.4 1e-06 
0.944444444444 -1.55555555556 0 -0.4 1e-06 
1.0 -1.55555555556 0 -0.4 1e-06 
0.5 -1.51515151515 0 -0.4 1e-06 
0.555555555556 -1.51515151515 0 -0.4 1e-06 
0.611111111111 -1.51515151515 0 -0.4 1e-06 
0.666666666667 -1.51515151515 0 -0.4 1e-06 
0.722222222222 -1.51515151515 0 -0.4 1e-06 
0.777777777778 -1.51515151515 0 -0.4 1e-06 
0.833333333333 -1.51515151515 0 -0.4 1e-06 
0.888888888889 -1.51515151515 0 -0.4 1e-06 
0.944444444444 -1.51515151515 0 -0.4 1e-06 
1.0 -1.51515151515 0 -0.4 1e-06 
0.5 -1.47474747475 0 -0.4 1e-06 
0.555555555556 -1.47474747475 0 -0.4 1e-06 
0.611111111111 -1.47474747475 0 -0.4 1e-06 
0.666666666667 -1.47474747475 0 -0.4 1e-06 
0.722222222222 -1.47474747475 0 -0.4 1e-06 
0.777777777778 -1.47474747475 0 -0.4 1e-06 
0.833333333333 -1.47474747475 0 -0.4 1e-06 
0.888888888889 -1.47474747475 0 -0.4 1e-06 
0.944444444444 -1.47474747475 0 -0.4 1e-06 
1.0 -1.47474747475 0 -0.4 1e-06 
0.5 -1.43434343434 0 -0.4 1e-06 
0.555555555556 -1.43434343434 0 -0.4 1e-06 
0.611111111111 -1.43434343434 0 -0.4 1e-06 
0.666666666667 -1.43434343434 0 -0.4 1e-06 
0.722222222222 -1.43434343434 0 -0.4 1e-06 
0.777777777778 -1.43434343434 0 -0.4 1e-06 
0.833333333333 -1.43434343434 0 -0.4 1e-06 
0.888888888889 -1.43434343434 0 -0.4 1e-06 
0.944444444444 -1.43434343434 0 -0.4 1e-06 
1.0 -1.43434343434 0 -0.4 1e-06 
0.5 -1.39393939394 0 -0.4 1e-06 
0.555555555556 -1.39393939394 0 -0.4 1e-06 
0.611111111111 -1.39393939394 0 -0.4 1e-06 
0.666666666667 -1.39393939394 0 -0.4 1e-06 
0.722222222222 -1.39393939394 0 -0.4 1e-06 
0.777777777778 -1.39393939394 0 -0.4 1e-06 
0.833333333333 -1.39393939394 0 -0.4 1e-06 
0.888888888889 -1.39393939394 0 -0.4 1e-06 
0.944444444444 -1.39393939394 0 -0.4 1e-06 
1.0 -1.39393939394 0 -0.4 1e-06 
0.5 -1.35353535354 0 -0.4 1e-06 
0.555555555556 -1.35353535354 0 -0.4 1e-06 
0.611111111111 -1.35353535354 0 -0.4 1e-06 
0.666666666667 -1.35353535354 0 -0.4 1e-06 
0.722222222222 -1.35353535354 0 -0.4 1e-06 
0.777777777778 -1.35353535354 0 -0.4 1e-06 
0.833333333333 -1.35353535354 0 -0.4 1e-06 
0.888888888889 -1.35353535354 0 -0.4 1e-06 
0.944444444444 -1.35353535354 0 -0.4 1e-06 
1.0 -1.35353535354 0 -0.4 1e-06 
0.5 -1.31313131313 0 -0.4 1e-06 
0.555555555556 -1.31313131313 0 -0.4 1e-06 
0.611111111111 -1.31313131313 0 -0.4 1e-06 
0.666666666667 -1.31313131313 0 -0.4 1e-06 
0.722222222222 -1.31313131313 0 -0.4 1e-06 
0.777777777778 -1.31313131313 0 -0.4 1e-06 
0.833333333333 -1.31313131313 0 -0.4 1e-06 
0.888888888889 -1.31313131313 0 -0.4 1e-06 
0.944444444444 -1.31313131313 0 -0.4 1e-06 
1.0 -1.31313131313 0 -0.4 1e-06 
0.5 -1.27272727273 0 -0.4 1e-06 
0.555555555556 -1.27272727273 0 -0.4 1e-06 
0.611111111111 -1.27272727273 0 -0.4 1e-06 
0.666666666667 -1.27272727273 0 -0.4 1e-06 
0.722222222222 -1.27272727273 0 -0.4 1e-06 
0.777777777778 -1.27272727273 0 -0.4 1e-06 
0.833333333333 -1.27272727273 0 -0.4 1e-06 
0.888888888889 -1.27272727273 0 -0.4 1e-06 
0.944444444444 -1.27272727273 0 -0.4 1e-06 
1.0 -1.27272727273 0 -0.4 1e-06 
0.5 -1.23232323232 0 -0.4 1e-06 
0.555555555556 -1.23232323232 0 -0.4 1e-06 
0.611111111111 -1.23232323232 0 -0.4 1e-06 
0.666666666667 -1.23232323232 0 -0.4 1e-06 
0.722222222222 -1.23232323232 0 -0.4 1e-06 
0.777777777778 -1.23232323232 0 -0.4 1e-06 
0.833333333333 -1.23232323232 0 -0.4 1e-06 
0.888888888889 -1.23232323232 0 -0.4 1e-06 
0.944444444444 -1.23232323232 0 -0.4 1e-06 
1.0 -1.23232323232 0 -0.4 1e-06 
0.5 -1.19191919192 0 -0.4 1e-06 
0.555555555556 -1.19191919192 0 -0.4 1e-06 
0.611111111111 -1.19191919192 0 -0.4 1e-06 
0.666666666667 -1.19191919192 0 -0.4 1e-06 
0.722222222222 -1.19191919192 0 -0.4 1e-06 
0.777777777778 -1.19191919192 0 -0.4 1e-06 
0.833333333333 -1.19191919192 0 -0.4 1e-06 
0.888888888889 -1.19191919192 0 -0.4 1e-06 
0.944444444444 -1.19191919192 0 -0.4 1e-06 
1.0 -1.19191919192 0 -0.4 1e-06 
0.5 -1.15151515152 0 -0.4 1e-06 
0.555555555556 -1.15151515152 0 -0.4 1e-06 
0.611111111111 -1.15151515152 0 -0.4 1e-06 
0.666666666667 -1.15151515152 0 -0.4 1e-06 
0.722222222222 -1.15151515152 0 -0.4 1e-06 
0.777777777778 -1.15151515152 0 -0.4 1e-06 
0.833333333333 -1.15151515152 0 -0.4 1e-06 
0.888888888889 -1.15151515152 0 -0.4 1e-06 
0.944444444444 -1.15151515152 0 -0.4 1e-06 
1.0 -1.15151515152 0 -0.4 1e-06 
0.5 -1.11111111111 0 -0.4 1e-06 
0.555555555556 -1.11111111111 0 -0.4 1e-06 
0.611111111111 -1.11111111111 0 -0.4 1e-06 
0.666666666667 -1.11111111111 0 -0.4 1e-06 
0.722222222222 -1.11111111111 0 -0.4 1e-06 
0.777777777778 -1.11111111111 0 -0.4 1e-06 
0.833333333333 -1.11111111111 0 -0.4 1e-06 
0.888888888889 -1.11111111111 0 -0.4 1e-06 
0.944444444444 -1.11111111111 0 -0.4 1e-06 
1.0 -1.11111111111 0 -0.4 1e-06 
0.5 -1.07070707071 0 -0.4 1e-06 
0.555555555556 -1.07070707071 0 -0.4 1e-06 
0.611111111111 -1.07070707071 0 -0.4 1e-06 
0.666666666667 -1.07070707071 0 -0.4 1e-06 
0.722222222222 -1.07070707071 0 -0.4 1e-06 
0.777777777778 -1.07070707071 0 -0.4 1e-06 
0.833333333333 -1.07070707071 0 -0.4 1e-06 
0.888888888889 -1.07070707071 0 -0.4 1e-06 
0.944444444444 -1.07070707071 0 -0.4 1e-06 
1.0 -1.07070707071 0 -0.4 1e-06 
0.5 -1.0303030303 0 -0.4 1e-06 
0.555555555556 -1.0303030303 0 -0.4 1e-06 
0.611111111111 -1.0303030303 0 -0.4 1e-06 
0.666666666667 -1.0303030303 0 -0.4 1e-06 
0.722222222222 -1.0303030303 0 -0.4 1e-06 
0.777777777778 -1.0303030303 0 -0.4 1e-06 
0.833333333333 -1.0303030303 0 -0.4 1e-06 
0.888888888889 -1.0303030303 0 -0.4 1e-06 
0.944444444444 -1.0303030303 0 -0.4 1e-06 
1.0 -1.0303030303 0 -0.4 1e-06 
0.5 -0.989898989899 0 -0.4 1e-06 
0.555555555556 -0.989898989899 0 -0.4 1e-06 
0.611111111111 -0.989898989899 0 -0.4 1e-06 
0.666666666667 -0.989898989899 0 -0.4 1e-06 
0.722222222222 -0.989898989899 0 -0.4 1e-06 
0.777777777778 -0.989898989899 0 -0.4 1e-06 
0.833333333333 -0.989898989899 0 -0.4 1e-06 
0.888888888889 -0.989898989899 0 -0.4 1e-06 
0.944444444444 -0.989898989899 0 -0.4 1e-06 
1.0 -0.989898989899 0 -0.4 1e-06 
0.5 -0.949494949495 0 -0.4 1e-06 
0.555555555556 -0.949494949495 0 -0.4 1e-06 
0.611111111111 -0.949494949495 0 -0.4 1e-06 
0.666666666667 -0.949494949495 0 -0.4 1e-06 
0.722222222222 -0.949494949495 0 -0.4 1e-06 
0.777777777778 -0.949494949495 0 -0.4 1e-06 
0.833333333333 -0.949494949495 0 -0.4 1e-06 
0.888888888889 -0.949494949495 0 -0.4 1e-06 
0.944444444444 -0.949494949495 0 -0.4 1e-06 
1.0 -0.949494949495 0 -0.4 1e-06 
0.5 -0.909090909091 0 -0.4 1e-06 
0.555555555556 -0.909090909091 0 -0.4 1e-06 
0.611111111111 -0.909090909091 0 -0.4 1e-06 
0.666666666667 -0.909090909091 0 -0.4 1e-06 
0.722222222222 -0.909090909091 0 -0.4 1e-06 
0.777777777778 -0.909090909091 0 -0.4 1e-06 
0.833333333333 -0.909090909091 0 -0.4 1e-06 
0.888888888889 -0.909090909091 0 -0.4 1e-06 
0.944444444444 -0.909090909091 0 -0.4 1e-06 
1.0 -0.909090909091 0 -0.4 1e-06 
0.5 -0.868686868687 0 -0.4 1e-06 
0.555555555556 -0.868686868687 0 -0.4 1e-06 
0.611111111111 -0.868686868687 0 -0.4 1e-06 
0.666666666667 -0.868686868687 0 -0.4 1e-06 
0.722222222222 -0.868686868687 0 -0.4 1e-06 
0.777777777778 -0.868686868687 0 -0.4 1e-06 
0.833333333333 -0.868686868687 0 -0.4 1e-06 
0.888888888889 -0.868686868687 0 -0.4 1e-06 
0.944444444444 -0.868686868687 0 -0.4 1e-06 
1.0 -0.868686868687 0 -0.4 1e-06 
0.5 -0.828282828283 0 -0.4 1e-06 
0.555555555556 -0.828282828283 0 -0.4 1e-06 
0.611111111111 -0.828282828283 0 -0.4 1e-06 
0.666666666667 -0.828282828283 0 -0.4 1e-06 
0.722222222222 -0.828282828283 0 -0.4 1e-06 
0.777777777778 -0.828282828283 0 -0.4 1e-06 
0.833333333333 -0.828282828283 0 -0.4 1e-06 
0.888888888889 -0.828282828283 0 -0.4 1e-06 
0.944444444444 -0.828282828283 0 -0.4 1e-06 
1.0 -0.828282828283 0 -0.4 1e-06 
0.5 -0.787878787879 0 -0.4 1e-06 
0.555555555556 -0.787878787879 0 -0.4 1e-06 
0.611111111111 -0.787878787879 0 -0.4 1e-06 
0.666666666667 -0.787878787879 0 -0.4 1e-06 
0.722222222222 -0.787878787879 0 -0.4 1e-06 
0.777777777778 -0.787878787879 0 -0.4 1e-06 
0.833333333333 -0.787878787879 0 -0.4 1e-06 
0.888888888889 -0.787878787879 0 -0.4 1e-06 
0.944444444444 -0.787878787879 0 -0.4 1e-06 
1.0 -0.787878787879 0 -0.4 1e-06 
0.5 -0.747474747475 0 -0.4 1e-06 
0.555555555556 -0.747474747475 0 -0.4 1e-06 
0.611111111111 -0.747474747475 0 -0.4 1e-06 
0.666666666667 -0.747474747475 0 -0.4 1e-06 
0.722222222222 -0.747474747475 0 -0.4 1e-06 
0.777777777778 -0.747474747475 0 -0.4 1e-06 
0.833333333333 -0.747474747475 0 -0.4 1e-06 
0.888888888889 -0.747474747475 0 -0.4 1e-06 
0.944444444444 -0.747474747475 0 -0.4 1e-06 
1.0 -0.747474747475 0 -0.4 1e-06 
0.5 -0.707070707071 0 -0.4 1e-06 
0.555555555556 -0.707070707071 0 -0.4 1e-06 
0.611111111111 -0.707070707071 0 -0.4 1e-06 
0.666666666667 -0.707070707071 0 -0.4 1e-06 
0.722222222222 -0.707070707071 0 -0.4 1e-06 
0.777777777778 -0.707070707071 0 -0.4 1e-06 
0.833333333333 -0.707070707071 0 -0.4 1e-06 
0.888888888889 -0.707070707071 0 -0.4 1e-06 
0.944444444444 -0.707070707071 0 -0.4 1e-06 
1.0 -0.707070707071 0 -0.4 1e-06 
0.5 -0.666666666667 0 -0.4 1e-06 
0.555555555556 -0.666666666667 0 -0.4 1e-06 
0.611111111111 -0.666666666667 0 -0.4 1e-06 
0.666666666667 -0.666666666667 0 -0.4 1e-06 
0.722222222222 -0.666666666667 0 -0.4 1e-06 
0.777777777778 -0.666666666667 0 -0.4 1e-06 
0.833333333333 -0.666666666667 0 -0.4 1e-06 
0.888888888889 -0.666666666667 0 -0.4 1e-06 
0.944444444444 -0.666666666667 0 -0.4 1e-06 
1.0 -0.666666666667 0 -0.4 1e-06 
0.5 -0.626262626263 0 -0.4 1e-06 
0.555555555556 -0.626262626263 0 -0.4 1e-06 
0.611111111111 -0.626262626263 0 -0.4 1e-06 
0.666666666667 -0.626262626263 0 -0.4 1e-06 
0.722222222222 -0.626262626263 0 -0.4 1e-06 
0.777777777778 -0.626262626263 0 -0.4 1e-06 
0.833333333333 -0.626262626263 0 -0.4 1e-06 
0.888888888889 -0.626262626263 0 -0.4 1e-06 
0.944444444444 -0.626262626263 0 -0.4 1e-06 
1.0 -0.626262626263 0 -0.4 1e-06 
0.5 -0.585858585859 0 -0.4 1e-06 
0.555555555556 -0.585858585859 0 -0.4 1e-06 
0.611111111111 -0.585858585859 0 -0.4 1e-06 
0.666666666667 -0.585858585859 0 -0.4 1e-06 
0.722222222222 -0.585858585859 0 -0.4 1e-06 
0.777777777778 -0.585858585859 0 -0.4 1e-06 
0.833333333333 -0.585858585859 0 -0.4 1e-06 
0.888888888889 -0.585858585859 0 -0.4 1e-06 
0.944444444444 -0.585858585859 0 -0.4 1e-06 
1.0 -0.585858585859 0 -0.4 1e-06 
0.5 -0.545454545455 0 -0.4 1e-06 
0.555555555556 -0.545454545455 0 -0.4 1e-06 
0.611111111111 -0.545454545455 0 -0.4 1e-06 
0.666666666667 -0.545454545455 0 -0.4 1e-06 
0.722222222222 -0.545454545455 0 -0.4 1e-06 
0.777777777778 -0.545454545455 0 -0.4 1e-06 
0.833333333333 -0.545454545455 0 -0.4 1e-06 
0.888888888889 -0.545454545455 0 -0.4 1e-06 
0.944444444444 -0.545454545455 0 -0.4 1e-06 
1.0 -0.545454545455 0 -0.4 1e-06 
0.5 -0.505050505051 0 -0.4 1e-06 
0.555555555556 -0.505050505051 0 -0.4 1e-06 
0.611111111111 -0.505050505051 0 -0.4 1e-06 
0.666666666667 -0.505050505051 0 -0.4 1e-06 
0.722222222222 -0.505050505051 0 -0.4 1e-06 
0.777777777778 -0.505050505051 0 -0.4 1e-06 
0.833333333333 -0.505050505051 0 -0.4 1e-06 
0.888888888889 -0.505050505051 0 -0.4 1e-06 
0.944444444444 -0.505050505051 0 -0.4 1e-06 
1.0 -0.505050505051 0 -0.4 1e-06 
0.5 -0.464646464646 0 -0.4 1e-06 
0.555555555556 -0.464646464646 0 -0.4 1e-06 
0.611111111111 -0.464646464646 0 -0.4 1e-06 
0.666666666667 -0.464646464646 0 -0.4 1e-06 
0.722222222222 -0.464646464646 0 -0.4 1e-06 
0.777777777778 -0.464646464646 0 -0.4 1e-06 
0.833333333333 -0.464646464646 0 -0.4 1e-06 
0.888888888889 -0.464646464646 0 -0.4 1e-06 
0.944444444444 -0.464646464646 0 -0.4 1e-06 
1.0 -0.464646464646 0 -0.4 1e-06 
0.5 -0.424242424242 0 -0.4 1e-06 
0.555555555556 -0.424242424242 0 -0.4 1e-06 
0.611111111111 -0.424242424242 0 -0.4 1e-06 
0.666666666667 -0.424242424242 0 -0.4 1e-06 
0.722222222222 -0.424242424242 0 -0.4 1e-06 
0.777777777778 -0.424242424242 0 -0.4 1e-06 
0.833333333333 -0.424242424242 0 -0.4 1e-06 
0.888888888889 -0.424242424242 0 -0.4 1e-06 
0.944444444444 -0.424242424242 0 -0.4 1e-06 
1.0 -0.424242424242 0 -0.4 1e-06 
0.5 -0.383838383838 0 -0.4 1e-06 
0.555555555556 -0.383838383838 0 -0.4 1e-06 
0.611111111111 -0.383838383838 0 -0.4 1e-06 
0.666666666667 -0.383838383838 0 -0.4 1e-06 
0.722222222222 -0.383838383838 0 -0.4 1e-06 
0.777777777778 -0.383838383838 0 -0.4 1e-06 
0.833333333333 -0.383838383838 0 -0.4 1e-06 
0.888888888889 -0.383838383838 0 -0.4 1e-06 
0.944444444444 -0.383838383838 0 -0.4 1e-06 
1.0 -0.383838383838 0 -0.4 1e-06 
0.5 -0.343434343434 0 -0.4 1e-06 
0.555555555556 -0.343434343434 0 -0.4 1e-06 
0.611111111111 -0.343434343434 0 -0.4 1e-06 
0.666666666667 -0.343434343434 0 -0.4 1e-06 
0.722222222222 -0.343434343434 0 -0.4 1e-06 
0.777777777778 -0.343434343434 0 -0.4 1e-06 
0.833333333333 -0.343434343434 0 -0.4 1e-06 
0.888888888889 -0.343434343434 0 -0.4 1e-06 
0.944444444444 -0.343434343434 0 -0.4 1e-06 
1.0 -0.343434343434 0 -0.4 1e-06 
0.5 -0.30303030303 0 -0.4 1e-06 
0.555555555556 -0.30303030303 0 -0.4 1e-06 
0.611111111111 -0.30303030303 0 -0.4 1e-06 
0.666666666667 -0.30303030303 0 -0.4 1e-06 
0.722222222222 -0.30303030303 0 -0.4 1e-06 
0.777777777778 -0.30303030303 0 -0.4 1e-06 
0.833333333333 -0.30303030303 0 -0.4 1e-06 
0.888888888889 -0.30303030303 0 -0.4 1e-06 
0.944444444444 -0.30303030303 0 -0.4 1e-06 
1.0 -0.30303030303 0 -0.4 1e-06 
0.5 -0.262626262626 0 -0.4 1e-06 
0.555555555556 -0.262626262626 0 -0.4 1e-06 
0.611111111111 -0.262626262626 0 -0.4 1e-06 
0.666666666667 -0.262626262626 0 -0.4 1e-06 
0.722222222222 -0.262626262626 0 -0.4 1e-06 
0.777777777778 -0.262626262626 0 -0.4 1e-06 
0.833333333333 -0.262626262626 0 -0.4 1e-06 
0.888888888889 -0.262626262626 0 -0.4 1e-06 
0.944444444444 -0.262626262626 0 -0.4 1e-06 
1.0 -0.262626262626 0 -0.4 1e-06 
0.5 -0.222222222222 0 -0.4 1e-06 
0.555555555556 -0.222222222222 0 -0.4 1e-06 
0.611111111111 -0.222222222222 0 -0.4 1e-06 
0.666666666667 -0.222222222222 0 -0.4 1e-06 
0.722222222222 -0.222222222222 0 -0.4 1e-06 
0.777777777778 -0.222222222222 0 -0.4 1e-06 
0.833333333333 -0.222222222222 0 -0.4 1e-06 
0.888888888889 -0.222222222222 0 -0.4 1e-06 
0.944444444444 -0.222222222222 0 -0.4 1e-06 
1.0 -0.222222222222 0 -0.4 1e-06 
0.5 -0.181818181818 0 -0.4 1e-06 
0.555555555556 -0.181818181818 0 -0.4 1e-06 
0.611111111111 -0.181818181818 0 -0.4 1e-06 
0.666666666667 -0.181818181818 0 -0.4 1e-06 
0.722222222222 -0.181818181818 0 -0.4 1e-06 
0.777777777778 -0.181818181818 0 -0.4 1e-06 
0.833333333333 -0.181818181818 0 -0.4 1e-06 
0.888888888889 -0.181818181818 0 -0.4 1e-06 
0.944444444444 -0.181818181818 0 -0.4 1e-06 
1.0 -0.181818181818 0 -0.4 1e-06 
0.5 -0.141414141414 0 -0.4 1e-06 
0.555555555556 -0.141414141414 0 -0.4 1e-06 
0.611111111111 -0.141414141414 0 -0.4 1e-06 
0.666666666667 -0.141414141414 0 -0.4 1e-06 
0.722222222222 -0.141414141414 0 -0.4 1e-06 
0.777777777778 -0.141414141414 0 -0.4 1e-06 
0.833333333333 -0.141414141414 0 -0.4 1e-06 
0.888888888889 -0.141414141414 0 -0.4 1e-06 
0.944444444444 -0.141414141414 0 -0.4 1e-06 
1.0 -0.141414141414 0 -0.4 1e-06 
0.5 -0.10101010101 0 -0.4 1e-06 
0.555555555556 -0.10101010101 0 -0.4 1e-06 
0.611111111111 -0.10101010101 0 -0.4 1e-06 
0.666666666667 -0.10101010101 0 -0.4 1e-06 
0.722222222222 -0.10101010101 0 -0.4 1e-06 
0.777777777778 -0.10101010101 0 -0.4 1e-06 
0.833333333333 -0.10101010101 0 -0.4 1e-06 
0.888888888889 -0.10101010101 0 -0.4 1e-06 
0.944444444444 -0.10101010101 0 -0.4 1e-06 
1.0 -0.10101010101 0 -0.4 1e-06 
0.5 -0.0606060606061 0 -0.4 1e-06 
0.555555555556 -0.0606060606061 0 -0.4 1e-06 
0.611111111111 -0.0606060606061 0 -0.4 1e-06 
0.666666666667 -0.0606060606061 0 -0.4 1e-06 
0.722222222222 -0.0606060606061 0 -0.4 1e-06 
0.777777777778 -0.0606060606061 0 -0.4 1e-06 
0.833333333333 -0.0606060606061 0 -0.4 1e-06 
0.888888888889 -0.0606060606061 0 -0.4 1e-06 
0.944444444444 -0.0606060606061 0 -0.4 1e-06 
1.0 -0.0606060606061 0 -0.4 1e-06 
0.5 -0.020202020202 0 -0.4 1e-06 
0.555555555556 -0.020202020202 0 -0.4 1e-06 
0.611111111111 -0.020202020202 0 -0.4 1e-06 
0.666666666667 -0.020202020202 0 -0.4 1e-06 
0.722222222222 -0.020202020202 0 -0.4 1e-06 
0.777777777778 -0.020202020202 0 -0.4 1e-06 
0.833333333333 -0.020202020202 0 -0.4 1e-06 
0.888888888889 -0.020202020202 0 -0.4 1e-06 
0.944444444444 -0.020202020202 0 -0.4 1e-06 
1.0 -0.020202020202 0 -0.4 1e-06 
0.5 0.020202020202 0 -0.4 1e-06 
0.555555555556 0.020202020202 0 -0.4 1e-06 
0.611111111111 0.020202020202 0 -0.4 1e-06 
0.666666666667 0.020202020202 0 -0.4 1e-06 
0.722222222222 0.020202020202 0 -0.4 1e-06 
0.777777777778 0.020202020202 0 -0.4 1e-06 
0.833333333333 0.020202020202 0 -0.4 1e-06 
0.888888888889 0.020202020202 0 -0.4 1e-06 
0.944444444444 0.020202020202 0 -0.4 1e-06 
1.0 0.020202020202 0 -0.4 1e-06 
0.5 0.0606060606061 0 -0.4 1e-06 
0.555555555556 0.0606060606061 0 -0.4 1e-06 
0.611111111111 0.0606060606061 0 -0.4 1e-06 
0.666666666667 0.0606060606061 0 -0.4 1e-06 
0.722222222222 0.0606060606061 0 -0.4 1e-06 
0.777777777778 0.0606060606061 0 -0.4 1e-06 
0.833333333333 0.0606060606061 0 -0.4 1e-06 
0.888888888889 0.0606060606061 0 -0.4 1e-06 
0.944444444444 0.0606060606061 0 -0.4 1e-06 
1.0 0.0606060606061 0 -0.4 1e-06 
0.5 0.10101010101 0 -0.4 1e-06 
0.555555555556 0.10101010101 0 -0.4 1e-06 
0.611111111111 0.10101010101 0 -0.4 1e-06 
0.666666666667 0.10101010101 0 -0.4 1e-06 
0.722222222222 0.10101010101 0 -0.4 1e-06 
0.777777777778 0.10101010101 0 -0.4 1e-06 
0.833333333333 0.10101010101 0 -0.4 1e-06 
0.888888888889 0.10101010101 0 -0.4 1e-06 
0.944444444444 0.10101010101 0 -0.4 1e-06 
1.0 0.10101010101 0 -0.4 1e-06 
0.5 0.141414141414 0 -0.4 1e-06 
0.555555555556 0.141414141414 0 -0.4 1e-06 
0.611111111111 0.141414141414 0 -0.4 1e-06 
0.666666666667 0.141414141414 0 -0.4 1e-06 
0.722222222222 0.141414141414 0 -0.4 1e-06 
0.777777777778 0.141414141414 0 -0.4 1e-06 
0.833333333333 0.141414141414 0 -0.4 1e-06 
0.888888888889 0.141414141414 0 -0.4 1e-06 
0.944444444444 0.141414141414 0 -0.4 1e-06 
1.0 0.141414141414 0 -0.4 1e-06 
0.5 0.181818181818 0 -0.4 1e-06 
0.555555555556 0.181818181818 0 -0.4 1e-06 
0.611111111111 0.181818181818 0 -0.4 1e-06 
0.666666666667 0.181818181818 0 -0.4 1e-06 
0.722222222222 0.181818181818 0 -0.4 1e-06 
0.777777777778 0.181818181818 0 -0.4 1e-06 
0.833333333333 0.181818181818 0 -0.4 1e-06 
0.888888888889 0.181818181818 0 -0.4 1e-06 
0.944444444444 0.181818181818 0 -0.4 1e-06 
1.0 0.181818181818 0 -0.4 1e-06 
0.5 0.222222222222 0 -0.4 1e-06 
0.555555555556 0.222222222222 0 -0.4 1e-06 
0.611111111111 0.222222222222 0 -0.4 1e-06 
0.666666666667 0.222222222222 0 -0.4 1e-06 
0.722222222222 0.222222222222 0 -0.4 1e-06 
0.777777777778 0.222222222222 0 -0.4 1e-06 
0.833333333333 0.222222222222 0 -0.4 1e-06 
0.888888888889 0.222222222222 0 -0.4 1e-06 
0.944444444444 0.222222222222 0 -0.4 1e-06 
1.0 0.222222222222 0 -0.4 1e-06 
0.5 0.262626262626 0 -0.4 1e-06 
0.555555555556 0.262626262626 0 -0.4 1e-06 
0.611111111111 0.262626262626 0 -0.4 1e-06 
0.666666666667 0.262626262626 0 -0.4 1e-06 
0.722222222222 0.262626262626 0 -0.4 1e-06 
0.777777777778 0.262626262626 0 -0.4 1e-06 
0.833333333333 0.262626262626 0 -0.4 1e-06 
0.888888888889 0.262626262626 0 -0.4 1e-06 
0.944444444444 0.262626262626 0 -0.4 1e-06 
1.0 0.262626262626 0 -0.4 1e-06 
0.5 0.30303030303 0 -0.4 1e-06 
0.555555555556 0.30303030303 0 -0.4 1e-06 
0.611111111111 0.30303030303 0 -0.4 1e-06 
0.666666666667 0.30303030303 0 -0.4 1e-06 
0.722222222222 0.30303030303 0 -0.4 1e-06 
0.777777777778 0.30303030303 0 -0.4 1e-06 
0.833333333333 0.30303030303 0 -0.4 1e-06 
0.888888888889 0.30303030303 0 -0.4 1e-06 
0.944444444444 0.30303030303 0 -0.4 1e-06 
1.0 0.30303030303 0 -0.4 1e-06 
0.5 0.343434343434 0 -0.4 1e-06 
0.555555555556 0.343434343434 0 -0.4 1e-06 
0.611111111111 0.343434343434 0 -0.4 1e-06 
0.666666666667 0.343434343434 0 -0.4 1e-06 
0.722222222222 0.343434343434 0 -0.4 1e-06 
0.777777777778 0.343434343434 0 -0.4 1e-06 
0.833333333333 0.343434343434 0 -0.4 1e-06 
0.888888888889 0.343434343434 0 -0.4 1e-06 
0.944444444444 0.343434343434 0 -0.4 1e-06 
1.0 0.343434343434 0 -0.4 1e-06 
0.5 0.383838383838 0 -0.4 1e-06 
0.555555555556 0.383838383838 0 -0.4 1e-06 
0.611111111111 0.383838383838 0 -0.4 1e-06 
0.666666666667 0.383838383838 0 -0.4 1e-06 
0.722222222222 0.383838383838 0 -0.4 1e-06 
0.777777777778 0.383838383838 0 -0.4 1e-06 
0.833333333333 0.383838383838 0 -0.4 1e-06 
0.888888888889 0.383838383838 0 -0.4 1e-06 
0.944444444444 0.383838383838 0 -0.4 1e-06 
1.0 0.383838383838 0 -0.4 1e-06 
0.5 0.424242424242 0 -0.4 1e-06 
0.555555555556 0.424242424242 0 -0.4 1e-06 
0.611111111111 0.424242424242 0 -0.4 1e-06 
0.666666666667 0.424242424242 0 -0.4 1e-06 
0.722222222222 0.424242424242 0 -0.4 1e-06 
0.777777777778 0.424242424242 0 -0.4 1e-06 
0.833333333333 0.424242424242 0 -0.4 1e-06 
0.888888888889 0.424242424242 0 -0.4 1e-06 
0.944444444444 0.424242424242 0 -0.4 1e-06 
1.0 0.424242424242 0 -0.4 1e-06 
0.5 0.464646464646 0 -0.4 1e-06 
0.555555555556 0.464646464646 0 -0.4 1e-06 
0.611111111111 0.464646464646 0 -0.4 1e-06 
0.666666666667 0.464646464646 0 -0.4 1e-06 
0.722222222222 0.464646464646 0 -0.4 1e-06 
0.777777777778 0.464646464646 0 -0.4 1e-06 
0.833333333333 0.464646464646 0 -0.4 1e-06 
0.888888888889 0.464646464646 0 -0.4 1e-06 
0.944444444444 0.464646464646 0 -0.4 1e-06 
1.0 0.464646464646 0 -0.4 1e-06 
0.5 0.505050505051 0 -0.4 1e-06 
0.555555555556 0.505050505051 0 -0.4 1e-06 
0.611111111111 0.505050505051 0 -0.4 1e-06 
0.666666666667 0.505050505051 0 -0.4 1e-06 
0.722222222222 0.505050505051 0 -0.4 1e-06 
0.777777777778 0.505050505051 0 -0.4 1e-06 
0.833333333333 0.505050505051 0 -0.4 1e-06 
0.888888888889 0.505050505051 0 -0.4 1e-06 
0.944444444444 0.505050505051 0 -0.4 1e-06 
1.0 0.505050505051 0 -0.4 1e-06 
0.5 0.545454545455 0 -0.4 1e-06 
0.555555555556 0.545454545455 0 -0.4 1e-06 
0.611111111111 0.545454545455 0 -0.4 1e-06 
0.666666666667 0.545454545455 0 -0.4 1e-06 
0.722222222222 0.545454545455 0 -0.4 1e-06 
0.777777777778 0.545454545455 0 -0.4 1e-06 
0.833333333333 0.545454545455 0 -0.4 1e-06 
0.888888888889 0.545454545455 0 -0.4 1e-06 
0.944444444444 0.545454545455 0 -0.4 1e-06 
1.0 0.545454545455 0 -0.4 1e-06 
0.5 0.585858585859 0 -0.4 1e-06 
0.555555555556 0.585858585859 0 -0.4 1e-06 
0.611111111111 0.585858585859 0 -0.4 1e-06 
0.666666666667 0.585858585859 0 -0.4 1e-06 
0.722222222222 0.585858585859 0 -0.4 1e-06 
0.777777777778 0.585858585859 0 -0.4 1e-06 
0.833333333333 0.585858585859 0 -0.4 1e-06 
0.888888888889 0.585858585859 0 -0.4 1e-06 
0.944444444444 0.585858585859 0 -0.4 1e-06 
1.0 0.585858585859 0 -0.4 1e-06 
0.5 0.626262626263 0 -0.4 1e-06 
0.555555555556 0.626262626263 0 -0.4 1e-06 
0.611111111111 0.626262626263 0 -0.4 1e-06 
0.666666666667 0.626262626263 0 -0.4 1e-06 
0.722222222222 0.626262626263 0 -0.4 1e-06 
0.777777777778 0.626262626263 0 -0.4 1e-06 
0.833333333333 0.626262626263 0 -0.4 1e-06 
0.888888888889 0.626262626263 0 -0.4 1e-06 
0.944444444444 0.626262626263 0 -0.4 1e-06 
1.0 0.626262626263 0 -0.4 1e-06 
0.5 0.666666666667 0 -0.4 1e-06 
0.555555555556 0.666666666667 0 -0.4 1e-06 
0.611111111111 0.666666666667 0 -0.4 1e-06 
0.666666666667 0.666666666667 0 -0.4 1e-06 
0.722222222222 0.666666666667 0 -0.4 1e-06 
0.777777777778 0.666666666667 0 -0.4 1e-06 
0.833333333333 0.666666666667 0 -0.4 1e-06 
0.888888888889 0.666666666667 0 -0.4 1e-06 
0.944444444444 0.666666666667 0 -0.4 1e-06 
1.0 0.666666666667 0 -0.4 1e-06 
0.5 0.707070707071 0 -0.4 1e-06 
0.555555555556 0.707070707071 0 -0.4 1e-06 
0.611111111111 0.707070707071 0 -0.4 1e-06 
0.666666666667 0.707070707071 0 -0.4 1e-06 
0.722222222222 0.707070707071 0 -0.4 1e-06 
0.777777777778 0.707070707071 0 -0.4 1e-06 
0.833333333333 0.707070707071 0 -0.4 1e-06 
0.888888888889 0.707070707071 0 -0.4 1e-06 
0.944444444444 0.707070707071 0 -0.4 1e-06 
1.0 0.707070707071 0 -0.4 1e-06 
0.5 0.747474747475 0 -0.4 1e-06 
0.555555555556 0.747474747475 0 -0.4 1e-06 
0.611111111111 0.747474747475 0 -0.4 1e-06 
0.666666666667 0.747474747475 0 -0.4 1e-06 
0.722222222222 0.747474747475 0 -0.4 1e-06 
0.777777777778 0.747474747475 0 -0.4 1e-06 
0.833333333333 0.747474747475 0 -0.4 1e-06 
0.888888888889 0.747474747475 0 -0.4 1e-06 
0.944444444444 0.747474747475 0 -0.4 1e-06 
1.0 0.747474747475 0 -0.4 1e-06 
0.5 0.787878787879 0 -0.4 1e-06 
0.555555555556 0.787878787879 0 -0.4 1e-06 
0.611111111111 0.787878787879 0 -0.4 1e-06 
0.666666666667 0.787878787879 0 -0.4 1e-06 
0.722222222222 0.787878787879 0 -0.4 1e-06 
0.777777777778 0.787878787879 0 -0.4 1e-06 
0.833333333333 0.787878787879 0 -0.4 1e-06 
0.888888888889 0.787878787879 0 -0.4 1e-06 
0.944444444444 0.787878787879 0 -0.4 1e-06 
1.0 0.787878787879 0 -0.4 1e-06 
0.5 0.828282828283 0 -0.4 1e-06 
0.555555555556 0.828282828283 0 -0.4 1e-06 
0.611111111111 0.828282828283 0 -0.4 1e-06 
0.666666666667 0.828282828283 0 -0.4 1e-06 
0.722222222222 0.828282828283 0 -0.4 1e-06 
0.777777777778 0.828282828283 0 -0.4 1e-06 
0.833333333333 0.828282828283 0 -0.4 1e-06 
0.888888888889 0.828282828283 0 -0.4 1e-06 
0.944444444444 0.828282828283 0 -0.4 1e-06 
1.0 0.828282828283 0 -0.4 1e-06 
0.5 0.868686868687 0 -0.4 1e-06 
0.555555555556 0.868686868687 0 -0.4 1e-06 
0.611111111111 0.868686868687 0 -0.4 1e-06 
0.666666666667 0.868686868687 0 -0.4 1e-06 
0.722222222222 0.868686868687 0 -0.4 1e-06 
0.777777777778 0.868686868687 0 -0.4 1e-06 
0.833333333333 0.868686868687 0 -0.4 1e-06 
0.888888888889 0.868686868687 0 -0.4 1e-06 
0.944444444444 0.868686868687 0 -0.4 1e-06 
1.0 0.868686868687 0 -0.4 1e-06 
0.5 0.909090909091 0 -0.4 1e-06 
0.555555555556 0.909090909091 0 -0.4 1e-06 
0.611111111111 0.909090909091 0 -0.4 1e-06 
0.666666666667 0.909090909091 0 -0.4 1e-06 
0.722222222222 0.909090909091 0 -0.4 1e-06 
0.777777777778 0.909090909091 0 -0.4 1e-06 
0.833333333333 0.909090909091 0 -0.4 1e-06 
0.888888888889 0.909090909091 0 -0.4 1e-06 
0.944444444444 0.909090909091 0 -0.4 1e-06 
1.0 0.909090909091 0 -0.4 1e-06 
0.5 0.949494949495 0 -0.4 1e-06 
0.555555555556 0.949494949495 0 -0.4 1e-06 
0.611111111111 0.949494949495 0 -0.4 1e-06 
0.666666666667 0.949494949495 0 -0.4 1e-06 
0.722222222222 0.949494949495 0 -0.4 1e-06 
0.777777777778 0.949494949495 0 -0.4 1e-06 
0.833333333333 0.949494949495 0 -0.4 1e-06 
0.888888888889 0.949494949495 0 -0.4 1e-06 
0.944444444444 0.949494949495 0 -0.4 1e-06 
1.0 0.949494949495 0 -0.4 1e-06 
0.5 0.989898989899 0 -0.4 1e-06 
0.555555555556 0.989898989899 0 -0.4 1e-06 
0.611111111111 0.989898989899 0 -0.4 1e-06 
0.666666666667 0.989898989899 0 -0.4 1e-06 
0.722222222222 0.989898989899 0 -0.4 1e-06 
0.777777777778 0.989898989899 0 -0.4 1e-06 
0.833333333333 0.989898989899 0 -0.4 1e-06 
0.888888888889 0.989898989899 0 -0.4 1e-06 
0.944444444444 0.989898989899 0 -0.4 1e-06 
1.0 0.989898989899 0 -0.4 1e-06 
0.5 1.0303030303 0 -0.4 1e-06 
0.555555555556 1.0303030303 0 -0.4 1e-06 
0.611111111111 1.0303030303 0 -0.4 1e-06 
0.666666666667 1.0303030303 0 -0.4 1e-06 
0.722222222222 1.0303030303 0 -0.4 1e-06 
0.777777777778 1.0303030303 0 -0.4 1e-06 
0.833333333333 1.0303030303 0 -0.4 1e-06 
0.888888888889 1.0303030303 0 -0.4 1e-06 
0.944444444444 1.0303030303 0 -0.4 1e-06 
1.0 1.0303030303 0 -0.4 1e-06 
0.5 1.07070707071 0 -0.4 1e-06 
0.555555555556 1.07070707071 0 -0.4 1e-06 
0.611111111111 1.07070707071 0 -0.4 1e-06 
0.666666666667 1.07070707071 0 -0.4 1e-06 
0.722222222222 1.07070707071 0 -0.4 1e-06 
0.777777777778 1.07070707071 0 -0.4 1e-06 
0.833333333333 1.07070707071 0 -0.4 1e-06 
0.888888888889 1.07070707071 0 -0.4 1e-06 
0.944444444444 1.07070707071 0 -0.4 1e-06 
1.0 1.07070707071 0 -0.4 1e-06 
0.5 1.11111111111 0 -0.4 1e-06 
0.555555555556 1.11111111111 0 -0.4 1e-06 
0.611111111111 1.11111111111 0 -0.4 1e-06 
0.666666666667 1.11111111111 0 -0.4 1e-06 
0.722222222222 1.11111111111 0 -0.4 1e-06 
0.777777777778 1.11111111111 0 -0.4 1e-06 
0.833333333333 1.11111111111 0 -0.4 1e-06 
0.888888888889 1.11111111111 0 -0.4 1e-06 
0.944444444444 1.11111111111 0 -0.4 1e-06 
1.0 1.11111111111 0 -0.4 1e-06 
0.5 1.15151515152 0 -0.4 1e-06 
0.555555555556 1.15151515152 0 -0.4 1e-06 
0.611111111111 1.15151515152 0 -0.4 1e-06 
0.666666666667 1.15151515152 0 -0.4 1e-06 
0.722222222222 1.15151515152 0 -0.4 1e-06 
0.777777777778 1.15151515152 0 -0.4 1e-06 
0.833333333333 1.15151515152 0 -0.4 1e-06 
0.888888888889 1.15151515152 0 -0.4 1e-06 
0.944444444444 1.15151515152 0 -0.4 1e-06 
1.0 1.15151515152 0 -0.4 1e-06 
0.5 1.19191919192 0 -0.4 1e-06 
0.555555555556 1.19191919192 0 -0.4 1e-06 
0.611111111111 1.19191919192 0 -0.4 1e-06 
0.666666666667 1.19191919192 0 -0.4 1e-06 
0.722222222222 1.19191919192 0 -0.4 1e-06 
0.777777777778 1.19191919192 0 -0.4 1e-06 
0.833333333333 1.19191919192 0 -0.4 1e-06 
0.888888888889 1.19191919192 0 -0.4 1e-06 
0.944444444444 1.19191919192 0 -0.4 1e-06 
1.0 1.19191919192 0 -0.4 1e-06 
0.5 1.23232323232 0 -0.4 1e-06 
0.555555555556 1.23232323232 0 -0.4 1e-06 
0.611111111111 1.23232323232 0 -0.4 1e-06 
0.666666666667 1.23232323232 0 -0.4 1e-06 
0.722222222222 1.23232323232 0 -0.4 1e-06 
0.777777777778 1.23232323232 0 -0.4 1e-06 
0.833333333333 1.23232323232 0 -0.4 1e-06 
0.888888888889 1.23232323232 0 -0.4 1e-06 
0.944444444444 1.23232323232 0 -0.4 1e-06 
1.0 1.23232323232 0 -0.4 1e-06 
0.5 1.27272727273 0 -0.4 1e-06 
0.555555555556 1.27272727273 0 -0.4 1e-06 
0.611111111111 1.27272727273 0 -0.4 1e-06 
0.666666666667 1.27272727273 0 -0.4 1e-06 
0.722222222222 1.27272727273 0 -0.4 1e-06 
0.777777777778 1.27272727273 0 -0.4 1e-06 
0.833333333333 1.27272727273 0 -0.4 1e-06 
0.888888888889 1.27272727273 0 -0.4 1e-06 
0.944444444444 1.27272727273 0 -0.4 1e-06 
1.0 1.27272727273 0 -0.4 1e-06 
0.5 1.31313131313 0 -0.4 1e-06 
0.555555555556 1.31313131313 0 -0.4 1e-06 
0.611111111111 1.31313131313 0 -0.4 1e-06 
0.666666666667 1.31313131313 0 -0.4 1e-06 
0.722222222222 1.31313131313 0 -0.4 1e-06 
0.777777777778 1.31313131313 0 -0.4 1e-06 
0.833333333333 1.31313131313 0 -0.4 1e-06 
0.888888888889 1.31313131313 0 -0.4 1e-06 
0.944444444444 1.31313131313 0 -0.4 1e-06 
1.0 1.31313131313 0 -0.4 1e-06 
0.5 1.35353535354 0 -0.4 1e-06 
0.555555555556 1.35353535354 0 -0.4 1e-06 
0.611111111111 1.35353535354 0 -0.4 1e-06 
0.666666666667 1.35353535354 0 -0.4 1e-06 
0.722222222222 1.35353535354 0 -0.4 1e-06 
0.777777777778 1.35353535354 0 -0.4 1e-06 
0.833333333333 1.35353535354 0 -0.4 1e-06 
0.888888888889 1.35353535354 0 -0.4 1e-06 
0.944444444444 1.35353535354 0 -0.4 1e-06 
1.0 1.35353535354 0 -0.4 1e-06 
0.5 1.39393939394 0 -0.4 1e-06 
0.555555555556 1.39393939394 0 -0.4 1e-06 
0.611111111111 1.39393939394 0 -0.4 1e-06 
0.666666666667 1.39393939394 0 -0.4 1e-06 
0.722222222222 1.39393939394 0 -0.4 1e-06 
0.777777777778 1.39393939394 0 -0.4 1e-06 
0.833333333333 1.39393939394 0 -0.4 1e-06 
0.888888888889 1.39393939394 0 -0.4 1e-06 
0.944444444444 1.39393939394 0 -0.4 1e-06 
1.0 1.39393939394 0 -0.4 1e-06 
0.5 1.43434343434 0 -0.4 1e-06 
0.555555555556 1.43434343434 0 -0.4 1e-06 
0.611111111111 1.43434343434 0 -0.4 1e-06 
0.666666666667 1.43434343434 0 -0.4 1e-06 
0.722222222222 1.43434343434 0 -0.4 1e-06 
0.777777777778 1.43434343434 0 -0.4 1e-06 
0.833333333333 1.43434343434 0 -0.4 1e-06 
0.888888888889 1.43434343434 0 -0.4 1e-06 
0.944444444444 1.43434343434 0 -0.4 1e-06 
1.0 1.43434343434 0 -0.4 1e-06 
0.5 1.47474747475 0 -0.4 1e-06 
0.555555555556 1.47474747475 0 -0.4 1e-06 
0.611111111111 1.47474747475 0 -0.4 1e-06 
0.666666666667 1.47474747475 0 -0.4 1e-06 
0.722222222222 1.47474747475 0 -0.4 1e-06 
0.777777777778 1.47474747475 0 -0.4 1e-06 
0.833333333333 1.47474747475 0 -0.4 1e-06 
0.888888888889 1.47474747475 0 -0.4 1e-06 
0.944444444444 1.47474747475 0 -0.4 1e-06 
1.0 1.47474747475 0 -0.4 1e-06 
0.5 1.51515151515 0 -0.4 1e-06 
0.555555555556 1.51515151515 0 -0.4 1e-06 
0.611111111111 1.51515151515 0 -0.4 1e-06 
0.666666666667 1.51515151515 0 -0.4 1e-06 
0.722222222222 1.51515151515 0 -0.4 1e-06 
0.777777777778 1.51515151515 0 -0.4 1e-06 
0.833333333333 1.51515151515 0 -0.4 1e-06 
0.888888888889 1.51515151515 0 -0.4 1e-06 
0.944444444444 1.51515151515 0 -0.4 1e-06 
1.0 1.51515151515 0 -0.4 1e-06 
0.5 1.55555555556 0 -0.4 1e-06 
0.555555555556 1.55555555556 0 -0.4 1e-06 
0.611111111111 1.55555555556 0 -0.4 1e-06 
0.666666666667 1.55555555556 0 -0.4 1e-06 
0.722222222222 1.55555555556 0 -0.4 1e-06 
0.777777777778 1.55555555556 0 -0.4 1e-06 
0.833333333333 1.55555555556 0 -0.4 1e-06 
0.888888888889 1.55555555556 0 -0.4 1e-06 
0.944444444444 1.55555555556 0 -0.4 1e-06 
1.0 1.55555555556 0 -0.4 1e-06 
0.5 1.59595959596 0 -0.4 1e-06 
0.555555555556 1.59595959596 0 -0.4 1e-06 
0.611111111111 1.59595959596 0 -0.4 1e-06 
0.666666666667 1.59595959596 0 -0.4 1e-06 
0.722222222222 1.59595959596 0 -0.4 1e-06 
0.777777777778 1.59595959596 0 -0.4 1e-06 
0.833333333333 1.59595959596 0 -0.4 1e-06 
0.888888888889 1.59595959596 0 -0.4 1e-06 
0.944444444444 1.59595959596 0 -0.4 1e-06 
1.0 1.59595959596 0 -0.4 1e-06 
0.5 1.63636363636 0 -0.4 1e-06 
0.555555555556 1.63636363636 0 -0.4 1e-06 
0.611111111111 1.63636363636 0 -0.4 1e-06 
0.666666666667 1.63636363636 0 -0.4 1e-06 
0.722222222222 1.63636363636 0 -0.4 1e-06 
0.777777777778 1.63636363636 0 -0.4 1e-06 
0.833333333333 1.63636363636 0 -0.4 1e-06 
0.888888888889 1.63636363636 0 -0.4 1e-06 
0.944444444444 1.63636363636 0 -0.4 1e-06 
1.0 1.63636363636 0 -0.4 1e-06 
0.5 1.67676767677 0 -0.4 1e-06 
0.555555555556 1.67676767677 0 -0.4 1e-06 
0.611111111111 1.67676767677 0 -0.4 1e-06 
0.666666666667 1.67676767677 0 -0.4 1e-06 
0.722222222222 1.67676767677 0 -0.4 1e-06 
0.777777777778 1.67676767677 0 -0.4 1e-06 
0.833333333333 1.67676767677 0 -0.4 1e-06 
0.888888888889 1.67676767677 0 -0.4 1e-06 
0.944444444444 1.67676767677 0 -0.4 1e-06 
1.0 1.67676767677 0 -0.4 1e-06 
0.5 1.71717171717 0 -0.4 1e-06 
0.555555555556 1.71717171717 0 -0.4 1e-06 
0.611111111111 1.71717171717 0 -0.4 1e-06 
0.666666666667 1.71717171717 0 -0.4 1e-06 
0.722222222222 1.71717171717 0 -0.4 1e-06 
0.777777777778 1.71717171717 0 -0.4 1e-06 
0.833333333333 1.71717171717 0 -0.4 1e-06 
0.888888888889 1.71717171717 0 -0.4 1e-06 
0.944444444444 1.71717171717 0 -0.4 1e-06 
1.0 1.71717171717 0 -0.4 1e-06 
0.5 1.75757575758 0 -0.4 1e-06 
0.555555555556 1.75757575758 0 -0.4 1e-06 
0.611111111111 1.75757575758 0 -0.4 1e-06 
0.666666666667 1.75757575758 0 -0.4 1e-06 
0.722222222222 1.75757575758 0 -0.4 1e-06 
0.777777777778 1.75757575758 0 -0.4 1e-06 
0.833333333333 1.75757575758 0 -0.4 1e-06 
0.888888888889 1.75757575758 0 -0.4 1e-06 
0.944444444444 1.75757575758 0 -0.4 1e-06 
1.0 1.75757575758 0 -0.4 1e-06 
0.5 1.79797979798 0 -0.4 1e-06 
0.555555555556 1.79797979798 0 -0.4 1e-06 
0.611111111111 1.79797979798 0 -0.4 1e-06 
0.666666666667 1.79797979798 0 -0.4 1e-06 
0.722222222222 1.79797979798 0 -0.4 1e-06 
0.777777777778 1.79797979798 0 -0.4 1e-06 
0.833333333333 1.79797979798 0 -0.4 1e-06 
0.888888888889 1.79797979798 0 -0.4 1e-06 
0.944444444444 1.79797979798 0 -0.4 1e-06 
1.0 1.79797979798 0 -0.4 1e-06 
0.5 1.83838383838 0 -0.4 1e-06 
0.555555555556 1.83838383838 0 -0.4 1e-06 
0.611111111111 1.83838383838 0 -0.4 1e-06 
0.666666666667 1.83838383838 0 -0.4 1e-06 
0.722222222222 1.83838383838 0 -0.4 1e-06 
0.777777777778 1.83838383838 0 -0.4 1e-06 
0.833333333333 1.83838383838 0 -0.4 1e-06 
0.888888888889 1.83838383838 0 -0.4 1e-06 
0.944444444444 1.83838383838 0 -0.4 1e-06 
1.0 1.83838383838 0 -0.4 1e-06 
0.5 1.87878787879 0 -0.4 1e-06 
0.555555555556 1.87878787879 0 -0.4 1e-06 
0.611111111111 1.87878787879 0 -0.4 1e-06 
0.666666666667 1.87878787879 0 -0.4 1e-06 
0.722222222222 1.87878787879 0 -0.4 1e-06 
0.777777777778 1.87878787879 0 -0.4 1e-06 
0.833333333333 1.87878787879 0 -0.4 1e-06 
0.888888888889 1.87878787879 0 -0.4 1e-06 
0.944444444444 1.87878787879 0 -0.4 1e-06 
1.0 1.87878787879 0 -0.4 1e-06 
0.5 1.91919191919 0 -0.4 1e-06 
0.555555555556 1.91919191919 0 -0.4 1e-06 
0.611111111111 1.91919191919 0 -0.4 1e-06 
0.666666666667 1.91919191919 0 -0.4 1e-06 
0.722222222222 1.91919191919 0 -0.4 1e-06 
0.777777777778 1.91919191919 0 -0.4 1e-06 
0.833333333333 1.91919191919 0 -0.4 1e-06 
0.888888888889 1.91919191919 0 -0.4 1e-06 
0.944444444444 1.91919191919 0 -0.4 1e-06 
1.0 1.91919191919 0 -0.4 1e-06 
0.5 1.9595959596 0 -0.4 1e-06 
0.555555555556 1.9595959596 0 -0.4 1e-06 
0.611111111111 1.9595959596 0 -0.4 1e-06 
0.666666666667 1.9595959596 0 -0.4 1e-06 
0.722222222222 1.9595959596 0 -0.4 1e-06 
0.777777777778 1.9595959596 0 -0.4 1e-06 
0.833333333333 1.9595959596 0 -0.4 1e-06 
0.888888888889 1.9595959596 0 -0.4 1e-06 
0.944444444444 1.9595959596 0 -0.4 1e-06 
1.0 1.9595959596 0 -0.4 1e-06 
0.5 2.0 0 -0.4 1e-06 
0.555555555556 2.0 0 -0.4 1e-06 
0.611111111111 2.0 0 -0.4 1e-06 
0.666666666667 2.0 0 -0.4 1e-06 
0.722222222222 2.0 0 -0.4 1e-06 
0.777777777778 2.0 0 -0.4 1e-06 
0.833333333333 2.0 0 -0.4 1e-06 
0.888888888889 2.0 0 -0.4 1e-06 
0.944444444444 2.0 0 -0.4 1e-06 
1.0 2.0 0 -0.4 1e-06 
0.5 -2.0 0 0.0 1e-06 
0.555555555556 -2.0 0 0.0 1e-06 
0.611111111111 -2.0 0 0.0 1e-06 
0.666666666667 -2.0 0 0.0 1e-06 
0.722222222222 -2.0 0 0.0 1e-06 
0.777777777778 -2.0 0 0.0 1e-06 
0.833333333333 -2.0 0 0.0 1e-06 
0.888888888889 -2.0 0 0.0 1e-06 
0.944444444444 -2.0 0 0.0 1e-06 
1.0 -2.0 0 0.0 1e-06 
0.5 -1.9595959596 0 0.0 1e-06 
0.555555555556 -1.9595959596 0 0.0 1e-06 
0.611111111111 -1.9595959596 0 0.0 1e-06 
0.666666666667 -1.9595959596 0 0.0 1e-06 
0.722222222222 -1.9595959596 0 0.0 1e-06 
0.777777777778 -1.9595959596 0 0.0 1e-06 
0.833333333333 -1.9595959596 0 0.0 1e-06 
0.888888888889 -1.9595959596 0 0.0 1e-06 
0.944444444444 -1.9595959596 0 0.0 1e-06 
1.0 -1.9595959596 0 0.0 1e-06 
0.5 -1.91919191919 0 0.0 1e-06 
0.555555555556 -1.91919191919 0 0.0 1e-06 
0.611111111111 -1.91919191919 0 0.0 1e-06 
0.666666666667 -1.91919191919 0 0.0 1e-06 
0.722222222222 -1.91919191919 0 0.0 1e-06 
0.777777777778 -1.91919191919 0 0.0 1e-06 
0.833333333333 -1.91919191919 0 0.0 1e-06 
0.888888888889 -1.91919191919 0 0.0 1e-06 
0.944444444444 -1.91919191919 0 0.0 1e-06 
1.0 -1.91919191919 0 0.0 1e-06 
0.5 -1.87878787879 0 0.0 1e-06 
0.555555555556 -1.87878787879 0 0.0 1e-06 
0.611111111111 -1.87878787879 0 0.0 1e-06 
0.666666666667 -1.87878787879 0 0.0 1e-06 
0.722222222222 -1.87878787879 0 0.0 1e-06 
0.777777777778 -1.87878787879 0 0.0 1e-06 
0.833333333333 -1.87878787879 0 0.0 1e-06 
0.888888888889 -1.87878787879 0 0.0 1e-06 
0.944444444444 -1.87878787879 0 0.0 1e-06 
1.0 -1.87878787879 0 0.0 1e-06 
0.5 -1.83838383838 0 0.0 1e-06 
0.555555555556 -1.83838383838 0 0.0 1e-06 
0.611111111111 -1.83838383838 0 0.0 1e-06 
0.666666666667 -1.83838383838 0 0.0 1e-06 
0.722222222222 -1.83838383838 0 0.0 1e-06 
0.777777777778 -1.83838383838 0 0.0 1e-06 
0.833333333333 -1.83838383838 0 0.0 1e-06 
0.888888888889 -1.83838383838 0 0.0 1e-06 
0.944444444444 -1.83838383838 0 0.0 1e-06 
1.0 -1.83838383838 0 0.0 1e-06 
0.5 -1.79797979798 0 0.0 1e-06 
0.555555555556 -1.79797979798 0 0.0 1e-06 
0.611111111111 -1.79797979798 0 0.0 1e-06 
0.666666666667 -1.79797979798 0 0.0 1e-06 
0.722222222222 -1.79797979798 0 0.0 1e-06 
0.777777777778 -1.79797979798 0 0.0 1e-06 
0.833333333333 -1.79797979798 0 0.0 1e-06 
0.888888888889 -1.79797979798 0 0.0 1e-06 
0.944444444444 -1.79797979798 0 0.0 1e-06 
1.0 -1.79797979798 0 0.0 1e-06 
0.5 -1.75757575758 0 0.0 1e-06 
0.555555555556 -1.75757575758 0 0.0 1e-06 
0.611111111111 -1.75757575758 0 0.0 1e-06 
0.666666666667 -1.75757575758 0 0.0 1e-06 
0.722222222222 -1.75757575758 0 0.0 1e-06 
0.777777777778 -1.75757575758 0 0.0 1e-06 
0.833333333333 -1.75757575758 0 0.0 1e-06 
0.888888888889 -1.75757575758 0 0.0 1e-06 
0.944444444444 -1.75757575758 0 0.0 1e-06 
1.0 -1.75757575758 0 0.0 1e-06 
0.5 -1.71717171717 0 0.0 1e-06 
0.555555555556 -1.71717171717 0 0.0 1e-06 
0.611111111111 -1.71717171717 0 0.0 1e-06 
0.666666666667 -1.71717171717 0 0.0 1e-06 
0.722222222222 -1.71717171717 0 0.0 1e-06 
0.777777777778 -1.71717171717 0 0.0 1e-06 
0.833333333333 -1.71717171717 0 0.0 1e-06 
0.888888888889 -1.71717171717 0 0.0 1e-06 
0.944444444444 -1.71717171717 0 0.0 1e-06 
1.0 -1.71717171717 0 0.0 1e-06 
0.5 -1.67676767677 0 0.0 1e-06 
0.555555555556 -1.67676767677 0 0.0 1e-06 
0.611111111111 -1.67676767677 0 0.0 1e-06 
0.666666666667 -1.67676767677 0 0.0 1e-06 
0.722222222222 -1.67676767677 0 0.0 1e-06 
0.777777777778 -1.67676767677 0 0.0 1e-06 
0.833333333333 -1.67676767677 0 0.0 1e-06 
0.888888888889 -1.67676767677 0 0.0 1e-06 
0.944444444444 -1.67676767677 0 0.0 1e-06 
1.0 -1.67676767677 0 0.0 1e-06 
0.5 -1.63636363636 0 0.0 1e-06 
0.555555555556 -1.63636363636 0 0.0 1e-06 
0.611111111111 -1.63636363636 0 0.0 1e-06 
0.666666666667 -1.63636363636 0 0.0 1e-06 
0.722222222222 -1.63636363636 0 0.0 1e-06 
0.777777777778 -1.63636363636 0 0.0 1e-06 
0.833333333333 -1.63636363636 0 0.0 1e-06 
0.888888888889 -1.63636363636 0 0.0 1e-06 
0.944444444444 -1.63636363636 0 0.0 1e-06 
1.0 -1.63636363636 0 0.0 1e-06 
0.5 -1.59595959596 0 0.0 1e-06 
0.555555555556 -1.59595959596 0 0.0 1e-06 
0.611111111111 -1.59595959596 0 0.0 1e-06 
0.666666666667 -1.59595959596 0 0.0 1e-06 
0.722222222222 -1.59595959596 0 0.0 1e-06 
0.777777777778 -1.59595959596 0 0.0 1e-06 
0.833333333333 -1.59595959596 0 0.0 1e-06 
0.888888888889 -1.59595959596 0 0.0 1e-06 
0.944444444444 -1.59595959596 0 0.0 1e-06 
1.0 -1.59595959596 0 0.0 1e-06 
0.5 -1.55555555556 0 0.0 1e-06 
0.555555555556 -1.55555555556 0 0.0 1e-06 
0.611111111111 -1.55555555556 0 0.0 1e-06 
0.666666666667 -1.55555555556 0 0.0 1e-06 
0.722222222222 -1.55555555556 0 0.0 1e-06 
0.777777777778 -1.55555555556 0 0.0 1e-06 
0.833333333333 -1.55555555556 0 0.0 1e-06 
0.888888888889 -1.55555555556 0 0.0 1e-06 
0.944444444444 -1.55555555556 0 0.0 1e-06 
1.0 -1.55555555556 0 0.0 1e-06 
0.5 -1.51515151515 0 0.0 1e-06 
0.555555555556 -1.51515151515 0 0.0 1e-06 
0.611111111111 -1.51515151515 0 0.0 1e-06 
0.666666666667 -1.51515151515 0 0.0 1e-06 
0.722222222222 -1.51515151515 0 0.0 1e-06 
0.777777777778 -1.51515151515 0 0.0 1e-06 
0.833333333333 -1.51515151515 0 0.0 1e-06 
0.888888888889 -1.51515151515 0 0.0 1e-06 
0.944444444444 -1.51515151515 0 0.0 1e-06 
1.0 -1.51515151515 0 0.0 1e-06 
0.5 -1.47474747475 0 0.0 1e-06 
0.555555555556 -1.47474747475 0 0.0 1e-06 
0.611111111111 -1.47474747475 0 0.0 1e-06 
0.666666666667 -1.47474747475 0 0.0 1e-06 
0.722222222222 -1.47474747475 0 0.0 1e-06 
0.777777777778 -1.47474747475 0 0.0 1e-06 
0.833333333333 -1.47474747475 0 0.0 1e-06 
0.888888888889 -1.47474747475 0 0.0 1e-06 
0.944444444444 -1.47474747475 0 0.0 1e-06 
1.0 -1.47474747475 0 0.0 1e-06 
0.5 -1.43434343434 0 0.0 1e-06 
0.555555555556 -1.43434343434 0 0.0 1e-06 
0.611111111111 -1.43434343434 0 0.0 1e-06 
0.666666666667 -1.43434343434 0 0.0 1e-06 
0.722222222222 -1.43434343434 0 0.0 1e-06 
0.777777777778 -1.43434343434 0 0.0 1e-06 
0.833333333333 -1.43434343434 0 0.0 1e-06 
0.888888888889 -1.43434343434 0 0.0 1e-06 
0.944444444444 -1.43434343434 0 0.0 1e-06 
1.0 -1.43434343434 0 0.0 1e-06 
0.5 -1.39393939394 0 0.0 1e-06 
0.555555555556 -1.39393939394 0 0.0 1e-06 
0.611111111111 -1.39393939394 0 0.0 1e-06 
0.666666666667 -1.39393939394 0 0.0 1e-06 
0.722222222222 -1.39393939394 0 0.0 1e-06 
0.777777777778 -1.39393939394 0 0.0 1e-06 
0.833333333333 -1.39393939394 0 0.0 1e-06 
0.888888888889 -1.39393939394 0 0.0 1e-06 
0.944444444444 -1.39393939394 0 0.0 1e-06 
1.0 -1.39393939394 0 0.0 1e-06 
0.5 -1.35353535354 0 0.0 1e-06 
0.555555555556 -1.35353535354 0 0.0 1e-06 
0.611111111111 -1.35353535354 0 0.0 1e-06 
0.666666666667 -1.35353535354 0 0.0 1e-06 
0.722222222222 -1.35353535354 0 0.0 1e-06 
0.777777777778 -1.35353535354 0 0.0 1e-06 
0.833333333333 -1.35353535354 0 0.0 1e-06 
0.888888888889 -1.35353535354 0 0.0 1e-06 
0.944444444444 -1.35353535354 0 0.0 1e-06 
1.0 -1.35353535354 0 0.0 1e-06 
0.5 -1.31313131313 0 0.0 1e-06 
0.555555555556 -1.31313131313 0 0.0 1e-06 
0.611111111111 -1.31313131313 0 0.0 1e-06 
0.666666666667 -1.31313131313 0 0.0 1e-06 
0.722222222222 -1.31313131313 0 0.0 1e-06 
0.777777777778 -1.31313131313 0 0.0 1e-06 
0.833333333333 -1.31313131313 0 0.0 1e-06 
0.888888888889 -1.31313131313 0 0.0 1e-06 
0.944444444444 -1.31313131313 0 0.0 1e-06 
1.0 -1.31313131313 0 0.0 1e-06 
0.5 -1.27272727273 0 0.0 1e-06 
0.555555555556 -1.27272727273 0 0.0 1e-06 
0.611111111111 -1.27272727273 0 0.0 1e-06 
0.666666666667 -1.27272727273 0 0.0 1e-06 
0.722222222222 -1.27272727273 0 0.0 1e-06 
0.777777777778 -1.27272727273 0 0.0 1e-06 
0.833333333333 -1.27272727273 0 0.0 1e-06 
0.888888888889 -1.27272727273 0 0.0 1e-06 
0.944444444444 -1.27272727273 0 0.0 1e-06 
1.0 -1.27272727273 0 0.0 1e-06 
0.5 -1.23232323232 0 0.0 1e-06 
0.555555555556 -1.23232323232 0 0.0 1e-06 
0.611111111111 -1.23232323232 0 0.0 1e-06 
0.666666666667 -1.23232323232 0 0.0 1e-06 
0.722222222222 -1.23232323232 0 0.0 1e-06 
0.777777777778 -1.23232323232 0 0.0 1e-06 
0.833333333333 -1.23232323232 0 0.0 1e-06 
0.888888888889 -1.23232323232 0 0.0 1e-06 
0.944444444444 -1.23232323232 0 0.0 1e-06 
1.0 -1.23232323232 0 0.0 1e-06 
0.5 -1.19191919192 0 0.0 1e-06 
0.555555555556 -1.19191919192 0 0.0 1e-06 
0.611111111111 -1.19191919192 0 0.0 1e-06 
0.666666666667 -1.19191919192 0 0.0 1e-06 
0.722222222222 -1.19191919192 0 0.0 1e-06 
0.777777777778 -1.19191919192 0 0.0 1e-06 
0.833333333333 -1.19191919192 0 0.0 1e-06 
0.888888888889 -1.19191919192 0 0.0 1e-06 
0.944444444444 -1.19191919192 0 0.0 1e-06 
1.0 -1.19191919192 0 0.0 1e-06 
0.5 -1.15151515152 0 0.0 1e-06 
0.555555555556 -1.15151515152 0 0.0 1e-06 
0.611111111111 -1.15151515152 0 0.0 1e-06 
0.666666666667 -1.15151515152 0 0.0 1e-06 
0.722222222222 -1.15151515152 0 0.0 1e-06 
0.777777777778 -1.15151515152 0 0.0 1e-06 
0.833333333333 -1.15151515152 0 0.0 1e-06 
0.888888888889 -1.15151515152 0 0.0 1e-06 
0.944444444444 -1.15151515152 0 0.0 1e-06 
1.0 -1.15151515152 0 0.0 1e-06 
0.5 -1.11111111111 0 0.0 1e-06 
0.555555555556 -1.11111111111 0 0.0 1e-06 
0.611111111111 -1.11111111111 0 0.0 1e-06 
0.666666666667 -1.11111111111 0 0.0 1e-06 
0.722222222222 -1.11111111111 0 0.0 1e-06 
0.777777777778 -1.11111111111 0 0.0 1e-06 
0.833333333333 -1.11111111111 0 0.0 1e-06 
0.888888888889 -1.11111111111 0 0.0 1e-06 
0.944444444444 -1.11111111111 0 0.0 1e-06 
1.0 -1.11111111111 0 0.0 1e-06 
0.5 -1.07070707071 0 0.0 1e-06 
0.555555555556 -1.07070707071 0 0.0 1e-06 
0.611111111111 -1.07070707071 0 0.0 1e-06 
0.666666666667 -1.07070707071 0 0.0 1e-06 
0.722222222222 -1.07070707071 0 0.0 1e-06 
0.777777777778 -1.07070707071 0 0.0 1e-06 
0.833333333333 -1.07070707071 0 0.0 1e-06 
0.888888888889 -1.07070707071 0 0.0 1e-06 
0.944444444444 -1.07070707071 0 0.0 1e-06 
1.0 -1.07070707071 0 0.0 1e-06 
0.5 -1.0303030303 0 0.0 1e-06 
0.555555555556 -1.0303030303 0 0.0 1e-06 
0.611111111111 -1.0303030303 0 0.0 1e-06 
0.666666666667 -1.0303030303 0 0.0 1e-06 
0.722222222222 -1.0303030303 0 0.0 1e-06 
0.777777777778 -1.0303030303 0 0.0 1e-06 
0.833333333333 -1.0303030303 0 0.0 1e-06 
0.888888888889 -1.0303030303 0 0.0 1e-06 
0.944444444444 -1.0303030303 0 0.0 1e-06 
1.0 -1.0303030303 0 0.0 1e-06 
0.5 -0.989898989899 0 0.0 1e-06 
0.555555555556 -0.989898989899 0 0.0 1e-06 
0.611111111111 -0.989898989899 0 0.0 1e-06 
0.666666666667 -0.989898989899 0 0.0 1e-06 
0.722222222222 -0.989898989899 0 0.0 1e-06 
0.777777777778 -0.989898989899 0 0.0 1e-06 
0.833333333333 -0.989898989899 0 0.0 1e-06 
0.888888888889 -0.989898989899 0 0.0 1e-06 
0.944444444444 -0.989898989899 0 0.0 1e-06 
1.0 -0.989898989899 0 0.0 1e-06 
0.5 -0.949494949495 0 0.0 1e-06 
0.555555555556 -0.949494949495 0 0.0 1e-06 
0.611111111111 -0.949494949495 0 0.0 1e-06 
0.666666666667 -0.949494949495 0 0.0 1e-06 
0.722222222222 -0.949494949495 0 0.0 1e-06 
0.777777777778 -0.949494949495 0 0.0 1e-06 
0.833333333333 -0.949494949495 0 0.0 1e-06 
0.888888888889 -0.949494949495 0 0.0 1e-06 
0.944444444444 -0.949494949495 0 0.0 1e-06 
1.0 -0.949494949495 0 0.0 1e-06 
0.5 -0.909090909091 0 0.0 1e-06 
0.555555555556 -0.909090909091 0 0.0 1e-06 
0.611111111111 -0.909090909091 0 0.0 1e-06 
0.666666666667 -0.909090909091 0 0.0 1e-06 
0.722222222222 -0.909090909091 0 0.0 1e-06 
0.777777777778 -0.909090909091 0 0.0 1e-06 
0.833333333333 -0.909090909091 0 0.0 1e-06 
0.888888888889 -0.909090909091 0 0.0 1e-06 
0.944444444444 -0.909090909091 0 0.0 1e-06 
1.0 -0.909090909091 0 0.0 1e-06 
0.5 -0.868686868687 0 0.0 1e-06 
0.555555555556 -0.868686868687 0 0.0 1e-06 
0.611111111111 -0.868686868687 0 0.0 1e-06 
0.666666666667 -0.868686868687 0 0.0 1e-06 
0.722222222222 -0.868686868687 0 0.0 1e-06 
0.777777777778 -0.868686868687 0 0.0 1e-06 
0.833333333333 -0.868686868687 0 0.0 1e-06 
0.888888888889 -0.868686868687 0 0.0 1e-06 
0.944444444444 -0.868686868687 0 0.0 1e-06 
1.0 -0.868686868687 0 0.0 1e-06 
0.5 -0.828282828283 0 0.0 1e-06 
0.555555555556 -0.828282828283 0 0.0 1e-06 
0.611111111111 -0.828282828283 0 0.0 1e-06 
0.666666666667 -0.828282828283 0 0.0 1e-06 
0.722222222222 -0.828282828283 0 0.0 1e-06 
0.777777777778 -0.828282828283 0 0.0 1e-06 
0.833333333333 -0.828282828283 0 0.0 1e-06 
0.888888888889 -0.828282828283 0 0.0 1e-06 
0.944444444444 -0.828282828283 0 0.0 1e-06 
1.0 -0.828282828283 0 0.0 1e-06 
0.5 -0.787878787879 0 0.0 1e-06 
0.555555555556 -0.787878787879 0 0.0 1e-06 
0.611111111111 -0.787878787879 0 0.0 1e-06 
0.666666666667 -0.787878787879 0 0.0 1e-06 
0.722222222222 -0.787878787879 0 0.0 1e-06 
0.777777777778 -0.787878787879 0 0.0 1e-06 
0.833333333333 -0.787878787879 0 0.0 1e-06 
0.888888888889 -0.787878787879 0 0.0 1e-06 
0.944444444444 -0.787878787879 0 0.0 1e-06 
1.0 -0.787878787879 0 0.0 1e-06 
0.5 -0.747474747475 0 0.0 1e-06 
0.555555555556 -0.747474747475 0 0.0 1e-06 
0.611111111111 -0.747474747475 0 0.0 1e-06 
0.666666666667 -0.747474747475 0 0.0 1e-06 
0.722222222222 -0.747474747475 0 0.0 1e-06 
0.777777777778 -0.747474747475 0 0.0 1e-06 
0.833333333333 -0.747474747475 0 0.0 1e-06 
0.888888888889 -0.747474747475 0 0.0 1e-06 
0.944444444444 -0.747474747475 0 0.0 1e-06 
1.0 -0.747474747475 0 0.0 1e-06 
0.5 -0.707070707071 0 0.0 1e-06 
0.555555555556 -0.707070707071 0 0.0 1e-06 
0.611111111111 -0.707070707071 0 0.0 1e-06 
0.666666666667 -0.707070707071 0 0.0 1e-06 
0.722222222222 -0.707070707071 0 0.0 1e-06 
0.777777777778 -0.707070707071 0 0.0 1e-06 
0.833333333333 -0.707070707071 0 0.0 1e-06 
0.888888888889 -0.707070707071 0 0.0 1e-06 
0.944444444444 -0.707070707071 0 0.0 1e-06 
1.0 -0.707070707071 0 0.0 1e-06 
0.5 -0.666666666667 0 0.0 1e-06 
0.555555555556 -0.666666666667 0 0.0 1e-06 
0.611111111111 -0.666666666667 0 0.0 1e-06 
0.666666666667 -0.666666666667 0 0.0 1e-06 
0.722222222222 -0.666666666667 0 0.0 1e-06 
0.777777777778 -0.666666666667 0 0.0 1e-06 
0.833333333333 -0.666666666667 0 0.0 1e-06 
0.888888888889 -0.666666666667 0 0.0 1e-06 
0.944444444444 -0.666666666667 0 0.0 1e-06 
1.0 -0.666666666667 0 0.0 1e-06 
0.5 -0.626262626263 0 0.0 1e-06 
0.555555555556 -0.626262626263 0 0.0 1e-06 
0.611111111111 -0.626262626263 0 0.0 1e-06 
0.666666666667 -0.626262626263 0 0.0 1e-06 
0.722222222222 -0.626262626263 0 0.0 1e-06 
0.777777777778 -0.626262626263 0 0.0 1e-06 
0.833333333333 -0.626262626263 0 0.0 1e-06 
0.888888888889 -0.626262626263 0 0.0 1e-06 
0.944444444444 -0.626262626263 0 0.0 1e-06 
1.0 -0.626262626263 0 0.0 1e-06 
0.5 -0.585858585859 0 0.0 1e-06 
0.555555555556 -0.585858585859 0 0.0 1e-06 
0.611111111111 -0.585858585859 0 0.0 1e-06 
0.666666666667 -0.585858585859 0 0.0 1e-06 
0.722222222222 -0.585858585859 0 0.0 1e-06 
0.777777777778 -0.585858585859 0 0.0 1e-06 
0.833333333333 -0.585858585859 0 0.0 1e-06 
0.888888888889 -0.585858585859 0 0.0 1e-06 
0.944444444444 -0.585858585859 0 0.0 1e-06 
1.0 -0.585858585859 0 0.0 1e-06 
0.5 -0.545454545455 0 0.0 1e-06 
0.555555555556 -0.545454545455 0 0.0 1e-06 
0.611111111111 -0.545454545455 0 0.0 1e-06 
0.666666666667 -0.545454545455 0 0.0 1e-06 
0.722222222222 -0.545454545455 0 0.0 1e-06 
0.777777777778 -0.545454545455 0 0.0 1e-06 
0.833333333333 -0.545454545455 0 0.0 1e-06 
0.888888888889 -0.545454545455 0 0.0 1e-06 
0.944444444444 -0.545454545455 0 0.0 1e-06 
1.0 -0.545454545455 0 0.0 1e-06 
0.5 -0.505050505051 0 0.0 1e-06 
0.555555555556 -0.505050505051 0 0.0 1e-06 
0.611111111111 -0.505050505051 0 0.0 1e-06 
0.666666666667 -0.505050505051 0 0.0 1e-06 
0.722222222222 -0.505050505051 0 0.0 1e-06 
0.777777777778 -0.505050505051 0 0.0 1e-06 
0.833333333333 -0.505050505051 0 0.0 1e-06 
0.888888888889 -0.505050505051 0 0.0 1e-06 
0.944444444444 -0.505050505051 0 0.0 1e-06 
1.0 -0.505050505051 0 0.0 1e-06 
0.5 -0.464646464646 0 0.0 1e-06 
0.555555555556 -0.464646464646 0 0.0 1e-06 
0.611111111111 -0.464646464646 0 0.0 1e-06 
0.666666666667 -0.464646464646 0 0.0 1e-06 
0.722222222222 -0.464646464646 0 0.0 1e-06 
0.777777777778 -0.464646464646 0 0.0 1e-06 
0.833333333333 -0.464646464646 0 0.0 1e-06 
0.888888888889 -0.464646464646 0 0.0 1e-06 
0.944444444444 -0.464646464646 0 0.0 1e-06 
1.0 -0.464646464646 0 0.0 1e-06 
0.5 -0.424242424242 0 0.0 1e-06 
0.555555555556 -0.424242424242 0 0.0 1e-06 
0.611111111111 -0.424242424242 0 0.0 1e-06 
0.666666666667 -0.424242424242 0 0.0 1e-06 
0.722222222222 -0.424242424242 0 0.0 1e-06 
0.777777777778 -0.424242424242 0 0.0 1e-06 
0.833333333333 -0.424242424242 0 0.0 1e-06 
0.888888888889 -0.424242424242 0 0.0 1e-06 
0.944444444444 -0.424242424242 0 0.0 1e-06 
1.0 -0.424242424242 0 0.0 1e-06 
0.5 -0.383838383838 0 0.0 1e-06 
0.555555555556 -0.383838383838 0 0.0 1e-06 
0.611111111111 -0.383838383838 0 0.0 1e-06 
0.666666666667 -0.383838383838 0 0.0 1e-06 
0.722222222222 -0.383838383838 0 0.0 1e-06 
0.777777777778 -0.383838383838 0 0.0 1e-06 
0.833333333333 -0.383838383838 0 0.0 1e-06 
0.888888888889 -0.383838383838 0 0.0 1e-06 
0.944444444444 -0.383838383838 0 0.0 1e-06 
1.0 -0.383838383838 0 0.0 1e-06 
0.5 -0.343434343434 0 0.0 1e-06 
0.555555555556 -0.343434343434 0 0.0 1e-06 
0.611111111111 -0.343434343434 0 0.0 1e-06 
0.666666666667 -0.343434343434 0 0.0 1e-06 
0.722222222222 -0.343434343434 0 0.0 1e-06 
0.777777777778 -0.343434343434 0 0.0 1e-06 
0.833333333333 -0.343434343434 0 0.0 1e-06 
0.888888888889 -0.343434343434 0 0.0 1e-06 
0.944444444444 -0.343434343434 0 0.0 1e-06 
1.0 -0.343434343434 0 0.0 1e-06 
0.5 -0.30303030303 0 0.0 1e-06 
0.555555555556 -0.30303030303 0 0.0 1e-06 
0.611111111111 -0.30303030303 0 0.0 1e-06 
0.666666666667 -0.30303030303 0 0.0 1e-06 
0.722222222222 -0.30303030303 0 0.0 1e-06 
0.777777777778 -0.30303030303 0 0.0 1e-06 
0.833333333333 -0.30303030303 0 0.0 1e-06 
0.888888888889 -0.30303030303 0 0.0 1e-06 
0.944444444444 -0.30303030303 0 0.0 1e-06 
1.0 -0.30303030303 0 0.0 1e-06 
0.5 -0.262626262626 0 0.0 1e-06 
0.555555555556 -0.262626262626 0 0.0 1e-06 
0.611111111111 -0.262626262626 0 0.0 1e-06 
0.666666666667 -0.262626262626 0 0.0 1e-06 
0.722222222222 -0.262626262626 0 0.0 1e-06 
0.777777777778 -0.262626262626 0 0.0 1e-06 
0.833333333333 -0.262626262626 0 0.0 1e-06 
0.888888888889 -0.262626262626 0 0.0 1e-06 
0.944444444444 -0.262626262626 0 0.0 1e-06 
1.0 -0.262626262626 0 0.0 1e-06 
0.5 -0.222222222222 0 0.0 1e-06 
0.555555555556 -0.222222222222 0 0.0 1e-06 
0.611111111111 -0.222222222222 0 0.0 1e-06 
0.666666666667 -0.222222222222 0 0.0 1e-06 
0.722222222222 -0.222222222222 0 0.0 1e-06 
0.777777777778 -0.222222222222 0 0.0 1e-06 
0.833333333333 -0.222222222222 0 0.0 1e-06 
0.888888888889 -0.222222222222 0 0.0 1e-06 
0.944444444444 -0.222222222222 0 0.0 1e-06 
1.0 -0.222222222222 0 0.0 1e-06 
0.5 -0.181818181818 0 0.0 1e-06 
0.555555555556 -0.181818181818 0 0.0 1e-06 
0.611111111111 -0.181818181818 0 0.0 1e-06 
0.666666666667 -0.181818181818 0 0.0 1e-06 
0.722222222222 -0.181818181818 0 0.0 1e-06 
0.777777777778 -0.181818181818 0 0.0 1e-06 
0.833333333333 -0.181818181818 0 0.0 1e-06 
0.888888888889 -0.181818181818 0 0.0 1e-06 
0.944444444444 -0.181818181818 0 0.0 1e-06 
1.0 -0.181818181818 0 0.0 1e-06 
0.5 -0.141414141414 0 0.0 1e-06 
0.555555555556 -0.141414141414 0 0.0 1e-06 
0.611111111111 -0.141414141414 0 0.0 1e-06 
0.666666666667 -0.141414141414 0 0.0 1e-06 
0.722222222222 -0.141414141414 0 0.0 1e-06 
0.777777777778 -0.141414141414 0 0.0 1e-06 
0.833333333333 -0.141414141414 0 0.0 1e-06 
0.888888888889 -0.141414141414 0 0.0 1e-06 
0.944444444444 -0.141414141414 0 0.0 1e-06 
1.0 -0.141414141414 0 0.0 1e-06 
0.5 -0.10101010101 0 0.0 1e-06 
0.555555555556 -0.10101010101 0 0.0 1e-06 
0.611111111111 -0.10101010101 0 0.0 1e-06 
0.666666666667 -0.10101010101 0 0.0 1e-06 
0.722222222222 -0.10101010101 0 0.0 1e-06 
0.777777777778 -0.10101010101 0 0.0 1e-06 
0.833333333333 -0.10101010101 0 0.0 1e-06 
0.888888888889 -0.10101010101 0 0.0 1e-06 
0.944444444444 -0.10101010101 0 0.0 1e-06 
1.0 -0.10101010101 0 0.0 1e-06 
0.5 -0.0606060606061 0 0.0 1e-06 
0.555555555556 -0.0606060606061 0 0.0 1e-06 
0.611111111111 -0.0606060606061 0 0.0 1e-06 
0.666666666667 -0.0606060606061 0 0.0 1e-06 
0.722222222222 -0.0606060606061 0 0.0 1e-06 
0.777777777778 -0.0606060606061 0 0.0 1e-06 
0.833333333333 -0.0606060606061 0 0.0 1e-06 
0.888888888889 -0.0606060606061 0 0.0 1e-06 
0.944444444444 -0.0606060606061 0 0.0 1e-06 
1.0 -0.0606060606061 0 0.0 1e-06 
0.5 -0.020202020202 0 0.0 1e-06 
0.555555555556 -0.020202020202 0 0.0 1e-06 
0.611111111111 -0.020202020202 0 0.0 1e-06 
0.666666666667 -0.020202020202 0 0.0 1e-06 
0.722222222222 -0.020202020202 0 0.0 1e-06 
0.777777777778 -0.020202020202 0 0.0 1e-06 
0.833333333333 -0.020202020202 0 0.0 1e-06 
0.888888888889 -0.020202020202 0 0.0 1e-06 
0.944444444444 -0.020202020202 0 0.0 1e-06 
1.0 -0.020202020202 0 0.0 1e-06 
0.5 0.020202020202 0 0.0 1e-06 
0.555555555556 0.020202020202 0 0.0 1e-06 
0.611111111111 0.020202020202 0 0.0 1e-06 
0.666666666667 0.020202020202 0 0.0 1e-06 
0.722222222222 0.020202020202 0 0.0 1e-06 
0.777777777778 0.020202020202 0 0.0 1e-06 
0.833333333333 0.020202020202 0 0.0 1e-06 
0.888888888889 0.020202020202 0 0.0 1e-06 
0.944444444444 0.020202020202 0 0.0 1e-06 
1.0 0.020202020202 0 0.0 1e-06 
0.5 0.0606060606061 0 0.0 1e-06 
0.555555555556 0.0606060606061 0 0.0 1e-06 
0.611111111111 0.0606060606061 0 0.0 1e-06 
0.666666666667 0.0606060606061 0 0.0 1e-06 
0.722222222222 0.0606060606061 0 0.0 1e-06 
0.777777777778 0.0606060606061 0 0.0 1e-06 
0.833333333333 0.0606060606061 0 0.0 1e-06 
0.888888888889 0.0606060606061 0 0.0 1e-06 
0.944444444444 0.0606060606061 0 0.0 1e-06 
1.0 0.0606060606061 0 0.0 1e-06 
0.5 0.10101010101 0 0.0 1e-06 
0.555555555556 0.10101010101 0 0.0 1e-06 
0.611111111111 0.10101010101 0 0.0 1e-06 
0.666666666667 0.10101010101 0 0.0 1e-06 
0.722222222222 0.10101010101 0 0.0 1e-06 
0.777777777778 0.10101010101 0 0.0 1e-06 
0.833333333333 0.10101010101 0 0.0 1e-06 
0.888888888889 0.10101010101 0 0.0 1e-06 
0.944444444444 0.10101010101 0 0.0 1e-06 
1.0 0.10101010101 0 0.0 1e-06 
0.5 0.141414141414 0 0.0 1e-06 
0.555555555556 0.141414141414 0 0.0 1e-06 
0.611111111111 0.141414141414 0 0.0 1e-06 
0.666666666667 0.141414141414 0 0.0 1e-06 
0.722222222222 0.141414141414 0 0.0 1e-06 
0.777777777778 0.141414141414 0 0.0 1e-06 
0.833333333333 0.141414141414 0 0.0 1e-06 
0.888888888889 0.141414141414 0 0.0 1e-06 
0.944444444444 0.141414141414 0 0.0 1e-06 
1.0 0.141414141414 0 0.0 1e-06 
0.5 0.181818181818 0 0.0 1e-06 
0.555555555556 0.181818181818 0 0.0 1e-06 
0.611111111111 0.181818181818 0 0.0 1e-06 
0.666666666667 0.181818181818 0 0.0 1e-06 
0.722222222222 0.181818181818 0 0.0 1e-06 
0.777777777778 0.181818181818 0 0.0 1e-06 
0.833333333333 0.181818181818 0 0.0 1e-06 
0.888888888889 0.181818181818 0 0.0 1e-06 
0.944444444444 0.181818181818 0 0.0 1e-06 
1.0 0.181818181818 0 0.0 1e-06 
0.5 0.222222222222 0 0.0 1e-06 
0.555555555556 0.222222222222 0 0.0 1e-06 
0.611111111111 0.222222222222 0 0.0 1e-06 
0.666666666667 0.222222222222 0 0.0 1e-06 
0.722222222222 0.222222222222 0 0.0 1e-06 
0.777777777778 0.222222222222 0 0.0 1e-06 
0.833333333333 0.222222222222 0 0.0 1e-06 
0.888888888889 0.222222222222 0 0.0 1e-06 
0.944444444444 0.222222222222 0 0.0 1e-06 
1.0 0.222222222222 0 0.0 1e-06 
0.5 0.262626262626 0 0.0 1e-06 
0.555555555556 0.262626262626 0 0.0 1e-06 
0.611111111111 0.262626262626 0 0.0 1e-06 
0.666666666667 0.262626262626 0 0.0 1e-06 
0.722222222222 0.262626262626 0 0.0 1e-06 
0.777777777778 0.262626262626 0 0.0 1e-06 
0.833333333333 0.262626262626 0 0.0 1e-06 
0.888888888889 0.262626262626 0 0.0 1e-06 
0.944444444444 0.262626262626 0 0.0 1e-06 
1.0 0.262626262626 0 0.0 1e-06 
0.5 0.30303030303 0 0.0 1e-06 
0.555555555556 0.30303030303 0 0.0 1e-06 
0.611111111111 0.30303030303 0 0.0 1e-06 
0.666666666667 0.30303030303 0 0.0 1e-06 
0.722222222222 0.30303030303 0 0.0 1e-06 
0.777777777778 0.30303030303 0 0.0 1e-06 
0.833333333333 0.30303030303 0 0.0 1e-06 
0.888888888889 0.30303030303 0 0.0 1e-06 
0.944444444444 0.30303030303 0 0.0 1e-06 
1.0 0.30303030303 0 0.0 1e-06 
0.5 0.343434343434 0 0.0 1e-06 
0.555555555556 0.343434343434 0 0.0 1e-06 
0.611111111111 0.343434343434 0 0.0 1e-06 
0.666666666667 0.343434343434 0 0.0 1e-06 
0.722222222222 0.343434343434 0 0.0 1e-06 
0.777777777778 0.343434343434 0 0.0 1e-06 
0.833333333333 0.343434343434 0 0.0 1e-06 
0.888888888889 0.343434343434 0 0.0 1e-06 
0.944444444444 0.343434343434 0 0.0 1e-06 
1.0 0.343434343434 0 0.0 1e-06 
0.5 0.383838383838 0 0.0 1e-06 
0.555555555556 0.383838383838 0 0.0 1e-06 
0.611111111111 0.383838383838 0 0.0 1e-06 
0.666666666667 0.383838383838 0 0.0 1e-06 
0.722222222222 0.383838383838 0 0.0 1e-06 
0.777777777778 0.383838383838 0 0.0 1e-06 
0.833333333333 0.383838383838 0 0.0 1e-06 
0.888888888889 0.383838383838 0 0.0 1e-06 
0.944444444444 0.383838383838 0 0.0 1e-06 
1.0 0.383838383838 0 0.0 1e-06 
0.5 0.424242424242 0 0.0 1e-06 
0.555555555556 0.424242424242 0 0.0 1e-06 
0.611111111111 0.424242424242 0 0.0 1e-06 
0.666666666667 0.424242424242 0 0.0 1e-06 
0.722222222222 0.424242424242 0 0.0 1e-06 
0.777777777778 0.424242424242 0 0.0 1e-06 
0.833333333333 0.424242424242 0 0.0 1e-06 
0.888888888889 0.424242424242 0 0.0 1e-06 
0.944444444444 0.424242424242 0 0.0 1e-06 
1.0 0.424242424242 0 0.0 1e-06 
0.5 0.464646464646 0 0.0 1e-06 
0.555555555556 0.464646464646 0 0.0 1e-06 
0.611111111111 0.464646464646 0 0.0 1e-06 
0.666666666667 0.464646464646 0 0.0 1e-06 
0.722222222222 0.464646464646 0 0.0 1e-06 
0.777777777778 0.464646464646 0 0.0 1e-06 
0.833333333333 0.464646464646 0 0.0 1e-06 
0.888888888889 0.464646464646 0 0.0 1e-06 
0.944444444444 0.464646464646 0 0.0 1e-06 
1.0 0.464646464646 0 0.0 1e-06 
0.5 0.505050505051 0 0.0 1e-06 
0.555555555556 0.505050505051 0 0.0 1e-06 
0.611111111111 0.505050505051 0 0.0 1e-06 
0.666666666667 0.505050505051 0 0.0 1e-06 
0.722222222222 0.505050505051 0 0.0 1e-06 
0.777777777778 0.505050505051 0 0.0 1e-06 
0.833333333333 0.505050505051 0 0.0 1e-06 
0.888888888889 0.505050505051 0 0.0 1e-06 
0.944444444444 0.505050505051 0 0.0 1e-06 
1.0 0.505050505051 0 0.0 1e-06 
0.5 0.545454545455 0 0.0 1e-06 
0.555555555556 0.545454545455 0 0.0 1e-06 
0.611111111111 0.545454545455 0 0.0 1e-06 
0.666666666667 0.545454545455 0 0.0 1e-06 
0.722222222222 0.545454545455 0 0.0 1e-06 
0.777777777778 0.545454545455 0 0.0 1e-06 
0.833333333333 0.545454545455 0 0.0 1e-06 
0.888888888889 0.545454545455 0 0.0 1e-06 
0.944444444444 0.545454545455 0 0.0 1e-06 
1.0 0.545454545455 0 0.0 1e-06 
0.5 0.585858585859 0 0.0 1e-06 
0.555555555556 0.585858585859 0 0.0 1e-06 
0.611111111111 0.585858585859 0 0.0 1e-06 
0.666666666667 0.585858585859 0 0.0 1e-06 
0.722222222222 0.585858585859 0 0.0 1e-06 
0.777777777778 0.585858585859 0 0.0 1e-06 
0.833333333333 0.585858585859 0 0.0 1e-06 
0.888888888889 0.585858585859 0 0.0 1e-06 
0.944444444444 0.585858585859 0 0.0 1e-06 
1.0 0.585858585859 0 0.0 1e-06 
0.5 0.626262626263 0 0.0 1e-06 
0.555555555556 0.626262626263 0 0.0 1e-06 
0.611111111111 0.626262626263 0 0.0 1e-06 
0.666666666667 0.626262626263 0 0.0 1e-06 
0.722222222222 0.626262626263 0 0.0 1e-06 
0.777777777778 0.626262626263 0 0.0 1e-06 
0.833333333333 0.626262626263 0 0.0 1e-06 
0.888888888889 0.626262626263 0 0.0 1e-06 
0.944444444444 0.626262626263 0 0.0 1e-06 
1.0 0.626262626263 0 0.0 1e-06 
0.5 0.666666666667 0 0.0 1e-06 
0.555555555556 0.666666666667 0 0.0 1e-06 
0.611111111111 0.666666666667 0 0.0 1e-06 
0.666666666667 0.666666666667 0 0.0 1e-06 
0.722222222222 0.666666666667 0 0.0 1e-06 
0.777777777778 0.666666666667 0 0.0 1e-06 
0.833333333333 0.666666666667 0 0.0 1e-06 
0.888888888889 0.666666666667 0 0.0 1e-06 
0.944444444444 0.666666666667 0 0.0 1e-06 
1.0 0.666666666667 0 0.0 1e-06 
0.5 0.707070707071 0 0.0 1e-06 
0.555555555556 0.707070707071 0 0.0 1e-06 
0.611111111111 0.707070707071 0 0.0 1e-06 
0.666666666667 0.707070707071 0 0.0 1e-06 
0.722222222222 0.707070707071 0 0.0 1e-06 
0.777777777778 0.707070707071 0 0.0 1e-06 
0.833333333333 0.707070707071 0 0.0 1e-06 
0.888888888889 0.707070707071 0 0.0 1e-06 
0.944444444444 0.707070707071 0 0.0 1e-06 
1.0 0.707070707071 0 0.0 1e-06 
0.5 0.747474747475 0 0.0 1e-06 
0.555555555556 0.747474747475 0 0.0 1e-06 
0.611111111111 0.747474747475 0 0.0 1e-06 
0.666666666667 0.747474747475 0 0.0 1e-06 
0.722222222222 0.747474747475 0 0.0 1e-06 
0.777777777778 0.747474747475 0 0.0 1e-06 
0.833333333333 0.747474747475 0 0.0 1e-06 
0.888888888889 0.747474747475 0 0.0 1e-06 
0.944444444444 0.747474747475 0 0.0 1e-06 
1.0 0.747474747475 0 0.0 1e-06 
0.5 0.787878787879 0 0.0 1e-06 
0.555555555556 0.787878787879 0 0.0 1e-06 
0.611111111111 0.787878787879 0 0.0 1e-06 
0.666666666667 0.787878787879 0 0.0 1e-06 
0.722222222222 0.787878787879 0 0.0 1e-06 
0.777777777778 0.787878787879 0 0.0 1e-06 
0.833333333333 0.787878787879 0 0.0 1e-06 
0.888888888889 0.787878787879 0 0.0 1e-06 
0.944444444444 0.787878787879 0 0.0 1e-06 
1.0 0.787878787879 0 0.0 1e-06 
0.5 0.828282828283 0 0.0 1e-06 
0.555555555556 0.828282828283 0 0.0 1e-06 
0.611111111111 0.828282828283 0 0.0 1e-06 
0.666666666667 0.828282828283 0 0.0 1e-06 
0.722222222222 0.828282828283 0 0.0 1e-06 
0.777777777778 0.828282828283 0 0.0 1e-06 
0.833333333333 0.828282828283 0 0.0 1e-06 
0.888888888889 0.828282828283 0 0.0 1e-06 
0.944444444444 0.828282828283 0 0.0 1e-06 
1.0 0.828282828283 0 0.0 1e-06 
0.5 0.868686868687 0 0.0 1e-06 
0.555555555556 0.868686868687 0 0.0 1e-06 
0.611111111111 0.868686868687 0 0.0 1e-06 
0.666666666667 0.868686868687 0 0.0 1e-06 
0.722222222222 0.868686868687 0 0.0 1e-06 
0.777777777778 0.868686868687 0 0.0 1e-06 
0.833333333333 0.868686868687 0 0.0 1e-06 
0.888888888889 0.868686868687 0 0.0 1e-06 
0.944444444444 0.868686868687 0 0.0 1e-06 
1.0 0.868686868687 0 0.0 1e-06 
0.5 0.909090909091 0 0.0 1e-06 
0.555555555556 0.909090909091 0 0.0 1e-06 
0.611111111111 0.909090909091 0 0.0 1e-06 
0.666666666667 0.909090909091 0 0.0 1e-06 
0.722222222222 0.909090909091 0 0.0 1e-06 
0.777777777778 0.909090909091 0 0.0 1e-06 
0.833333333333 0.909090909091 0 0.0 1e-06 
0.888888888889 0.909090909091 0 0.0 1e-06 
0.944444444444 0.909090909091 0 0.0 1e-06 
1.0 0.909090909091 0 0.0 1e-06 
0.5 0.949494949495 0 0.0 1e-06 
0.555555555556 0.949494949495 0 0.0 1e-06 
0.611111111111 0.949494949495 0 0.0 1e-06 
0.666666666667 0.949494949495 0 0.0 1e-06 
0.722222222222 0.949494949495 0 0.0 1e-06 
0.777777777778 0.949494949495 0 0.0 1e-06 
0.833333333333 0.949494949495 0 0.0 1e-06 
0.888888888889 0.949494949495 0 0.0 1e-06 
0.944444444444 0.949494949495 0 0.0 1e-06 
1.0 0.949494949495 0 0.0 1e-06 
0.5 0.989898989899 0 0.0 1e-06 
0.555555555556 0.989898989899 0 0.0 1e-06 
0.611111111111 0.989898989899 0 0.0 1e-06 
0.666666666667 0.989898989899 0 0.0 1e-06 
0.722222222222 0.989898989899 0 0.0 1e-06 
0.777777777778 0.989898989899 0 0.0 1e-06 
0.833333333333 0.989898989899 0 0.0 1e-06 
0.888888888889 0.989898989899 0 0.0 1e-06 
0.944444444444 0.989898989899 0 0.0 1e-06 
1.0 0.989898989899 0 0.0 1e-06 
0.5 1.0303030303 0 0.0 1e-06 
0.555555555556 1.0303030303 0 0.0 1e-06 
0.611111111111 1.0303030303 0 0.0 1e-06 
0.666666666667 1.0303030303 0 0.0 1e-06 
0.722222222222 1.0303030303 0 0.0 1e-06 
0.777777777778 1.0303030303 0 0.0 1e-06 
0.833333333333 1.0303030303 0 0.0 1e-06 
0.888888888889 1.0303030303 0 0.0 1e-06 
0.944444444444 1.0303030303 0 0.0 1e-06 
1.0 1.0303030303 0 0.0 1e-06 
0.5 1.07070707071 0 0.0 1e-06 
0.555555555556 1.07070707071 0 0.0 1e-06 
0.611111111111 1.07070707071 0 0.0 1e-06 
0.666666666667 1.07070707071 0 0.0 1e-06 
0.722222222222 1.07070707071 0 0.0 1e-06 
0.777777777778 1.07070707071 0 0.0 1e-06 
0.833333333333 1.07070707071 0 0.0 1e-06 
0.888888888889 1.07070707071 0 0.0 1e-06 
0.944444444444 1.07070707071 0 0.0 1e-06 
1.0 1.07070707071 0 0.0 1e-06 
0.5 1.11111111111 0 0.0 1e-06 
0.555555555556 1.11111111111 0 0.0 1e-06 
0.611111111111 1.11111111111 0 0.0 1e-06 
0.666666666667 1.11111111111 0 0.0 1e-06 
0.722222222222 1.11111111111 0 0.0 1e-06 
0.777777777778 1.11111111111 0 0.0 1e-06 
0.833333333333 1.11111111111 0 0.0 1e-06 
0.888888888889 1.11111111111 0 0.0 1e-06 
0.944444444444 1.11111111111 0 0.0 1e-06 
1.0 1.11111111111 0 0.0 1e-06 
0.5 1.15151515152 0 0.0 1e-06 
0.555555555556 1.15151515152 0 0.0 1e-06 
0.611111111111 1.15151515152 0 0.0 1e-06 
0.666666666667 1.15151515152 0 0.0 1e-06 
0.722222222222 1.15151515152 0 0.0 1e-06 
0.777777777778 1.15151515152 0 0.0 1e-06 
0.833333333333 1.15151515152 0 0.0 1e-06 
0.888888888889 1.15151515152 0 0.0 1e-06 
0.944444444444 1.15151515152 0 0.0 1e-06 
1.0 1.15151515152 0 0.0 1e-06 
0.5 1.19191919192 0 0.0 1e-06 
0.555555555556 1.19191919192 0 0.0 1e-06 
0.611111111111 1.19191919192 0 0.0 1e-06 
0.666666666667 1.19191919192 0 0.0 1e-06 
0.722222222222 1.19191919192 0 0.0 1e-06 
0.777777777778 1.19191919192 0 0.0 1e-06 
0.833333333333 1.19191919192 0 0.0 1e-06 
0.888888888889 1.19191919192 0 0.0 1e-06 
0.944444444444 1.19191919192 0 0.0 1e-06 
1.0 1.19191919192 0 0.0 1e-06 
0.5 1.23232323232 0 0.0 1e-06 
0.555555555556 1.23232323232 0 0.0 1e-06 
0.611111111111 1.23232323232 0 0.0 1e-06 
0.666666666667 1.23232323232 0 0.0 1e-06 
0.722222222222 1.23232323232 0 0.0 1e-06 
0.777777777778 1.23232323232 0 0.0 1e-06 
0.833333333333 1.23232323232 0 0.0 1e-06 
0.888888888889 1.23232323232 0 0.0 1e-06 
0.944444444444 1.23232323232 0 0.0 1e-06 
1.0 1.23232323232 0 0.0 1e-06 
0.5 1.27272727273 0 0.0 1e-06 
0.555555555556 1.27272727273 0 0.0 1e-06 
0.611111111111 1.27272727273 0 0.0 1e-06 
0.666666666667 1.27272727273 0 0.0 1e-06 
0.722222222222 1.27272727273 0 0.0 1e-06 
0.777777777778 1.27272727273 0 0.0 1e-06 
0.833333333333 1.27272727273 0 0.0 1e-06 
0.888888888889 1.27272727273 0 0.0 1e-06 
0.944444444444 1.27272727273 0 0.0 1e-06 
1.0 1.27272727273 0 0.0 1e-06 
0.5 1.31313131313 0 0.0 1e-06 
0.555555555556 1.31313131313 0 0.0 1e-06 
0.611111111111 1.31313131313 0 0.0 1e-06 
0.666666666667 1.31313131313 0 0.0 1e-06 
0.722222222222 1.31313131313 0 0.0 1e-06 
0.777777777778 1.31313131313 0 0.0 1e-06 
0.833333333333 1.31313131313 0 0.0 1e-06 
0.888888888889 1.31313131313 0 0.0 1e-06 
0.944444444444 1.31313131313 0 0.0 1e-06 
1.0 1.31313131313 0 0.0 1e-06 
0.5 1.35353535354 0 0.0 1e-06 
0.555555555556 1.35353535354 0 0.0 1e-06 
0.611111111111 1.35353535354 0 0.0 1e-06 
0.666666666667 1.35353535354 0 0.0 1e-06 
0.722222222222 1.35353535354 0 0.0 1e-06 
0.777777777778 1.35353535354 0 0.0 1e-06 
0.833333333333 1.35353535354 0 0.0 1e-06 
0.888888888889 1.35353535354 0 0.0 1e-06 
0.944444444444 1.35353535354 0 0.0 1e-06 
1.0 1.35353535354 0 0.0 1e-06 
0.5 1.39393939394 0 0.0 1e-06 
0.555555555556 1.39393939394 0 0.0 1e-06 
0.611111111111 1.39393939394 0 0.0 1e-06 
0.666666666667 1.39393939394 0 0.0 1e-06 
0.722222222222 1.39393939394 0 0.0 1e-06 
0.777777777778 1.39393939394 0 0.0 1e-06 
0.833333333333 1.39393939394 0 0.0 1e-06 
0.888888888889 1.39393939394 0 0.0 1e-06 
0.944444444444 1.39393939394 0 0.0 1e-06 
1.0 1.39393939394 0 0.0 1e-06 
0.5 1.43434343434 0 0.0 1e-06 
0.555555555556 1.43434343434 0 0.0 1e-06 
0.611111111111 1.43434343434 0 0.0 1e-06 
0.666666666667 1.43434343434 0 0.0 1e-06 
0.722222222222 1.43434343434 0 0.0 1e-06 
0.777777777778 1.43434343434 0 0.0 1e-06 
0.833333333333 1.43434343434 0 0.0 1e-06 
0.888888888889 1.43434343434 0 0.0 1e-06 
0.944444444444 1.43434343434 0 0.0 1e-06 
1.0 1.43434343434 0 0.0 1e-06 
0.5 1.47474747475 0 0.0 1e-06 
0.555555555556 1.47474747475 0 0.0 1e-06 
0.611111111111 1.47474747475 0 0.0 1e-06 
0.666666666667 1.47474747475 0 0.0 1e-06 
0.722222222222 1.47474747475 0 0.0 1e-06 
0.777777777778 1.47474747475 0 0.0 1e-06 
0.833333333333 1.47474747475 0 0.0 1e-06 
0.888888888889 1.47474747475 0 0.0 1e-06 
0.944444444444 1.47474747475 0 0.0 1e-06 
1.0 1.47474747475 0 0.0 1e-06 
0.5 1.51515151515 0 0.0 1e-06 
0.555555555556 1.51515151515 0 0.0 1e-06 
0.611111111111 1.51515151515 0 0.0 1e-06 
0.666666666667 1.51515151515 0 0.0 1e-06 
0.722222222222 1.51515151515 0 0.0 1e-06 
0.777777777778 1.51515151515 0 0.0 1e-06 
0.833333333333 1.51515151515 0 0.0 1e-06 
0.888888888889 1.51515151515 0 0.0 1e-06 
0.944444444444 1.51515151515 0 0.0 1e-06 
1.0 1.51515151515 0 0.0 1e-06 
0.5 1.55555555556 0 0.0 1e-06 
0.555555555556 1.55555555556 0 0.0 1e-06 
0.611111111111 1.55555555556 0 0.0 1e-06 
0.666666666667 1.55555555556 0 0.0 1e-06 
0.722222222222 1.55555555556 0 0.0 1e-06 
0.777777777778 1.55555555556 0 0.0 1e-06 
0.833333333333 1.55555555556 0 0.0 1e-06 
0.888888888889 1.55555555556 0 0.0 1e-06 
0.944444444444 1.55555555556 0 0.0 1e-06 
1.0 1.55555555556 0 0.0 1e-06 
0.5 1.59595959596 0 0.0 1e-06 
0.555555555556 1.59595959596 0 0.0 1e-06 
0.611111111111 1.59595959596 0 0.0 1e-06 
0.666666666667 1.59595959596 0 0.0 1e-06 
0.722222222222 1.59595959596 0 0.0 1e-06 
0.777777777778 1.59595959596 0 0.0 1e-06 
0.833333333333 1.59595959596 0 0.0 1e-06 
0.888888888889 1.59595959596 0 0.0 1e-06 
0.944444444444 1.59595959596 0 0.0 1e-06 
1.0 1.59595959596 0 0.0 1e-06 
0.5 1.63636363636 0 0.0 1e-06 
0.555555555556 1.63636363636 0 0.0 1e-06 
0.611111111111 1.63636363636 0 0.0 1e-06 
0.666666666667 1.63636363636 0 0.0 1e-06 
0.722222222222 1.63636363636 0 0.0 1e-06 
0.777777777778 1.63636363636 0 0.0 1e-06 
0.833333333333 1.63636363636 0 0.0 1e-06 
0.888888888889 1.63636363636 0 0.0 1e-06 
0.944444444444 1.63636363636 0 0.0 1e-06 
1.0 1.63636363636 0 0.0 1e-06 
0.5 1.67676767677 0 0.0 1e-06 
0.555555555556 1.67676767677 0 0.0 1e-06 
0.611111111111 1.67676767677 0 0.0 1e-06 
0.666666666667 1.67676767677 0 0.0 1e-06 
0.722222222222 1.67676767677 0 0.0 1e-06 
0.777777777778 1.67676767677 0 0.0 1e-06 
0.833333333333 1.67676767677 0 0.0 1e-06 
0.888888888889 1.67676767677 0 0.0 1e-06 
0.944444444444 1.67676767677 0 0.0 1e-06 
1.0 1.67676767677 0 0.0 1e-06 
0.5 1.71717171717 0 0.0 1e-06 
0.555555555556 1.71717171717 0 0.0 1e-06 
0.611111111111 1.71717171717 0 0.0 1e-06 
0.666666666667 1.71717171717 0 0.0 1e-06 
0.722222222222 1.71717171717 0 0.0 1e-06 
0.777777777778 1.71717171717 0 0.0 1e-06 
0.833333333333 1.71717171717 0 0.0 1e-06 
0.888888888889 1.71717171717 0 0.0 1e-06 
0.944444444444 1.71717171717 0 0.0 1e-06 
1.0 1.71717171717 0 0.0 1e-06 
0.5 1.75757575758 0 0.0 1e-06 
0.555555555556 1.75757575758 0 0.0 1e-06 
0.611111111111 1.75757575758 0 0.0 1e-06 
0.666666666667 1.75757575758 0 0.0 1e-06 
0.722222222222 1.75757575758 0 0.0 1e-06 
0.777777777778 1.75757575758 0 0.0 1e-06 
0.833333333333 1.75757575758 0 0.0 1e-06 
0.888888888889 1.75757575758 0 0.0 1e-06 
0.944444444444 1.75757575758 0 0.0 1e-06 
1.0 1.75757575758 0 0.0 1e-06 
0.5 1.79797979798 0 0.0 1e-06 
0.555555555556 1.79797979798 0 0.0 1e-06 
0.611111111111 1.79797979798 0 0.0 1e-06 
0.666666666667 1.79797979798 0 0.0 1e-06 
0.722222222222 1.79797979798 0 0.0 1e-06 
0.777777777778 1.79797979798 0 0.0 1e-06 
0.833333333333 1.79797979798 0 0.0 1e-06 
0.888888888889 1.79797979798 0 0.0 1e-06 
0.944444444444 1.79797979798 0 0.0 1e-06 
1.0 1.79797979798 0 0.0 1e-06 
0.5 1.83838383838 0 0.0 1e-06 
0.555555555556 1.83838383838 0 0.0 1e-06 
0.611111111111 1.83838383838 0 0.0 1e-06 
0.666666666667 1.83838383838 0 0.0 1e-06 
0.722222222222 1.83838383838 0 0.0 1e-06 
0.777777777778 1.83838383838 0 0.0 1e-06 
0.833333333333 1.83838383838 0 0.0 1e-06 
0.888888888889 1.83838383838 0 0.0 1e-06 
0.944444444444 1.83838383838 0 0.0 1e-06 
1.0 1.83838383838 0 0.0 1e-06 
0.5 1.87878787879 0 0.0 1e-06 
0.555555555556 1.87878787879 0 0.0 1e-06 
0.611111111111 1.87878787879 0 0.0 1e-06 
0.666666666667 1.87878787879 0 0.0 1e-06 
0.722222222222 1.87878787879 0 0.0 1e-06 
0.777777777778 1.87878787879 0 0.0 1e-06 
0.833333333333 1.87878787879 0 0.0 1e-06 
0.888888888889 1.87878787879 0 0.0 1e-06 
0.944444444444 1.87878787879 0 0.0 1e-06 
1.0 1.87878787879 0 0.0 1e-06 
0.5 1.91919191919 0 0.0 1e-06 
0.555555555556 1.91919191919 0 0.0 1e-06 
0.611111111111 1.91919191919 0 0.0 1e-06 
0.666666666667 1.91919191919 0 0.0 1e-06 
0.722222222222 1.91919191919 0 0.0 1e-06 
0.777777777778 1.91919191919 0 0.0 1e-06 
0.833333333333 1.91919191919 0 0.0 1e-06 
0.888888888889 1.91919191919 0 0.0 1e-06 
0.944444444444 1.91919191919 0 0.0 1e-06 
1.0 1.91919191919 0 0.0 1e-06 
0.5 1.9595959596 0 0.0 1e-06 
0.555555555556 1.9595959596 0 0.0 1e-06 
0.611111111111 1.9595959596 0 0.0 1e-06 
0.666666666667 1.9595959596 0 0.0 1e-06 
0.722222222222 1.9595959596 0 0.0 1e-06 
0.777777777778 1.9595959596 0 0.0 1e-06 
0.833333333333 1.9595959596 0 0.0 1e-06 
0.888888888889 1.9595959596 0 0.0 1e-06 
0.944444444444 1.9595959596 0 0.0 1e-06 
1.0 1.9595959596 0 0.0 1e-06 
0.5 2.0 0 0.0 1e-06 
0.555555555556 2.0 0 0.0 1e-06 
0.611111111111 2.0 0 0.0 1e-06 
0.666666666667 2.0 0 0.0 1e-06 
0.722222222222 2.0 0 0.0 1e-06 
0.777777777778 2.0 0 0.0 1e-06 
0.833333333333 2.0 0 0.0 1e-06 
0.888888888889 2.0 0 0.0 1e-06 
0.944444444444 2.0 0 0.0 1e-06 
1.0 2.0 0 0.0 1e-06 
0.5 -2.0 0 0.4 1e-06 
0.555555555556 -2.0 0 0.4 1e-06 
0.611111111111 -2.0 0 0.4 1e-06 
0.666666666667 -2.0 0 0.4 1e-06 
0.722222222222 -2.0 0 0.4 1e-06 
0.777777777778 -2.0 0 0.4 1e-06 
0.833333333333 -2.0 0 0.4 1e-06 
0.888888888889 -2.0 0 0.4 1e-06 
0.944444444444 -2.0 0 0.4 1e-06 
1.0 -2.0 0 0.4 1e-06 
0.5 -1.9595959596 0 0.4 1e-06 
0.555555555556 -1.9595959596 0 0.4 1e-06 
0.611111111111 -1.9595959596 0 0.4 1e-06 
0.666666666667 -1.9595959596 0 0.4 1e-06 
0.722222222222 -1.9595959596 0 0.4 1e-06 
0.777777777778 -1.9595959596 0 0.4 1e-06 
0.833333333333 -1.9595959596 0 0.4 1e-06 
0.888888888889 -1.9595959596 0 0.4 1e-06 
0.944444444444 -1.9595959596 0 0.4 1e-06 
1.0 -1.9595959596 0 0.4 1e-06 
0.5 -1.91919191919 0 0.4 1e-06 
0.555555555556 -1.91919191919 0 0.4 1e-06 
0.611111111111 -1.91919191919 0 0.4 1e-06 
0.666666666667 -1.91919191919 0 0.4 1e-06 
0.722222222222 -1.91919191919 0 0.4 1e-06 
0.777777777778 -1.91919191919 0 0.4 1e-06 
0.833333333333 -1.91919191919 0 0.4 1e-06 
0.888888888889 -1.91919191919 0 0.4 1e-06 
0.944444444444 -1.91919191919 0 0.4 1e-06 
1.0 -1.91919191919 0 0.4 1e-06 
0.5 -1.87878787879 0 0.4 1e-06 
0.555555555556 -1.87878787879 0 0.4 1e-06 
0.611111111111 -1.87878787879 0 0.4 1e-06 
0.666666666667 -1.87878787879 0 0.4 1e-06 
0.722222222222 -1.87878787879 0 0.4 1e-06 
0.777777777778 -1.87878787879 0 0.4 1e-06 
0.833333333333 -1.87878787879 0 0.4 1e-06 
0.888888888889 -1.87878787879 0 0.4 1e-06 
0.944444444444 -1.87878787879 0 0.4 1e-06 
1.0 -1.87878787879 0 0.4 1e-06 
0.5 -1.83838383838 0 0.4 1e-06 
0.555555555556 -1.83838383838 0 0.4 1e-06 
0.611111111111 -1.83838383838 0 0.4 1e-06 
0.666666666667 -1.83838383838 0 0.4 1e-06 
0.722222222222 -1.83838383838 0 0.4 1e-06 
0.777777777778 -1.83838383838 0 0.4 1e-06 
0.833333333333 -1.83838383838 0 0.4 1e-06 
0.888888888889 -1.83838383838 0 0.4 1e-06 
0.944444444444 -1.83838383838 0 0.4 1e-06 
1.0 -1.83838383838 0 0.4 1e-06 
0.5 -1.79797979798 0 0.4 1e-06 
0.555555555556 -1.79797979798 0 0.4 1e-06 
0.611111111111 -1.79797979798 0 0.4 1e-06 
0.666666666667 -1.79797979798 0 0.4 1e-06 
0.722222222222 -1.79797979798 0 0.4 1e-06 
0.777777777778 -1.79797979798 0 0.4 1e-06 
0.833333333333 -1.79797979798 0 0.4 1e-06 
0.888888888889 -1.79797979798 0 0.4 1e-06 
0.944444444444 -1.79797979798 0 0.4 1e-06 
1.0 -1.79797979798 0 0.4 1e-06 
0.5 -1.75757575758 0 0.4 1e-06 
0.555555555556 -1.75757575758 0 0.4 1e-06 
0.611111111111 -1.75757575758 0 0.4 1e-06 
0.666666666667 -1.75757575758 0 0.4 1e-06 
0.722222222222 -1.75757575758 0 0.4 1e-06 
0.777777777778 -1.75757575758 0 0.4 1e-06 
0.833333333333 -1.75757575758 0 0.4 1e-06 
0.888888888889 -1.75757575758 0 0.4 1e-06 
0.944444444444 -1.75757575758 0 0.4 1e-06 
1.0 -1.75757575758 0 0.4 1e-06 
0.5 -1.71717171717 0 0.4 1e-06 
0.555555555556 -1.71717171717 0 0.4 1e-06 
0.611111111111 -1.71717171717 0 0.4 1e-06 
0.666666666667 -1.71717171717 0 0.4 1e-06 
0.722222222222 -1.71717171717 0 0.4 1e-06 
0.777777777778 -1.71717171717 0 0.4 1e-06 
0.833333333333 -1.71717171717 0 0.4 1e-06 
0.888888888889 -1.71717171717 0 0.4 1e-06 
0.944444444444 -1.71717171717 0 0.4 1e-06 
1.0 -1.71717171717 0 0.4 1e-06 
0.5 -1.67676767677 0 0.4 1e-06 
0.555555555556 -1.67676767677 0 0.4 1e-06 
0.611111111111 -1.67676767677 0 0.4 1e-06 
0.666666666667 -1.67676767677 0 0.4 1e-06 
0.722222222222 -1.67676767677 0 0.4 1e-06 
0.777777777778 -1.67676767677 0 0.4 1e-06 
0.833333333333 -1.67676767677 0 0.4 1e-06 
0.888888888889 -1.67676767677 0 0.4 1e-06 
0.944444444444 -1.67676767677 0 0.4 1e-06 
1.0 -1.67676767677 0 0.4 1e-06 
0.5 -1.63636363636 0 0.4 1e-06 
0.555555555556 -1.63636363636 0 0.4 1e-06 
0.611111111111 -1.63636363636 0 0.4 1e-06 
0.666666666667 -1.63636363636 0 0.4 1e-06 
0.722222222222 -1.63636363636 0 0.4 1e-06 
0.777777777778 -1.63636363636 0 0.4 1e-06 
0.833333333333 -1.63636363636 0 0.4 1e-06 
0.888888888889 -1.63636363636 0 0.4 1e-06 
0.944444444444 -1.63636363636 0 0.4 1e-06 
1.0 -1.63636363636 0 0.4 1e-06 
0.5 -1.59595959596 0 0.4 1e-06 
0.555555555556 -1.59595959596 0 0.4 1e-06 
0.611111111111 -1.59595959596 0 0.4 1e-06 
0.666666666667 -1.59595959596 0 0.4 1e-06 
0.722222222222 -1.59595959596 0 0.4 1e-06 
0.777777777778 -1.59595959596 0 0.4 1e-06 
0.833333333333 -1.59595959596 0 0.4 1e-06 
0.888888888889 -1.59595959596 0 0.4 1e-06 
0.944444444444 -1.59595959596 0 0.4 1e-06 
1.0 -1.59595959596 0 0.4 1e-06 
0.5 -1.55555555556 0 0.4 1e-06 
0.555555555556 -1.55555555556 0 0.4 1e-06 
0.611111111111 -1.55555555556 0 0.4 1e-06 
0.666666666667 -1.55555555556 0 0.4 1e-06 
0.722222222222 -1.55555555556 0 0.4 1e-06 
0.777777777778 -1.55555555556 0 0.4 1e-06 
0.833333333333 -1.55555555556 0 0.4 1e-06 
0.888888888889 -1.55555555556 0 0.4 1e-06 
0.944444444444 -1.55555555556 0 0.4 1e-06 
1.0 -1.55555555556 0 0.4 1e-06 
0.5 -1.51515151515 0 0.4 1e-06 
0.555555555556 -1.51515151515 0 0.4 1e-06 
0.611111111111 -1.51515151515 0 0.4 1e-06 
0.666666666667 -1.51515151515 0 0.4 1e-06 
0.722222222222 -1.51515151515 0 0.4 1e-06 
0.777777777778 -1.51515151515 0 0.4 1e-06 
0.833333333333 -1.51515151515 0 0.4 1e-06 
0.888888888889 -1.51515151515 0 0.4 1e-06 
0.944444444444 -1.51515151515 0 0.4 1e-06 
1.0 -1.51515151515 0 0.4 1e-06 
0.5 -1.47474747475 0 0.4 1e-06 
0.555555555556 -1.47474747475 0 0.4 1e-06 
0.611111111111 -1.47474747475 0 0.4 1e-06 
0.666666666667 -1.47474747475 0 0.4 1e-06 
0.722222222222 -1.47474747475 0 0.4 1e-06 
0.777777777778 -1.47474747475 0 0.4 1e-06 
0.833333333333 -1.47474747475 0 0.4 1e-06 
0.888888888889 -1.47474747475 0 0.4 1e-06 
0.944444444444 -1.47474747475 0 0.4 1e-06 
1.0 -1.47474747475 0 0.4 1e-06 
0.5 -1.43434343434 0 0.4 1e-06 
0.555555555556 -1.43434343434 0 0.4 1e-06 
0.611111111111 -1.43434343434 0 0.4 1e-06 
0.666666666667 -1.43434343434 0 0.4 1e-06 
0.722222222222 -1.43434343434 0 0.4 1e-06 
0.777777777778 -1.43434343434 0 0.4 1e-06 
0.833333333333 -1.43434343434 0 0.4 1e-06 
0.888888888889 -1.43434343434 0 0.4 1e-06 
0.944444444444 -1.43434343434 0 0.4 1e-06 
1.0 -1.43434343434 0 0.4 1e-06 
0.5 -1.39393939394 0 0.4 1e-06 
0.555555555556 -1.39393939394 0 0.4 1e-06 
0.611111111111 -1.39393939394 0 0.4 1e-06 
0.666666666667 -1.39393939394 0 0.4 1e-06 
0.722222222222 -1.39393939394 0 0.4 1e-06 
0.777777777778 -1.39393939394 0 0.4 1e-06 
0.833333333333 -1.39393939394 0 0.4 1e-06 
0.888888888889 -1.39393939394 0 0.4 1e-06 
0.944444444444 -1.39393939394 0 0.4 1e-06 
1.0 -1.39393939394 0 0.4 1e-06 
0.5 -1.35353535354 0 0.4 1e-06 
0.555555555556 -1.35353535354 0 0.4 1e-06 
0.611111111111 -1.35353535354 0 0.4 1e-06 
0.666666666667 -1.35353535354 0 0.4 1e-06 
0.722222222222 -1.35353535354 0 0.4 1e-06 
0.777777777778 -1.35353535354 0 0.4 1e-06 
0.833333333333 -1.35353535354 0 0.4 1e-06 
0.888888888889 -1.35353535354 0 0.4 1e-06 
0.944444444444 -1.35353535354 0 0.4 1e-06 
1.0 -1.35353535354 0 0.4 1e-06 
0.5 -1.31313131313 0 0.4 1e-06 
0.555555555556 -1.31313131313 0 0.4 1e-06 
0.611111111111 -1.31313131313 0 0.4 1e-06 
0.666666666667 -1.31313131313 0 0.4 1e-06 
0.722222222222 -1.31313131313 0 0.4 1e-06 
0.777777777778 -1.31313131313 0 0.4 1e-06 
0.833333333333 -1.31313131313 0 0.4 1e-06 
0.888888888889 -1.31313131313 0 0.4 1e-06 
0.944444444444 -1.31313131313 0 0.4 1e-06 
1.0 -1.31313131313 0 0.4 1e-06 
0.5 -1.27272727273 0 0.4 1e-06 
0.555555555556 -1.27272727273 0 0.4 1e-06 
0.611111111111 -1.27272727273 0 0.4 1e-06 
0.666666666667 -1.27272727273 0 0.4 1e-06 
0.722222222222 -1.27272727273 0 0.4 1e-06 
0.777777777778 -1.27272727273 0 0.4 1e-06 
0.833333333333 -1.27272727273 0 0.4 1e-06 
0.888888888889 -1.27272727273 0 0.4 1e-06 
0.944444444444 -1.27272727273 0 0.4 1e-06 
1.0 -1.27272727273 0 0.4 1e-06 
0.5 -1.23232323232 0 0.4 1e-06 
0.555555555556 -1.23232323232 0 0.4 1e-06 
0.611111111111 -1.23232323232 0 0.4 1e-06 
0.666666666667 -1.23232323232 0 0.4 1e-06 
0.722222222222 -1.23232323232 0 0.4 1e-06 
0.777777777778 -1.23232323232 0 0.4 1e-06 
0.833333333333 -1.23232323232 0 0.4 1e-06 
0.888888888889 -1.23232323232 0 0.4 1e-06 
0.944444444444 -1.23232323232 0 0.4 1e-06 
1.0 -1.23232323232 0 0.4 1e-06 
0.5 -1.19191919192 0 0.4 1e-06 
0.555555555556 -1.19191919192 0 0.4 1e-06 
0.611111111111 -1.19191919192 0 0.4 1e-06 
0.666666666667 -1.19191919192 0 0.4 1e-06 
0.722222222222 -1.19191919192 0 0.4 1e-06 
0.777777777778 -1.19191919192 0 0.4 1e-06 
0.833333333333 -1.19191919192 0 0.4 1e-06 
0.888888888889 -1.19191919192 0 0.4 1e-06 
0.944444444444 -1.19191919192 0 0.4 1e-06 
1.0 -1.19191919192 0 0.4 1e-06 
0.5 -1.15151515152 0 0.4 1e-06 
0.555555555556 -1.15151515152 0 0.4 1e-06 
0.611111111111 -1.15151515152 0 0.4 1e-06 
0.666666666667 -1.15151515152 0 0.4 1e-06 
0.722222222222 -1.15151515152 0 0.4 1e-06 
0.777777777778 -1.15151515152 0 0.4 1e-06 
0.833333333333 -1.15151515152 0 0.4 1e-06 
0.888888888889 -1.15151515152 0 0.4 1e-06 
0.944444444444 -1.15151515152 0 0.4 1e-06 
1.0 -1.15151515152 0 0.4 1e-06 
0.5 -1.11111111111 0 0.4 1e-06 
0.555555555556 -1.11111111111 0 0.4 1e-06 
0.611111111111 -1.11111111111 0 0.4 1e-06 
0.666666666667 -1.11111111111 0 0.4 1e-06 
0.722222222222 -1.11111111111 0 0.4 1e-06 
0.777777777778 -1.11111111111 0 0.4 1e-06 
0.833333333333 -1.11111111111 0 0.4 1e-06 
0.888888888889 -1.11111111111 0 0.4 1e-06 
0.944444444444 -1.11111111111 0 0.4 1e-06 
1.0 -1.11111111111 0 0.4 1e-06 
0.5 -1.07070707071 0 0.4 1e-06 
0.555555555556 -1.07070707071 0 0.4 1e-06 
0.611111111111 -1.07070707071 0 0.4 1e-06 
0.666666666667 -1.07070707071 0 0.4 1e-06 
0.722222222222 -1.07070707071 0 0.4 1e-06 
0.777777777778 -1.07070707071 0 0.4 1e-06 
0.833333333333 -1.07070707071 0 0.4 1e-06 
0.888888888889 -1.07070707071 0 0.4 1e-06 
0.944444444444 -1.07070707071 0 0.4 1e-06 
1.0 -1.07070707071 0 0.4 1e-06 
0.5 -1.0303030303 0 0.4 1e-06 
0.555555555556 -1.0303030303 0 0.4 1e-06 
0.611111111111 -1.0303030303 0 0.4 1e-06 
0.666666666667 -1.0303030303 0 0.4 1e-06 
0.722222222222 -1.0303030303 0 0.4 1e-06 
0.777777777778 -1.0303030303 0 0.4 1e-06 
0.833333333333 -1.0303030303 0 0.4 1e-06 
0.888888888889 -1.0303030303 0 0.4 1e-06 
0.944444444444 -1.0303030303 0 0.4 1e-06 
1.0 -1.0303030303 0 0.4 1e-06 
0.5 -0.989898989899 0 0.4 1e-06 
0.555555555556 -0.989898989899 0 0.4 1e-06 
0.611111111111 -0.989898989899 0 0.4 1e-06 
0.666666666667 -0.989898989899 0 0.4 1e-06 
0.722222222222 -0.989898989899 0 0.4 1e-06 
0.777777777778 -0.989898989899 0 0.4 1e-06 
0.833333333333 -0.989898989899 0 0.4 1e-06 
0.888888888889 -0.989898989899 0 0.4 1e-06 
0.944444444444 -0.989898989899 0 0.4 1e-06 
1.0 -0.989898989899 0 0.4 1e-06 
0.5 -0.949494949495 0 0.4 1e-06 
0.555555555556 -0.949494949495 0 0.4 1e-06 
0.611111111111 -0.949494949495 0 0.4 1e-06 
0.666666666667 -0.949494949495 0 0.4 1e-06 
0.722222222222 -0.949494949495 0 0.4 1e-06 
0.777777777778 -0.949494949495 0 0.4 1e-06 
0.833333333333 -0.949494949495 0 0.4 1e-06 
0.888888888889 -0.949494949495 0 0.4 1e-06 
0.944444444444 -0.949494949495 0 0.4 1e-06 
1.0 -0.949494949495 0 0.4 1e-06 
0.5 -0.909090909091 0 0.4 1e-06 
0.555555555556 -0.909090909091 0 0.4 1e-06 
0.611111111111 -0.909090909091 0 0.4 1e-06 
0.666666666667 -0.909090909091 0 0.4 1e-06 
0.722222222222 -0.909090909091 0 0.4 1e-06 
0.777777777778 -0.909090909091 0 0.4 1e-06 
0.833333333333 -0.909090909091 0 0.4 1e-06 
0.888888888889 -0.909090909091 0 0.4 1e-06 
0.944444444444 -0.909090909091 0 0.4 1e-06 
1.0 -0.909090909091 0 0.4 1e-06 
0.5 -0.868686868687 0 0.4 1e-06 
0.555555555556 -0.868686868687 0 0.4 1e-06 
0.611111111111 -0.868686868687 0 0.4 1e-06 
0.666666666667 -0.868686868687 0 0.4 1e-06 
0.722222222222 -0.868686868687 0 0.4 1e-06 
0.777777777778 -0.868686868687 0 0.4 1e-06 
0.833333333333 -0.868686868687 0 0.4 1e-06 
0.888888888889 -0.868686868687 0 0.4 1e-06 
0.944444444444 -0.868686868687 0 0.4 1e-06 
1.0 -0.868686868687 0 0.4 1e-06 
0.5 -0.828282828283 0 0.4 1e-06 
0.555555555556 -0.828282828283 0 0.4 1e-06 
0.611111111111 -0.828282828283 0 0.4 1e-06 
0.666666666667 -0.828282828283 0 0.4 1e-06 
0.722222222222 -0.828282828283 0 0.4 1e-06 
0.777777777778 -0.828282828283 0 0.4 1e-06 
0.833333333333 -0.828282828283 0 0.4 1e-06 
0.888888888889 -0.828282828283 0 0.4 1e-06 
0.944444444444 -0.828282828283 0 0.4 1e-06 
1.0 -0.828282828283 0 0.4 1e-06 
0.5 -0.787878787879 0 0.4 1e-06 
0.555555555556 -0.787878787879 0 0.4 1e-06 
0.611111111111 -0.787878787879 0 0.4 1e-06 
0.666666666667 -0.787878787879 0 0.4 1e-06 
0.722222222222 -0.787878787879 0 0.4 1e-06 
0.777777777778 -0.787878787879 0 0.4 1e-06 
0.833333333333 -0.787878787879 0 0.4 1e-06 
0.888888888889 -0.787878787879 0 0.4 1e-06 
0.944444444444 -0.787878787879 0 0.4 1e-06 
1.0 -0.787878787879 0 0.4 1e-06 
0.5 -0.747474747475 0 0.4 1e-06 
0.555555555556 -0.747474747475 0 0.4 1e-06 
0.611111111111 -0.747474747475 0 0.4 1e-06 
0.666666666667 -0.747474747475 0 0.4 1e-06 
0.722222222222 -0.747474747475 0 0.4 1e-06 
0.777777777778 -0.747474747475 0 0.4 1e-06 
0.833333333333 -0.747474747475 0 0.4 1e-06 
0.888888888889 -0.747474747475 0 0.4 1e-06 
0.944444444444 -0.747474747475 0 0.4 1e-06 
1.0 -0.747474747475 0 0.4 1e-06 
0.5 -0.707070707071 0 0.4 1e-06 
0.555555555556 -0.707070707071 0 0.4 1e-06 
0.611111111111 -0.707070707071 0 0.4 1e-06 
0.666666666667 -0.707070707071 0 0.4 1e-06 
0.722222222222 -0.707070707071 0 0.4 1e-06 
0.777777777778 -0.707070707071 0 0.4 1e-06 
0.833333333333 -0.707070707071 0 0.4 1e-06 
0.888888888889 -0.707070707071 0 0.4 1e-06 
0.944444444444 -0.707070707071 0 0.4 1e-06 
1.0 -0.707070707071 0 0.4 1e-06 
0.5 -0.666666666667 0 0.4 1e-06 
0.555555555556 -0.666666666667 0 0.4 1e-06 
0.611111111111 -0.666666666667 0 0.4 1e-06 
0.666666666667 -0.666666666667 0 0.4 1e-06 
0.722222222222 -0.666666666667 0 0.4 1e-06 
0.777777777778 -0.666666666667 0 0.4 1e-06 
0.833333333333 -0.666666666667 0 0.4 1e-06 
0.888888888889 -0.666666666667 0 0.4 1e-06 
0.944444444444 -0.666666666667 0 0.4 1e-06 
1.0 -0.666666666667 0 0.4 1e-06 
0.5 -0.626262626263 0 0.4 1e-06 
0.555555555556 -0.626262626263 0 0.4 1e-06 
0.611111111111 -0.626262626263 0 0.4 1e-06 
0.666666666667 -0.626262626263 0 0.4 1e-06 
0.722222222222 -0.626262626263 0 0.4 1e-06 
0.777777777778 -0.626262626263 0 0.4 1e-06 
0.833333333333 -0.626262626263 0 0.4 1e-06 
0.888888888889 -0.626262626263 0 0.4 1e-06 
0.944444444444 -0.626262626263 0 0.4 1e-06 
1.0 -0.626262626263 0 0.4 1e-06 
0.5 -0.585858585859 0 0.4 1e-06 
0.555555555556 -0.585858585859 0 0.4 1e-06 
0.611111111111 -0.585858585859 0 0.4 1e-06 
0.666666666667 -0.585858585859 0 0.4 1e-06 
0.722222222222 -0.585858585859 0 0.4 1e-06 
0.777777777778 -0.585858585859 0 0.4 1e-06 
0.833333333333 -0.585858585859 0 0.4 1e-06 
0.888888888889 -0.585858585859 0 0.4 1e-06 
0.944444444444 -0.585858585859 0 0.4 1e-06 
1.0 -0.585858585859 0 0.4 1e-06 
0.5 -0.545454545455 0 0.4 1e-06 
0.555555555556 -0.545454545455 0 0.4 1e-06 
0.611111111111 -0.545454545455 0 0.4 1e-06 
0.666666666667 -0.545454545455 0 0.4 1e-06 
0.722222222222 -0.545454545455 0 0.4 1e-06 
0.777777777778 -0.545454545455 0 0.4 1e-06 
0.833333333333 -0.545454545455 0 0.4 1e-06 
0.888888888889 -0.545454545455 0 0.4 1e-06 
0.944444444444 -0.545454545455 0 0.4 1e-06 
1.0 -0.545454545455 0 0.4 1e-06 
0.5 -0.505050505051 0 0.4 1e-06 
0.555555555556 -0.505050505051 0 0.4 1e-06 
0.611111111111 -0.505050505051 0 0.4 1e-06 
0.666666666667 -0.505050505051 0 0.4 1e-06 
0.722222222222 -0.505050505051 0 0.4 1e-06 
0.777777777778 -0.505050505051 0 0.4 1e-06 
0.833333333333 -0.505050505051 0 0.4 1e-06 
0.888888888889 -0.505050505051 0 0.4 1e-06 
0.944444444444 -0.505050505051 0 0.4 1e-06 
1.0 -0.505050505051 0 0.4 1e-06 
0.5 -0.464646464646 0 0.4 1e-06 
0.555555555556 -0.464646464646 0 0.4 1e-06 
0.611111111111 -0.464646464646 0 0.4 1e-06 
0.666666666667 -0.464646464646 0 0.4 1e-06 
0.722222222222 -0.464646464646 0 0.4 1e-06 
0.777777777778 -0.464646464646 0 0.4 1e-06 
0.833333333333 -0.464646464646 0 0.4 1e-06 
0.888888888889 -0.464646464646 0 0.4 1e-06 
0.944444444444 -0.464646464646 0 0.4 1e-06 
1.0 -0.464646464646 0 0.4 1e-06 
0.5 -0.424242424242 0 0.4 1e-06 
0.555555555556 -0.424242424242 0 0.4 1e-06 
0.611111111111 -0.424242424242 0 0.4 1e-06 
0.666666666667 -0.424242424242 0 0.4 1e-06 
0.722222222222 -0.424242424242 0 0.4 1e-06 
0.777777777778 -0.424242424242 0 0.4 1e-06 
0.833333333333 -0.424242424242 0 0.4 1e-06 
0.888888888889 -0.424242424242 0 0.4 1e-06 
0.944444444444 -0.424242424242 0 0.4 1e-06 
1.0 -0.424242424242 0 0.4 1e-06 
0.5 -0.383838383838 0 0.4 1e-06 
0.555555555556 -0.383838383838 0 0.4 1e-06 
0.611111111111 -0.383838383838 0 0.4 1e-06 
0.666666666667 -0.383838383838 0 0.4 1e-06 
0.722222222222 -0.383838383838 0 0.4 1e-06 
0.777777777778 -0.383838383838 0 0.4 1e-06 
0.833333333333 -0.383838383838 0 0.4 1e-06 
0.888888888889 -0.383838383838 0 0.4 1e-06 
0.944444444444 -0.383838383838 0 0.4 1e-06 
1.0 -0.383838383838 0 0.4 1e-06 
0.5 -0.343434343434 0 0.4 1e-06 
0.555555555556 -0.343434343434 0 0.4 1e-06 
0.611111111111 -0.343434343434 0 0.4 1e-06 
0.666666666667 -0.343434343434 0 0.4 1e-06 
0.722222222222 -0.343434343434 0 0.4 1e-06 
0.777777777778 -0.343434343434 0 0.4 1e-06 
0.833333333333 -0.343434343434 0 0.4 1e-06 
0.888888888889 -0.343434343434 0 0.4 1e-06 
0.944444444444 -0.343434343434 0 0.4 1e-06 
1.0 -0.343434343434 0 0.4 1e-06 
0.5 -0.30303030303 0 0.4 1e-06 
0.555555555556 -0.30303030303 0 0.4 1e-06 
0.611111111111 -0.30303030303 0 0.4 1e-06 
0.666666666667 -0.30303030303 0 0.4 1e-06 
0.722222222222 -0.30303030303 0 0.4 1e-06 
0.777777777778 -0.30303030303 0 0.4 1e-06 
0.833333333333 -0.30303030303 0 0.4 1e-06 
0.888888888889 -0.30303030303 0 0.4 1e-06 
0.944444444444 -0.30303030303 0 0.4 1e-06 
1.0 -0.30303030303 0 0.4 1e-06 
0.5 -0.262626262626 0 0.4 1e-06 
0.555555555556 -0.262626262626 0 0.4 1e-06 
0.611111111111 -0.262626262626 0 0.4 1e-06 
0.666666666667 -0.262626262626 0 0.4 1e-06 
0.722222222222 -0.262626262626 0 0.4 1e-06 
0.777777777778 -0.262626262626 0 0.4 1e-06 
0.833333333333 -0.262626262626 0 0.4 1e-06 
0.888888888889 -0.262626262626 0 0.4 1e-06 
0.944444444444 -0.262626262626 0 0.4 1e-06 
1.0 -0.262626262626 0 0.4 1e-06 
0.5 -0.222222222222 0 0.4 1e-06 
0.555555555556 -0.222222222222 0 0.4 1e-06 
0.611111111111 -0.222222222222 0 0.4 1e-06 
0.666666666667 -0.222222222222 0 0.4 1e-06 
0.722222222222 -0.222222222222 0 0.4 1e-06 
0.777777777778 -0.222222222222 0 0.4 1e-06 
0.833333333333 -0.222222222222 0 0.4 1e-06 
0.888888888889 -0.222222222222 0 0.4 1e-06 
0.944444444444 -0.222222222222 0 0.4 1e-06 
1.0 -0.222222222222 0 0.4 1e-06 
0.5 -0.181818181818 0 0.4 1e-06 
0.555555555556 -0.181818181818 0 0.4 1e-06 
0.611111111111 -0.181818181818 0 0.4 1e-06 
0.666666666667 -0.181818181818 0 0.4 1e-06 
0.722222222222 -0.181818181818 0 0.4 1e-06 
0.777777777778 -0.181818181818 0 0.4 1e-06 
0.833333333333 -0.181818181818 0 0.4 1e-06 
0.888888888889 -0.181818181818 0 0.4 1e-06 
0.944444444444 -0.181818181818 0 0.4 1e-06 
1.0 -0.181818181818 0 0.4 1e-06 
0.5 -0.141414141414 0 0.4 1e-06 
0.555555555556 -0.141414141414 0 0.4 1e-06 
0.611111111111 -0.141414141414 0 0.4 1e-06 
0.666666666667 -0.141414141414 0 0.4 1e-06 
0.722222222222 -0.141414141414 0 0.4 1e-06 
0.777777777778 -0.141414141414 0 0.4 1e-06 
0.833333333333 -0.141414141414 0 0.4 1e-06 
0.888888888889 -0.141414141414 0 0.4 1e-06 
0.944444444444 -0.141414141414 0 0.4 1e-06 
1.0 -0.141414141414 0 0.4 1e-06 
0.5 -0.10101010101 0 0.4 1e-06 
0.555555555556 -0.10101010101 0 0.4 1e-06 
0.611111111111 -0.10101010101 0 0.4 1e-06 
0.666666666667 -0.10101010101 0 0.4 1e-06 
0.722222222222 -0.10101010101 0 0.4 1e-06 
0.777777777778 -0.10101010101 0 0.4 1e-06 
0.833333333333 -0.10101010101 0 0.4 1e-06 
0.888888888889 -0.10101010101 0 0.4 1e-06 
0.944444444444 -0.10101010101 0 0.4 1e-06 
1.0 -0.10101010101 0 0.4 1e-06 
0.5 -0.0606060606061 0 0.4 1e-06 
0.555555555556 -0.0606060606061 0 0.4 1e-06 
0.611111111111 -0.0606060606061 0 0.4 1e-06 
0.666666666667 -0.0606060606061 0 0.4 1e-06 
0.722222222222 -0.0606060606061 0 0.4 1e-06 
0.777777777778 -0.0606060606061 0 0.4 1e-06 
0.833333333333 -0.0606060606061 0 0.4 1e-06 
0.888888888889 -0.0606060606061 0 0.4 1e-06 
0.944444444444 -0.0606060606061 0 0.4 1e-06 
1.0 -0.0606060606061 0 0.4 1e-06 
0.5 -0.020202020202 0 0.4 1e-06 
0.555555555556 -0.020202020202 0 0.4 1e-06 
0.611111111111 -0.020202020202 0 0.4 1e-06 
0.666666666667 -0.020202020202 0 0.4 1e-06 
0.722222222222 -0.020202020202 0 0.4 1e-06 
0.777777777778 -0.020202020202 0 0.4 1e-06 
0.833333333333 -0.020202020202 0 0.4 1e-06 
0.888888888889 -0.020202020202 0 0.4 1e-06 
0.944444444444 -0.020202020202 0 0.4 1e-06 
1.0 -0.020202020202 0 0.4 1e-06 
0.5 0.020202020202 0 0.4 1e-06 
0.555555555556 0.020202020202 0 0.4 1e-06 
0.611111111111 0.020202020202 0 0.4 1e-06 
0.666666666667 0.020202020202 0 0.4 1e-06 
0.722222222222 0.020202020202 0 0.4 1e-06 
0.777777777778 0.020202020202 0 0.4 1e-06 
0.833333333333 0.020202020202 0 0.4 1e-06 
0.888888888889 0.020202020202 0 0.4 1e-06 
0.944444444444 0.020202020202 0 0.4 1e-06 
1.0 0.020202020202 0 0.4 1e-06 
0.5 0.0606060606061 0 0.4 1e-06 
0.555555555556 0.0606060606061 0 0.4 1e-06 
0.611111111111 0.0606060606061 0 0.4 1e-06 
0.666666666667 0.0606060606061 0 0.4 1e-06 
0.722222222222 0.0606060606061 0 0.4 1e-06 
0.777777777778 0.0606060606061 0 0.4 1e-06 
0.833333333333 0.0606060606061 0 0.4 1e-06 
0.888888888889 0.0606060606061 0 0.4 1e-06 
0.944444444444 0.0606060606061 0 0.4 1e-06 
1.0 0.0606060606061 0 0.4 1e-06 
0.5 0.10101010101 0 0.4 1e-06 
0.555555555556 0.10101010101 0 0.4 1e-06 
0.611111111111 0.10101010101 0 0.4 1e-06 
0.666666666667 0.10101010101 0 0.4 1e-06 
0.722222222222 0.10101010101 0 0.4 1e-06 
0.777777777778 0.10101010101 0 0.4 1e-06 
0.833333333333 0.10101010101 0 0.4 1e-06 
0.888888888889 0.10101010101 0 0.4 1e-06 
0.944444444444 0.10101010101 0 0.4 1e-06 
1.0 0.10101010101 0 0.4 1e-06 
0.5 0.141414141414 0 0.4 1e-06 
0.555555555556 0.141414141414 0 0.4 1e-06 
0.611111111111 0.141414141414 0 0.4 1e-06 
0.666666666667 0.141414141414 0 0.4 1e-06 
0.722222222222 0.141414141414 0 0.4 1e-06 
0.777777777778 0.141414141414 0 0.4 1e-06 
0.833333333333 0.141414141414 0 0.4 1e-06 
0.888888888889 0.141414141414 0 0.4 1e-06 
0.944444444444 0.141414141414 0 0.4 1e-06 
1.0 0.141414141414 0 0.4 1e-06 
0.5 0.181818181818 0 0.4 1e-06 
0.555555555556 0.181818181818 0 0.4 1e-06 
0.611111111111 0.181818181818 0 0.4 1e-06 
0.666666666667 0.181818181818 0 0.4 1e-06 
0.722222222222 0.181818181818 0 0.4 1e-06 
0.777777777778 0.181818181818 0 0.4 1e-06 
0.833333333333 0.181818181818 0 0.4 1e-06 
0.888888888889 0.181818181818 0 0.4 1e-06 
0.944444444444 0.181818181818 0 0.4 1e-06 
1.0 0.181818181818 0 0.4 1e-06 
0.5 0.222222222222 0 0.4 1e-06 
0.555555555556 0.222222222222 0 0.4 1e-06 
0.611111111111 0.222222222222 0 0.4 1e-06 
0.666666666667 0.222222222222 0 0.4 1e-06 
0.722222222222 0.222222222222 0 0.4 1e-06 
0.777777777778 0.222222222222 0 0.4 1e-06 
0.833333333333 0.222222222222 0 0.4 1e-06 
0.888888888889 0.222222222222 0 0.4 1e-06 
0.944444444444 0.222222222222 0 0.4 1e-06 
1.0 0.222222222222 0 0.4 1e-06 
0.5 0.262626262626 0 0.4 1e-06 
0.555555555556 0.262626262626 0 0.4 1e-06 
0.611111111111 0.262626262626 0 0.4 1e-06 
0.666666666667 0.262626262626 0 0.4 1e-06 
0.722222222222 0.262626262626 0 0.4 1e-06 
0.777777777778 0.262626262626 0 0.4 1e-06 
0.833333333333 0.262626262626 0 0.4 1e-06 
0.888888888889 0.262626262626 0 0.4 1e-06 
0.944444444444 0.262626262626 0 0.4 1e-06 
1.0 0.262626262626 0 0.4 1e-06 
0.5 0.30303030303 0 0.4 1e-06 
0.555555555556 0.30303030303 0 0.4 1e-06 
0.611111111111 0.30303030303 0 0.4 1e-06 
0.666666666667 0.30303030303 0 0.4 1e-06 
0.722222222222 0.30303030303 0 0.4 1e-06 
0.777777777778 0.30303030303 0 0.4 1e-06 
0.833333333333 0.30303030303 0 0.4 1e-06 
0.888888888889 0.30303030303 0 0.4 1e-06 
0.944444444444 0.30303030303 0 0.4 1e-06 
1.0 0.30303030303 0 0.4 1e-06 
0.5 0.343434343434 0 0.4 1e-06 
0.555555555556 0.343434343434 0 0.4 1e-06 
0.611111111111 0.343434343434 0 0.4 1e-06 
0.666666666667 0.343434343434 0 0.4 1e-06 
0.722222222222 0.343434343434 0 0.4 1e-06 
0.777777777778 0.343434343434 0 0.4 1e-06 
0.833333333333 0.343434343434 0 0.4 1e-06 
0.888888888889 0.343434343434 0 0.4 1e-06 
0.944444444444 0.343434343434 0 0.4 1e-06 
1.0 0.343434343434 0 0.4 1e-06 
0.5 0.383838383838 0 0.4 1e-06 
0.555555555556 0.383838383838 0 0.4 1e-06 
0.611111111111 0.383838383838 0 0.4 1e-06 
0.666666666667 0.383838383838 0 0.4 1e-06 
0.722222222222 0.383838383838 0 0.4 1e-06 
0.777777777778 0.383838383838 0 0.4 1e-06 
0.833333333333 0.383838383838 0 0.4 1e-06 
0.888888888889 0.383838383838 0 0.4 1e-06 
0.944444444444 0.383838383838 0 0.4 1e-06 
1.0 0.383838383838 0 0.4 1e-06 
0.5 0.424242424242 0 0.4 1e-06 
0.555555555556 0.424242424242 0 0.4 1e-06 
0.611111111111 0.424242424242 0 0.4 1e-06 
0.666666666667 0.424242424242 0 0.4 1e-06 
0.722222222222 0.424242424242 0 0.4 1e-06 
0.777777777778 0.424242424242 0 0.4 1e-06 
0.833333333333 0.424242424242 0 0.4 1e-06 
0.888888888889 0.424242424242 0 0.4 1e-06 
0.944444444444 0.424242424242 0 0.4 1e-06 
1.0 0.424242424242 0 0.4 1e-06 
0.5 0.464646464646 0 0.4 1e-06 
0.555555555556 0.464646464646 0 0.4 1e-06 
0.611111111111 0.464646464646 0 0.4 1e-06 
0.666666666667 0.464646464646 0 0.4 1e-06 
0.722222222222 0.464646464646 0 0.4 1e-06 
0.777777777778 0.464646464646 0 0.4 1e-06 
0.833333333333 0.464646464646 0 0.4 1e-06 
0.888888888889 0.464646464646 0 0.4 1e-06 
0.944444444444 0.464646464646 0 0.4 1e-06 
1.0 0.464646464646 0 0.4 1e-06 
0.5 0.505050505051 0 0.4 1e-06 
0.555555555556 0.505050505051 0 0.4 1e-06 
0.611111111111 0.505050505051 0 0.4 1e-06 
0.666666666667 0.505050505051 0 0.4 1e-06 
0.722222222222 0.505050505051 0 0.4 1e-06 
0.777777777778 0.505050505051 0 0.4 1e-06 
0.833333333333 0.505050505051 0 0.4 1e-06 
0.888888888889 0.505050505051 0 0.4 1e-06 
0.944444444444 0.505050505051 0 0.4 1e-06 
1.0 0.505050505051 0 0.4 1e-06 
0.5 0.545454545455 0 0.4 1e-06 
0.555555555556 0.545454545455 0 0.4 1e-06 
0.611111111111 0.545454545455 0 0.4 1e-06 
0.666666666667 0.545454545455 0 0.4 1e-06 
0.722222222222 0.545454545455 0 0.4 1e-06 
0.777777777778 0.545454545455 0 0.4 1e-06 
0.833333333333 0.545454545455 0 0.4 1e-06 
0.888888888889 0.545454545455 0 0.4 1e-06 
0.944444444444 0.545454545455 0 0.4 1e-06 
1.0 0.545454545455 0 0.4 1e-06 
0.5 0.585858585859 0 0.4 1e-06 
0.555555555556 0.585858585859 0 0.4 1e-06 
0.611111111111 0.585858585859 0 0.4 1e-06 
0.666666666667 0.585858585859 0 0.4 1e-06 
0.722222222222 0.585858585859 0 0.4 1e-06 
0.777777777778 0.585858585859 0 0.4 1e-06 
0.833333333333 0.585858585859 0 0.4 1e-06 
0.888888888889 0.585858585859 0 0.4 1e-06 
0.944444444444 0.585858585859 0 0.4 1e-06 
1.0 0.585858585859 0 0.4 1e-06 
0.5 0.626262626263 0 0.4 1e-06 
0.555555555556 0.626262626263 0 0.4 1e-06 
0.611111111111 0.626262626263 0 0.4 1e-06 
0.666666666667 0.626262626263 0 0.4 1e-06 
0.722222222222 0.626262626263 0 0.4 1e-06 
0.777777777778 0.626262626263 0 0.4 1e-06 
0.833333333333 0.626262626263 0 0.4 1e-06 
0.888888888889 0.626262626263 0 0.4 1e-06 
0.944444444444 0.626262626263 0 0.4 1e-06 
1.0 0.626262626263 0 0.4 1e-06 
0.5 0.666666666667 0 0.4 1e-06 
0.555555555556 0.666666666667 0 0.4 1e-06 
0.611111111111 0.666666666667 0 0.4 1e-06 
0.666666666667 0.666666666667 0 0.4 1e-06 
0.722222222222 0.666666666667 0 0.4 1e-06 
0.777777777778 0.666666666667 0 0.4 1e-06 
0.833333333333 0.666666666667 0 0.4 1e-06 
0.888888888889 0.666666666667 0 0.4 1e-06 
0.944444444444 0.666666666667 0 0.4 1e-06 
1.0 0.666666666667 0 0.4 1e-06 
0.5 0.707070707071 0 0.4 1e-06 
0.555555555556 0.707070707071 0 0.4 1e-06 
0.611111111111 0.707070707071 0 0.4 1e-06 
0.666666666667 0.707070707071 0 0.4 1e-06 
0.722222222222 0.707070707071 0 0.4 1e-06 
0.777777777778 0.707070707071 0 0.4 1e-06 
0.833333333333 0.707070707071 0 0.4 1e-06 
0.888888888889 0.707070707071 0 0.4 1e-06 
0.944444444444 0.707070707071 0 0.4 1e-06 
1.0 0.707070707071 0 0.4 1e-06 
0.5 0.747474747475 0 0.4 1e-06 
0.555555555556 0.747474747475 0 0.4 1e-06 
0.611111111111 0.747474747475 0 0.4 1e-06 
0.666666666667 0.747474747475 0 0.4 1e-06 
0.722222222222 0.747474747475 0 0.4 1e-06 
0.777777777778 0.747474747475 0 0.4 1e-06 
0.833333333333 0.747474747475 0 0.4 1e-06 
0.888888888889 0.747474747475 0 0.4 1e-06 
0.944444444444 0.747474747475 0 0.4 1e-06 
1.0 0.747474747475 0 0.4 1e-06 
0.5 0.787878787879 0 0.4 1e-06 
0.555555555556 0.787878787879 0 0.4 1e-06 
0.611111111111 0.787878787879 0 0.4 1e-06 
0.666666666667 0.787878787879 0 0.4 1e-06 
0.722222222222 0.787878787879 0 0.4 1e-06 
0.777777777778 0.787878787879 0 0.4 1e-06 
0.833333333333 0.787878787879 0 0.4 1e-06 
0.888888888889 0.787878787879 0 0.4 1e-06 
0.944444444444 0.787878787879 0 0.4 1e-06 
1.0 0.787878787879 0 0.4 1e-06 
0.5 0.828282828283 0 0.4 1e-06 
0.555555555556 0.828282828283 0 0.4 1e-06 
0.611111111111 0.828282828283 0 0.4 1e-06 
0.666666666667 0.828282828283 0 0.4 1e-06 
0.722222222222 0.828282828283 0 0.4 1e-06 
0.777777777778 0.828282828283 0 0.4 1e-06 
0.833333333333 0.828282828283 0 0.4 1e-06 
0.888888888889 0.828282828283 0 0.4 1e-06 
0.944444444444 0.828282828283 0 0.4 1e-06 
1.0 0.828282828283 0 0.4 1e-06 
0.5 0.868686868687 0 0.4 1e-06 
0.555555555556 0.868686868687 0 0.4 1e-06 
0.611111111111 0.868686868687 0 0.4 1e-06 
0.666666666667 0.868686868687 0 0.4 1e-06 
0.722222222222 0.868686868687 0 0.4 1e-06 
0.777777777778 0.868686868687 0 0.4 1e-06 
0.833333333333 0.868686868687 0 0.4 1e-06 
0.888888888889 0.868686868687 0 0.4 1e-06 
0.944444444444 0.868686868687 0 0.4 1e-06 
1.0 0.868686868687 0 0.4 1e-06 
0.5 0.909090909091 0 0.4 1e-06 
0.555555555556 0.909090909091 0 0.4 1e-06 
0.611111111111 0.909090909091 0 0.4 1e-06 
0.666666666667 0.909090909091 0 0.4 1e-06 
0.722222222222 0.909090909091 0 0.4 1e-06 
0.777777777778 0.909090909091 0 0.4 1e-06 
0.833333333333 0.909090909091 0 0.4 1e-06 
0.888888888889 0.909090909091 0 0.4 1e-06 
0.944444444444 0.909090909091 0 0.4 1e-06 
1.0 0.909090909091 0 0.4 1e-06 
0.5 0.949494949495 0 0.4 1e-06 
0.555555555556 0.949494949495 0 0.4 1e-06 
0.611111111111 0.949494949495 0 0.4 1e-06 
0.666666666667 0.949494949495 0 0.4 1e-06 
0.722222222222 0.949494949495 0 0.4 1e-06 
0.777777777778 0.949494949495 0 0.4 1e-06 
0.833333333333 0.949494949495 0 0.4 1e-06 
0.888888888889 0.949494949495 0 0.4 1e-06 
0.944444444444 0.949494949495 0 0.4 1e-06 
1.0 0.949494949495 0 0.4 1e-06 
0.5 0.989898989899 0 0.4 1e-06 
0.555555555556 0.989898989899 0 0.4 1e-06 
0.611111111111 0.989898989899 0 0.4 1e-06 
0.666666666667 0.989898989899 0 0.4 1e-06 
0.722222222222 0.989898989899 0 0.4 1e-06 
0.777777777778 0.989898989899 0 0.4 1e-06 
0.833333333333 0.989898989899 0 0.4 1e-06 
0.888888888889 0.989898989899 0 0.4 1e-06 
0.944444444444 0.989898989899 0 0.4 1e-06 
1.0 0.989898989899 0 0.4 1e-06 
0.5 1.0303030303 0 0.4 1e-06 
0.555555555556 1.0303030303 0 0.4 1e-06 
0.611111111111 1.0303030303 0 0.4 1e-06 
0.666666666667 1.0303030303 0 0.4 1e-06 
0.722222222222 1.0303030303 0 0.4 1e-06 
0.777777777778 1.0303030303 0 0.4 1e-06 
0.833333333333 1.0303030303 0 0.4 1e-06 
0.888888888889 1.0303030303 0 0.4 1e-06 
0.944444444444 1.0303030303 0 0.4 1e-06 
1.0 1.0303030303 0 0.4 1e-06 
0.5 1.07070707071 0 0.4 1e-06 
0.555555555556 1.07070707071 0 0.4 1e-06 
0.611111111111 1.07070707071 0 0.4 1e-06 
0.666666666667 1.07070707071 0 0.4 1e-06 
0.722222222222 1.07070707071 0 0.4 1e-06 
0.777777777778 1.07070707071 0 0.4 1e-06 
0.833333333333 1.07070707071 0 0.4 1e-06 
0.888888888889 1.07070707071 0 0.4 1e-06 
0.944444444444 1.07070707071 0 0.4 1e-06 
1.0 1.07070707071 0 0.4 1e-06 
0.5 1.11111111111 0 0.4 1e-06 
0.555555555556 1.11111111111 0 0.4 1e-06 
0.611111111111 1.11111111111 0 0.4 1e-06 
0.666666666667 1.11111111111 0 0.4 1e-06 
0.722222222222 1.11111111111 0 0.4 1e-06 
0.777777777778 1.11111111111 0 0.4 1e-06 
0.833333333333 1.11111111111 0 0.4 1e-06 
0.888888888889 1.11111111111 0 0.4 1e-06 
0.944444444444 1.11111111111 0 0.4 1e-06 
1.0 1.11111111111 0 0.4 1e-06 
0.5 1.15151515152 0 0.4 1e-06 
0.555555555556 1.15151515152 0 0.4 1e-06 
0.611111111111 1.15151515152 0 0.4 1e-06 
0.666666666667 1.15151515152 0 0.4 1e-06 
0.722222222222 1.15151515152 0 0.4 1e-06 
0.777777777778 1.15151515152 0 0.4 1e-06 
0.833333333333 1.15151515152 0 0.4 1e-06 
0.888888888889 1.15151515152 0 0.4 1e-06 
0.944444444444 1.15151515152 0 0.4 1e-06 
1.0 1.15151515152 0 0.4 1e-06 
0.5 1.19191919192 0 0.4 1e-06 
0.555555555556 1.19191919192 0 0.4 1e-06 
0.611111111111 1.19191919192 0 0.4 1e-06 
0.666666666667 1.19191919192 0 0.4 1e-06 
0.722222222222 1.19191919192 0 0.4 1e-06 
0.777777777778 1.19191919192 0 0.4 1e-06 
0.833333333333 1.19191919192 0 0.4 1e-06 
0.888888888889 1.19191919192 0 0.4 1e-06 
0.944444444444 1.19191919192 0 0.4 1e-06 
1.0 1.19191919192 0 0.4 1e-06 
0.5 1.23232323232 0 0.4 1e-06 
0.555555555556 1.23232323232 0 0.4 1e-06 
0.611111111111 1.23232323232 0 0.4 1e-06 
0.666666666667 1.23232323232 0 0.4 1e-06 
0.722222222222 1.23232323232 0 0.4 1e-06 
0.777777777778 1.23232323232 0 0.4 1e-06 
0.833333333333 1.23232323232 0 0.4 1e-06 
0.888888888889 1.23232323232 0 0.4 1e-06 
0.944444444444 1.23232323232 0 0.4 1e-06 
1.0 1.23232323232 0 0.4 1e-06 
0.5 1.27272727273 0 0.4 1e-06 
0.555555555556 1.27272727273 0 0.4 1e-06 
0.611111111111 1.27272727273 0 0.4 1e-06 
0.666666666667 1.27272727273 0 0.4 1e-06 
0.722222222222 1.27272727273 0 0.4 1e-06 
0.777777777778 1.27272727273 0 0.4 1e-06 
0.833333333333 1.27272727273 0 0.4 1e-06 
0.888888888889 1.27272727273 0 0.4 1e-06 
0.944444444444 1.27272727273 0 0.4 1e-06 
1.0 1.27272727273 0 0.4 1e-06 
0.5 1.31313131313 0 0.4 1e-06 
0.555555555556 1.31313131313 0 0.4 1e-06 
0.611111111111 1.31313131313 0 0.4 1e-06 
0.666666666667 1.31313131313 0 0.4 1e-06 
0.722222222222 1.31313131313 0 0.4 1e-06 
0.777777777778 1.31313131313 0 0.4 1e-06 
0.833333333333 1.31313131313 0 0.4 1e-06 
0.888888888889 1.31313131313 0 0.4 1e-06 
0.944444444444 1.31313131313 0 0.4 1e-06 
1.0 1.31313131313 0 0.4 1e-06 
0.5 1.35353535354 0 0.4 1e-06 
0.555555555556 1.35353535354 0 0.4 1e-06 
0.611111111111 1.35353535354 0 0.4 1e-06 
0.666666666667 1.35353535354 0 0.4 1e-06 
0.722222222222 1.35353535354 0 0.4 1e-06 
0.777777777778 1.35353535354 0 0.4 1e-06 
0.833333333333 1.35353535354 0 0.4 1e-06 
0.888888888889 1.35353535354 0 0.4 1e-06 
0.944444444444 1.35353535354 0 0.4 1e-06 
1.0 1.35353535354 0 0.4 1e-06 
0.5 1.39393939394 0 0.4 1e-06 
0.555555555556 1.39393939394 0 0.4 1e-06 
0.611111111111 1.39393939394 0 0.4 1e-06 
0.666666666667 1.39393939394 0 0.4 1e-06 
0.722222222222 1.39393939394 0 0.4 1e-06 
0.777777777778 1.39393939394 0 0.4 1e-06 
0.833333333333 1.39393939394 0 0.4 1e-06 
0.888888888889 1.39393939394 0 0.4 1e-06 
0.944444444444 1.39393939394 0 0.4 1e-06 
1.0 1.39393939394 0 0.4 1e-06 
0.5 1.43434343434 0 0.4 1e-06 
0.555555555556 1.43434343434 0 0.4 1e-06 
0.611111111111 1.43434343434 0 0.4 1e-06 
0.666666666667 1.43434343434 0 0.4 1e-06 
0.722222222222 1.43434343434 0 0.4 1e-06 
0.777777777778 1.43434343434 0 0.4 1e-06 
0.833333333333 1.43434343434 0 0.4 1e-06 
0.888888888889 1.43434343434 0 0.4 1e-06 
0.944444444444 1.43434343434 0 0.4 1e-06 
1.0 1.43434343434 0 0.4 1e-06 
0.5 1.47474747475 0 0.4 1e-06 
0.555555555556 1.47474747475 0 0.4 1e-06 
0.611111111111 1.47474747475 0 0.4 1e-06 
0.666666666667 1.47474747475 0 0.4 1e-06 
0.722222222222 1.47474747475 0 0.4 1e-06 
0.777777777778 1.47474747475 0 0.4 1e-06 
0.833333333333 1.47474747475 0 0.4 1e-06 
0.888888888889 1.47474747475 0 0.4 1e-06 
0.944444444444 1.47474747475 0 0.4 1e-06 
1.0 1.47474747475 0 0.4 1e-06 
0.5 1.51515151515 0 0.4 1e-06 
0.555555555556 1.51515151515 0 0.4 1e-06 
0.611111111111 1.51515151515 0 0.4 1e-06 
0.666666666667 1.51515151515 0 0.4 1e-06 
0.722222222222 1.51515151515 0 0.4 1e-06 
0.777777777778 1.51515151515 0 0.4 1e-06 
0.833333333333 1.51515151515 0 0.4 1e-06 
0.888888888889 1.51515151515 0 0.4 1e-06 
0.944444444444 1.51515151515 0 0.4 1e-06 
1.0 1.51515151515 0 0.4 1e-06 
0.5 1.55555555556 0 0.4 1e-06 
0.555555555556 1.55555555556 0 0.4 1e-06 
0.611111111111 1.55555555556 0 0.4 1e-06 
0.666666666667 1.55555555556 0 0.4 1e-06 
0.722222222222 1.55555555556 0 0.4 1e-06 
0.777777777778 1.55555555556 0 0.4 1e-06 
0.833333333333 1.55555555556 0 0.4 1e-06 
0.888888888889 1.55555555556 0 0.4 1e-06 
0.944444444444 1.55555555556 0 0.4 1e-06 
1.0 1.55555555556 0 0.4 1e-06 
0.5 1.59595959596 0 0.4 1e-06 
0.555555555556 1.59595959596 0 0.4 1e-06 
0.611111111111 1.59595959596 0 0.4 1e-06 
0.666666666667 1.59595959596 0 0.4 1e-06 
0.722222222222 1.59595959596 0 0.4 1e-06 
0.777777777778 1.59595959596 0 0.4 1e-06 
0.833333333333 1.59595959596 0 0.4 1e-06 
0.888888888889 1.59595959596 0 0.4 1e-06 
0.944444444444 1.59595959596 0 0.4 1e-06 
1.0 1.59595959596 0 0.4 1e-06 
0.5 1.63636363636 0 0.4 1e-06 
0.555555555556 1.63636363636 0 0.4 1e-06 
0.611111111111 1.63636363636 0 0.4 1e-06 
0.666666666667 1.63636363636 0 0.4 1e-06 
0.722222222222 1.63636363636 0 0.4 1e-06 
0.777777777778 1.63636363636 0 0.4 1e-06 
0.833333333333 1.63636363636 0 0.4 1e-06 
0.888888888889 1.63636363636 0 0.4 1e-06 
0.944444444444 1.63636363636 0 0.4 1e-06 
1.0 1.63636363636 0 0.4 1e-06 
0.5 1.67676767677 0 0.4 1e-06 
0.555555555556 1.67676767677 0 0.4 1e-06 
0.611111111111 1.67676767677 0 0.4 1e-06 
0.666666666667 1.67676767677 0 0.4 1e-06 
0.722222222222 1.67676767677 0 0.4 1e-06 
0.777777777778 1.67676767677 0 0.4 1e-06 
0.833333333333 1.67676767677 0 0.4 1e-06 
0.888888888889 1.67676767677 0 0.4 1e-06 
0.944444444444 1.67676767677 0 0.4 1e-06 
1.0 1.67676767677 0 0.4 1e-06 
0.5 1.71717171717 0 0.4 1e-06 
0.555555555556 1.71717171717 0 0.4 1e-06 
0.611111111111 1.71717171717 0 0.4 1e-06 
0.666666666667 1.71717171717 0 0.4 1e-06 
0.722222222222 1.71717171717 0 0.4 1e-06 
0.777777777778 1.71717171717 0 0.4 1e-06 
0.833333333333 1.71717171717 0 0.4 1e-06 
0.888888888889 1.71717171717 0 0.4 1e-06 
0.944444444444 1.71717171717 0 0.4 1e-06 
1.0 1.71717171717 0 0.4 1e-06 
0.5 1.75757575758 0 0.4 1e-06 
0.555555555556 1.75757575758 0 0.4 1e-06 
0.611111111111 1.75757575758 0 0.4 1e-06 
0.666666666667 1.75757575758 0 0.4 1e-06 
0.722222222222 1.75757575758 0 0.4 1e-06 
0.777777777778 1.75757575758 0 0.4 1e-06 
0.833333333333 1.75757575758 0 0.4 1e-06 
0.888888888889 1.75757575758 0 0.4 1e-06 
0.944444444444 1.75757575758 0 0.4 1e-06 
1.0 1.75757575758 0 0.4 1e-06 
0.5 1.79797979798 0 0.4 1e-06 
0.555555555556 1.79797979798 0 0.4 1e-06 
0.611111111111 1.79797979798 0 0.4 1e-06 
0.666666666667 1.79797979798 0 0.4 1e-06 
0.722222222222 1.79797979798 0 0.4 1e-06 
0.777777777778 1.79797979798 0 0.4 1e-06 
0.833333333333 1.79797979798 0 0.4 1e-06 
0.888888888889 1.79797979798 0 0.4 1e-06 
0.944444444444 1.79797979798 0 0.4 1e-06 
1.0 1.79797979798 0 0.4 1e-06 
0.5 1.83838383838 0 0.4 1e-06 
0.555555555556 1.83838383838 0 0.4 1e-06 
0.611111111111 1.83838383838 0 0.4 1e-06 
0.666666666667 1.83838383838 0 0.4 1e-06 
0.722222222222 1.83838383838 0 0.4 1e-06 
0.777777777778 1.83838383838 0 0.4 1e-06 
0.833333333333 1.83838383838 0 0.4 1e-06 
0.888888888889 1.83838383838 0 0.4 1e-06 
0.944444444444 1.83838383838 0 0.4 1e-06 
1.0 1.83838383838 0 0.4 1e-06 
0.5 1.87878787879 0 0.4 1e-06 
0.555555555556 1.87878787879 0 0.4 1e-06 
0.611111111111 1.87878787879 0 0.4 1e-06 
0.666666666667 1.87878787879 0 0.4 1e-06 
0.722222222222 1.87878787879 0 0.4 1e-06 
0.777777777778 1.87878787879 0 0.4 1e-06 
0.833333333333 1.87878787879 0 0.4 1e-06 
0.888888888889 1.87878787879 0 0.4 1e-06 
0.944444444444 1.87878787879 0 0.4 1e-06 
1.0 1.87878787879 0 0.4 1e-06 
0.5 1.91919191919 0 0.4 1e-06 
0.555555555556 1.91919191919 0 0.4 1e-06 
0.611111111111 1.91919191919 0 0.4 1e-06 
0.666666666667 1.91919191919 0 0.4 1e-06 
0.722222222222 1.91919191919 0 0.4 1e-06 
0.777777777778 1.91919191919 0 0.4 1e-06 
0.833333333333 1.91919191919 0 0.4 1e-06 
0.888888888889 1.91919191919 0 0.4 1e-06 
0.944444444444 1.91919191919 0 0.4 1e-06 
1.0 1.91919191919 0 0.4 1e-06 
0.5 1.9595959596 0 0.4 1e-06 
0.555555555556 1.9595959596 0 0.4 1e-06 
0.611111111111 1.9595959596 0 0.4 1e-06 
0.666666666667 1.9595959596 0 0.4 1e-06 
0.722222222222 1.9595959596 0 0.4 1e-06 
0.777777777778 1.9595959596 0 0.4 1e-06 
0.833333333333 1.9595959596 0 0.4 1e-06 
0.888888888889 1.9595959596 0 0.4 1e-06 
0.944444444444 1.9595959596 0 0.4 1e-06 
1.0 1.9595959596 0 0.4 1e-06 
0.5 2.0 0 0.4 1e-06 
0.555555555556 2.0 0 0.4 1e-06 
0.611111111111 2.0 0 0.4 1e-06 
0.666666666667 2.0 0 0.4 1e-06 
0.722222222222 2.0 0 0.4 1e-06 
0.777777777778 2.0 0 0.4 1e-06 
0.833333333333 2.0 0 0.4 1e-06 
0.888888888889 2.0 0 0.4 1e-06 
0.944444444444 2.0 0 0.4 1e-06 
1.0 2.0 0 0.4 1e-06 
0.5 -2.0 0 0.8 1e-06 
0.555555555556 -2.0 0 0.8 1e-06 
0.611111111111 -2.0 0 0.8 1e-06 
0.666666666667 -2.0 0 0.8 1e-06 
0.722222222222 -2.0 0 0.8 1e-06 
0.777777777778 -2.0 0 0.8 1e-06 
0.833333333333 -2.0 0 0.8 1e-06 
0.888888888889 -2.0 0 0.8 1e-06 
0.944444444444 -2.0 0 0.8 1e-06 
1.0 -2.0 0 0.8 1e-06 
0.5 -1.9595959596 0 0.8 1e-06 
0.555555555556 -1.9595959596 0 0.8 1e-06 
0.611111111111 -1.9595959596 0 0.8 1e-06 
0.666666666667 -1.9595959596 0 0.8 1e-06 
0.722222222222 -1.9595959596 0 0.8 1e-06 
0.777777777778 -1.9595959596 0 0.8 1e-06 
0.833333333333 -1.9595959596 0 0.8 1e-06 
0.888888888889 -1.9595959596 0 0.8 1e-06 
0.944444444444 -1.9595959596 0 0.8 1e-06 
1.0 -1.9595959596 0 0.8 1e-06 
0.5 -1.91919191919 0 0.8 1e-06 
0.555555555556 -1.91919191919 0 0.8 1e-06 
0.611111111111 -1.91919191919 0 0.8 1e-06 
0.666666666667 -1.91919191919 0 0.8 1e-06 
0.722222222222 -1.91919191919 0 0.8 1e-06 
0.777777777778 -1.91919191919 0 0.8 1e-06 
0.833333333333 -1.91919191919 0 0.8 1e-06 
0.888888888889 -1.91919191919 0 0.8 1e-06 
0.944444444444 -1.91919191919 0 0.8 1e-06 
1.0 -1.91919191919 0 0.8 1e-06 
0.5 -1.87878787879 0 0.8 1e-06 
0.555555555556 -1.87878787879 0 0.8 1e-06 
0.611111111111 -1.87878787879 0 0.8 1e-06 
0.666666666667 -1.87878787879 0 0.8 1e-06 
0.722222222222 -1.87878787879 0 0.8 1e-06 
0.777777777778 -1.87878787879 0 0.8 1e-06 
0.833333333333 -1.87878787879 0 0.8 1e-06 
0.888888888889 -1.87878787879 0 0.8 1e-06 
0.944444444444 -1.87878787879 0 0.8 1e-06 
1.0 -1.87878787879 0 0.8 1e-06 
0.5 -1.83838383838 0 0.8 1e-06 
0.555555555556 -1.83838383838 0 0.8 1e-06 
0.611111111111 -1.83838383838 0 0.8 1e-06 
0.666666666667 -1.83838383838 0 0.8 1e-06 
0.722222222222 -1.83838383838 0 0.8 1e-06 
0.777777777778 -1.83838383838 0 0.8 1e-06 
0.833333333333 -1.83838383838 0 0.8 1e-06 
0.888888888889 -1.83838383838 0 0.8 1e-06 
0.944444444444 -1.83838383838 0 0.8 1e-06 
1.0 -1.83838383838 0 0.8 1e-06 
0.5 -1.79797979798 0 0.8 1e-06 
0.555555555556 -1.79797979798 0 0.8 1e-06 
0.611111111111 -1.79797979798 0 0.8 1e-06 
0.666666666667 -1.79797979798 0 0.8 1e-06 
0.722222222222 -1.79797979798 0 0.8 1e-06 
0.777777777778 -1.79797979798 0 0.8 1e-06 
0.833333333333 -1.79797979798 0 0.8 1e-06 
0.888888888889 -1.79797979798 0 0.8 1e-06 
0.944444444444 -1.79797979798 0 0.8 1e-06 
1.0 -1.79797979798 0 0.8 1e-06 
0.5 -1.75757575758 0 0.8 1e-06 
0.555555555556 -1.75757575758 0 0.8 1e-06 
0.611111111111 -1.75757575758 0 0.8 1e-06 
0.666666666667 -1.75757575758 0 0.8 1e-06 
0.722222222222 -1.75757575758 0 0.8 1e-06 
0.777777777778 -1.75757575758 0 0.8 1e-06 
0.833333333333 -1.75757575758 0 0.8 1e-06 
0.888888888889 -1.75757575758 0 0.8 1e-06 
0.944444444444 -1.75757575758 0 0.8 1e-06 
1.0 -1.75757575758 0 0.8 1e-06 
0.5 -1.71717171717 0 0.8 1e-06 
0.555555555556 -1.71717171717 0 0.8 1e-06 
0.611111111111 -1.71717171717 0 0.8 1e-06 
0.666666666667 -1.71717171717 0 0.8 1e-06 
0.722222222222 -1.71717171717 0 0.8 1e-06 
0.777777777778 -1.71717171717 0 0.8 1e-06 
0.833333333333 -1.71717171717 0 0.8 1e-06 
0.888888888889 -1.71717171717 0 0.8 1e-06 
0.944444444444 -1.71717171717 0 0.8 1e-06 
1.0 -1.71717171717 0 0.8 1e-06 
0.5 -1.67676767677 0 0.8 1e-06 
0.555555555556 -1.67676767677 0 0.8 1e-06 
0.611111111111 -1.67676767677 0 0.8 1e-06 
0.666666666667 -1.67676767677 0 0.8 1e-06 
0.722222222222 -1.67676767677 0 0.8 1e-06 
0.777777777778 -1.67676767677 0 0.8 1e-06 
0.833333333333 -1.67676767677 0 0.8 1e-06 
0.888888888889 -1.67676767677 0 0.8 1e-06 
0.944444444444 -1.67676767677 0 0.8 1e-06 
1.0 -1.67676767677 0 0.8 1e-06 
0.5 -1.63636363636 0 0.8 1e-06 
0.555555555556 -1.63636363636 0 0.8 1e-06 
0.611111111111 -1.63636363636 0 0.8 1e-06 
0.666666666667 -1.63636363636 0 0.8 1e-06 
0.722222222222 -1.63636363636 0 0.8 1e-06 
0.777777777778 -1.63636363636 0 0.8 1e-06 
0.833333333333 -1.63636363636 0 0.8 1e-06 
0.888888888889 -1.63636363636 0 0.8 1e-06 
0.944444444444 -1.63636363636 0 0.8 1e-06 
1.0 -1.63636363636 0 0.8 1e-06 
0.5 -1.59595959596 0 0.8 1e-06 
0.555555555556 -1.59595959596 0 0.8 1e-06 
0.611111111111 -1.59595959596 0 0.8 1e-06 
0.666666666667 -1.59595959596 0 0.8 1e-06 
0.722222222222 -1.59595959596 0 0.8 1e-06 
0.777777777778 -1.59595959596 0 0.8 1e-06 
0.833333333333 -1.59595959596 0 0.8 1e-06 
0.888888888889 -1.59595959596 0 0.8 1e-06 
0.944444444444 -1.59595959596 0 0.8 1e-06 
1.0 -1.59595959596 0 0.8 1e-06 
0.5 -1.55555555556 0 0.8 1e-06 
0.555555555556 -1.55555555556 0 0.8 1e-06 
0.611111111111 -1.55555555556 0 0.8 1e-06 
0.666666666667 -1.55555555556 0 0.8 1e-06 
0.722222222222 -1.55555555556 0 0.8 1e-06 
0.777777777778 -1.55555555556 0 0.8 1e-06 
0.833333333333 -1.55555555556 0 0.8 1e-06 
0.888888888889 -1.55555555556 0 0.8 1e-06 
0.944444444444 -1.55555555556 0 0.8 1e-06 
1.0 -1.55555555556 0 0.8 1e-06 
0.5 -1.51515151515 0 0.8 1e-06 
0.555555555556 -1.51515151515 0 0.8 1e-06 
0.611111111111 -1.51515151515 0 0.8 1e-06 
0.666666666667 -1.51515151515 0 0.8 1e-06 
0.722222222222 -1.51515151515 0 0.8 1e-06 
0.777777777778 -1.51515151515 0 0.8 1e-06 
0.833333333333 -1.51515151515 0 0.8 1e-06 
0.888888888889 -1.51515151515 0 0.8 1e-06 
0.944444444444 -1.51515151515 0 0.8 1e-06 
1.0 -1.51515151515 0 0.8 1e-06 
0.5 -1.47474747475 0 0.8 1e-06 
0.555555555556 -1.47474747475 0 0.8 1e-06 
0.611111111111 -1.47474747475 0 0.8 1e-06 
0.666666666667 -1.47474747475 0 0.8 1e-06 
0.722222222222 -1.47474747475 0 0.8 1e-06 
0.777777777778 -1.47474747475 0 0.8 1e-06 
0.833333333333 -1.47474747475 0 0.8 1e-06 
0.888888888889 -1.47474747475 0 0.8 1e-06 
0.944444444444 -1.47474747475 0 0.8 1e-06 
1.0 -1.47474747475 0 0.8 1e-06 
0.5 -1.43434343434 0 0.8 1e-06 
0.555555555556 -1.43434343434 0 0.8 1e-06 
0.611111111111 -1.43434343434 0 0.8 1e-06 
0.666666666667 -1.43434343434 0 0.8 1e-06 
0.722222222222 -1.43434343434 0 0.8 1e-06 
0.777777777778 -1.43434343434 0 0.8 1e-06 
0.833333333333 -1.43434343434 0 0.8 1e-06 
0.888888888889 -1.43434343434 0 0.8 1e-06 
0.944444444444 -1.43434343434 0 0.8 1e-06 
1.0 -1.43434343434 0 0.8 1e-06 
0.5 -1.39393939394 0 0.8 1e-06 
0.555555555556 -1.39393939394 0 0.8 1e-06 
0.611111111111 -1.39393939394 0 0.8 1e-06 
0.666666666667 -1.39393939394 0 0.8 1e-06 
0.722222222222 -1.39393939394 0 0.8 1e-06 
0.777777777778 -1.39393939394 0 0.8 1e-06 
0.833333333333 -1.39393939394 0 0.8 1e-06 
0.888888888889 -1.39393939394 0 0.8 1e-06 
0.944444444444 -1.39393939394 0 0.8 1e-06 
1.0 -1.39393939394 0 0.8 1e-06 
0.5 -1.35353535354 0 0.8 1e-06 
0.555555555556 -1.35353535354 0 0.8 1e-06 
0.611111111111 -1.35353535354 0 0.8 1e-06 
0.666666666667 -1.35353535354 0 0.8 1e-06 
0.722222222222 -1.35353535354 0 0.8 1e-06 
0.777777777778 -1.35353535354 0 0.8 1e-06 
0.833333333333 -1.35353535354 0 0.8 1e-06 
0.888888888889 -1.35353535354 0 0.8 1e-06 
0.944444444444 -1.35353535354 0 0.8 1e-06 
1.0 -1.35353535354 0 0.8 1e-06 
0.5 -1.31313131313 0 0.8 1e-06 
0.555555555556 -1.31313131313 0 0.8 1e-06 
0.611111111111 -1.31313131313 0 0.8 1e-06 
0.666666666667 -1.31313131313 0 0.8 1e-06 
0.722222222222 -1.31313131313 0 0.8 1e-06 
0.777777777778 -1.31313131313 0 0.8 1e-06 
0.833333333333 -1.31313131313 0 0.8 1e-06 
0.888888888889 -1.31313131313 0 0.8 1e-06 
0.944444444444 -1.31313131313 0 0.8 1e-06 
1.0 -1.31313131313 0 0.8 1e-06 
0.5 -1.27272727273 0 0.8 1e-06 
0.555555555556 -1.27272727273 0 0.8 1e-06 
0.611111111111 -1.27272727273 0 0.8 1e-06 
0.666666666667 -1.27272727273 0 0.8 1e-06 
0.722222222222 -1.27272727273 0 0.8 1e-06 
0.777777777778 -1.27272727273 0 0.8 1e-06 
0.833333333333 -1.27272727273 0 0.8 1e-06 
0.888888888889 -1.27272727273 0 0.8 1e-06 
0.944444444444 -1.27272727273 0 0.8 1e-06 
1.0 -1.27272727273 0 0.8 1e-06 
0.5 -1.23232323232 0 0.8 1e-06 
0.555555555556 -1.23232323232 0 0.8 1e-06 
0.611111111111 -1.23232323232 0 0.8 1e-06 
0.666666666667 -1.23232323232 0 0.8 1e-06 
0.722222222222 -1.23232323232 0 0.8 1e-06 
0.777777777778 -1.23232323232 0 0.8 1e-06 
0.833333333333 -1.23232323232 0 0.8 1e-06 
0.888888888889 -1.23232323232 0 0.8 1e-06 
0.944444444444 -1.23232323232 0 0.8 1e-06 
1.0 -1.23232323232 0 0.8 1e-06 
0.5 -1.19191919192 0 0.8 1e-06 
0.555555555556 -1.19191919192 0 0.8 1e-06 
0.611111111111 -1.19191919192 0 0.8 1e-06 
0.666666666667 -1.19191919192 0 0.8 1e-06 
0.722222222222 -1.19191919192 0 0.8 1e-06 
0.777777777778 -1.19191919192 0 0.8 1e-06 
0.833333333333 -1.19191919192 0 0.8 1e-06 
0.888888888889 -1.19191919192 0 0.8 1e-06 
0.944444444444 -1.19191919192 0 0.8 1e-06 
1.0 -1.19191919192 0 0.8 1e-06 
0.5 -1.15151515152 0 0.8 1e-06 
0.555555555556 -1.15151515152 0 0.8 1e-06 
0.611111111111 -1.15151515152 0 0.8 1e-06 
0.666666666667 -1.15151515152 0 0.8 1e-06 
0.722222222222 -1.15151515152 0 0.8 1e-06 
0.777777777778 -1.15151515152 0 0.8 1e-06 
0.833333333333 -1.15151515152 0 0.8 1e-06 
0.888888888889 -1.15151515152 0 0.8 1e-06 
0.944444444444 -1.15151515152 0 0.8 1e-06 
1.0 -1.15151515152 0 0.8 1e-06 
0.5 -1.11111111111 0 0.8 1e-06 
0.555555555556 -1.11111111111 0 0.8 1e-06 
0.611111111111 -1.11111111111 0 0.8 1e-06 
0.666666666667 -1.11111111111 0 0.8 1e-06 
0.722222222222 -1.11111111111 0 0.8 1e-06 
0.777777777778 -1.11111111111 0 0.8 1e-06 
0.833333333333 -1.11111111111 0 0.8 1e-06 
0.888888888889 -1.11111111111 0 0.8 1e-06 
0.944444444444 -1.11111111111 0 0.8 1e-06 
1.0 -1.11111111111 0 0.8 1e-06 
0.5 -1.07070707071 0 0.8 1e-06 
0.555555555556 -1.07070707071 0 0.8 1e-06 
0.611111111111 -1.07070707071 0 0.8 1e-06 
0.666666666667 -1.07070707071 0 0.8 1e-06 
0.722222222222 -1.07070707071 0 0.8 1e-06 
0.777777777778 -1.07070707071 0 0.8 1e-06 
0.833333333333 -1.07070707071 0 0.8 1e-06 
0.888888888889 -1.07070707071 0 0.8 1e-06 
0.944444444444 -1.07070707071 0 0.8 1e-06 
1.0 -1.07070707071 0 0.8 1e-06 
0.5 -1.0303030303 0 0.8 1e-06 
0.555555555556 -1.0303030303 0 0.8 1e-06 
0.611111111111 -1.0303030303 0 0.8 1e-06 
0.666666666667 -1.0303030303 0 0.8 1e-06 
0.722222222222 -1.0303030303 0 0.8 1e-06 
0.777777777778 -1.0303030303 0 0.8 1e-06 
0.833333333333 -1.0303030303 0 0.8 1e-06 
0.888888888889 -1.0303030303 0 0.8 1e-06 
0.944444444444 -1.0303030303 0 0.8 1e-06 
1.0 -1.0303030303 0 0.8 1e-06 
0.5 -0.989898989899 0 0.8 1e-06 
0.555555555556 -0.989898989899 0 0.8 1e-06 
0.611111111111 -0.989898989899 0 0.8 1e-06 
0.666666666667 -0.989898989899 0 0.8 1e-06 
0.722222222222 -0.989898989899 0 0.8 1e-06 
0.777777777778 -0.989898989899 0 0.8 1e-06 
0.833333333333 -0.989898989899 0 0.8 1e-06 
0.888888888889 -0.989898989899 0 0.8 1e-06 
0.944444444444 -0.989898989899 0 0.8 1e-06 
1.0 -0.989898989899 0 0.8 1e-06 
0.5 -0.949494949495 0 0.8 1e-06 
0.555555555556 -0.949494949495 0 0.8 1e-06 
0.611111111111 -0.949494949495 0 0.8 1e-06 
0.666666666667 -0.949494949495 0 0.8 1e-06 
0.722222222222 -0.949494949495 0 0.8 1e-06 
0.777777777778 -0.949494949495 0 0.8 1e-06 
0.833333333333 -0.949494949495 0 0.8 1e-06 
0.888888888889 -0.949494949495 0 0.8 1e-06 
0.944444444444 -0.949494949495 0 0.8 1e-06 
1.0 -0.949494949495 0 0.8 1e-06 
0.5 -0.909090909091 0 0.8 1e-06 
0.555555555556 -0.909090909091 0 0.8 1e-06 
0.611111111111 -0.909090909091 0 0.8 1e-06 
0.666666666667 -0.909090909091 0 0.8 1e-06 
0.722222222222 -0.909090909091 0 0.8 1e-06 
0.777777777778 -0.909090909091 0 0.8 1e-06 
0.833333333333 -0.909090909091 0 0.8 1e-06 
0.888888888889 -0.909090909091 0 0.8 1e-06 
0.944444444444 -0.909090909091 0 0.8 1e-06 
1.0 -0.909090909091 0 0.8 1e-06 
0.5 -0.868686868687 0 0.8 1e-06 
0.555555555556 -0.868686868687 0 0.8 1e-06 
0.611111111111 -0.868686868687 0 0.8 1e-06 
0.666666666667 -0.868686868687 0 0.8 1e-06 
0.722222222222 -0.868686868687 0 0.8 1e-06 
0.777777777778 -0.868686868687 0 0.8 1e-06 
0.833333333333 -0.868686868687 0 0.8 1e-06 
0.888888888889 -0.868686868687 0 0.8 1e-06 
0.944444444444 -0.868686868687 0 0.8 1e-06 
1.0 -0.868686868687 0 0.8 1e-06 
0.5 -0.828282828283 0 0.8 1e-06 
0.555555555556 -0.828282828283 0 0.8 1e-06 
0.611111111111 -0.828282828283 0 0.8 1e-06 
0.666666666667 -0.828282828283 0 0.8 1e-06 
0.722222222222 -0.828282828283 0 0.8 1e-06 
0.777777777778 -0.828282828283 0 0.8 1e-06 
0.833333333333 -0.828282828283 0 0.8 1e-06 
0.888888888889 -0.828282828283 0 0.8 1e-06 
0.944444444444 -0.828282828283 0 0.8 1e-06 
1.0 -0.828282828283 0 0.8 1e-06 
0.5 -0.787878787879 0 0.8 1e-06 
0.555555555556 -0.787878787879 0 0.8 1e-06 
0.611111111111 -0.787878787879 0 0.8 1e-06 
0.666666666667 -0.787878787879 0 0.8 1e-06 
0.722222222222 -0.787878787879 0 0.8 1e-06 
0.777777777778 -0.787878787879 0 0.8 1e-06 
0.833333333333 -0.787878787879 0 0.8 1e-06 
0.888888888889 -0.787878787879 0 0.8 1e-06 
0.944444444444 -0.787878787879 0 0.8 1e-06 
1.0 -0.787878787879 0 0.8 1e-06 
0.5 -0.747474747475 0 0.8 1e-06 
0.555555555556 -0.747474747475 0 0.8 1e-06 
0.611111111111 -0.747474747475 0 0.8 1e-06 
0.666666666667 -0.747474747475 0 0.8 1e-06 
0.722222222222 -0.747474747475 0 0.8 1e-06 
0.777777777778 -0.747474747475 0 0.8 1e-06 
0.833333333333 -0.747474747475 0 0.8 1e-06 
0.888888888889 -0.747474747475 0 0.8 1e-06 
0.944444444444 -0.747474747475 0 0.8 1e-06 
1.0 -0.747474747475 0 0.8 1e-06 
0.5 -0.707070707071 0 0.8 1e-06 
0.555555555556 -0.707070707071 0 0.8 1e-06 
0.611111111111 -0.707070707071 0 0.8 1e-06 
0.666666666667 -0.707070707071 0 0.8 1e-06 
0.722222222222 -0.707070707071 0 0.8 1e-06 
0.777777777778 -0.707070707071 0 0.8 1e-06 
0.833333333333 -0.707070707071 0 0.8 1e-06 
0.888888888889 -0.707070707071 0 0.8 1e-06 
0.944444444444 -0.707070707071 0 0.8 1e-06 
1.0 -0.707070707071 0 0.8 1e-06 
0.5 -0.666666666667 0 0.8 1e-06 
0.555555555556 -0.666666666667 0 0.8 1e-06 
0.611111111111 -0.666666666667 0 0.8 1e-06 
0.666666666667 -0.666666666667 0 0.8 1e-06 
0.722222222222 -0.666666666667 0 0.8 1e-06 
0.777777777778 -0.666666666667 0 0.8 1e-06 
0.833333333333 -0.666666666667 0 0.8 1e-06 
0.888888888889 -0.666666666667 0 0.8 1e-06 
0.944444444444 -0.666666666667 0 0.8 1e-06 
1.0 -0.666666666667 0 0.8 1e-06 
0.5 -0.626262626263 0 0.8 1e-06 
0.555555555556 -0.626262626263 0 0.8 1e-06 
0.611111111111 -0.626262626263 0 0.8 1e-06 
0.666666666667 -0.626262626263 0 0.8 1e-06 
0.722222222222 -0.626262626263 0 0.8 1e-06 
0.777777777778 -0.626262626263 0 0.8 1e-06 
0.833333333333 -0.626262626263 0 0.8 1e-06 
0.888888888889 -0.626262626263 0 0.8 1e-06 
0.944444444444 -0.626262626263 0 0.8 1e-06 
1.0 -0.626262626263 0 0.8 1e-06 
0.5 -0.585858585859 0 0.8 1e-06 
0.555555555556 -0.585858585859 0 0.8 1e-06 
0.611111111111 -0.585858585859 0 0.8 1e-06 
0.666666666667 -0.585858585859 0 0.8 1e-06 
0.722222222222 -0.585858585859 0 0.8 1e-06 
0.777777777778 -0.585858585859 0 0.8 1e-06 
0.833333333333 -0.585858585859 0 0.8 1e-06 
0.888888888889 -0.585858585859 0 0.8 1e-06 
0.944444444444 -0.585858585859 0 0.8 1e-06 
1.0 -0.585858585859 0 0.8 1e-06 
0.5 -0.545454545455 0 0.8 1e-06 
0.555555555556 -0.545454545455 0 0.8 1e-06 
0.611111111111 -0.545454545455 0 0.8 1e-06 
0.666666666667 -0.545454545455 0 0.8 1e-06 
0.722222222222 -0.545454545455 0 0.8 1e-06 
0.777777777778 -0.545454545455 0 0.8 1e-06 
0.833333333333 -0.545454545455 0 0.8 1e-06 
0.888888888889 -0.545454545455 0 0.8 1e-06 
0.944444444444 -0.545454545455 0 0.8 1e-06 
1.0 -0.545454545455 0 0.8 1e-06 
0.5 -0.505050505051 0 0.8 1e-06 
0.555555555556 -0.505050505051 0 0.8 1e-06 
0.611111111111 -0.505050505051 0 0.8 1e-06 
0.666666666667 -0.505050505051 0 0.8 1e-06 
0.722222222222 -0.505050505051 0 0.8 1e-06 
0.777777777778 -0.505050505051 0 0.8 1e-06 
0.833333333333 -0.505050505051 0 0.8 1e-06 
0.888888888889 -0.505050505051 0 0.8 1e-06 
0.944444444444 -0.505050505051 0 0.8 1e-06 
1.0 -0.505050505051 0 0.8 1e-06 
0.5 -0.464646464646 0 0.8 1e-06 
0.555555555556 -0.464646464646 0 0.8 1e-06 
0.611111111111 -0.464646464646 0 0.8 1e-06 
0.666666666667 -0.464646464646 0 0.8 1e-06 
0.722222222222 -0.464646464646 0 0.8 1e-06 
0.777777777778 -0.464646464646 0 0.8 1e-06 
0.833333333333 -0.464646464646 0 0.8 1e-06 
0.888888888889 -0.464646464646 0 0.8 1e-06 
0.944444444444 -0.464646464646 0 0.8 1e-06 
1.0 -0.464646464646 0 0.8 1e-06 
0.5 -0.424242424242 0 0.8 1e-06 
0.555555555556 -0.424242424242 0 0.8 1e-06 
0.611111111111 -0.424242424242 0 0.8 1e-06 
0.666666666667 -0.424242424242 0 0.8 1e-06 
0.722222222222 -0.424242424242 0 0.8 1e-06 
0.777777777778 -0.424242424242 0 0.8 1e-06 
0.833333333333 -0.424242424242 0 0.8 1e-06 
0.888888888889 -0.424242424242 0 0.8 1e-06 
0.944444444444 -0.424242424242 0 0.8 1e-06 
1.0 -0.424242424242 0 0.8 1e-06 
0.5 -0.383838383838 0 0.8 1e-06 
0.555555555556 -0.383838383838 0 0.8 1e-06 
0.611111111111 -0.383838383838 0 0.8 1e-06 
0.666666666667 -0.383838383838 0 0.8 1e-06 
0.722222222222 -0.383838383838 0 0.8 1e-06 
0.777777777778 -0.383838383838 0 0.8 1e-06 
0.833333333333 -0.383838383838 0 0.8 1e-06 
0.888888888889 -0.383838383838 0 0.8 1e-06 
0.944444444444 -0.383838383838 0 0.8 1e-06 
1.0 -0.383838383838 0 0.8 1e-06 
0.5 -0.343434343434 0 0.8 1e-06 
0.555555555556 -0.343434343434 0 0.8 1e-06 
0.611111111111 -0.343434343434 0 0.8 1e-06 
0.666666666667 -0.343434343434 0 0.8 1e-06 
0.722222222222 -0.343434343434 0 0.8 1e-06 
0.777777777778 -0.343434343434 0 0.8 1e-06 
0.833333333333 -0.343434343434 0 0.8 1e-06 
0.888888888889 -0.343434343434 0 0.8 1e-06 
0.944444444444 -0.343434343434 0 0.8 1e-06 
1.0 -0.343434343434 0 0.8 1e-06 
0.5 -0.30303030303 0 0.8 1e-06 
0.555555555556 -0.30303030303 0 0.8 1e-06 
0.611111111111 -0.30303030303 0 0.8 1e-06 
0.666666666667 -0.30303030303 0 0.8 1e-06 
0.722222222222 -0.30303030303 0 0.8 1e-06 
0.777777777778 -0.30303030303 0 0.8 1e-06 
0.833333333333 -0.30303030303 0 0.8 1e-06 
0.888888888889 -0.30303030303 0 0.8 1e-06 
0.944444444444 -0.30303030303 0 0.8 1e-06 
1.0 -0.30303030303 0 0.8 1e-06 
0.5 -0.262626262626 0 0.8 1e-06 
0.555555555556 -0.262626262626 0 0.8 1e-06 
0.611111111111 -0.262626262626 0 0.8 1e-06 
0.666666666667 -0.262626262626 0 0.8 1e-06 
0.722222222222 -0.262626262626 0 0.8 1e-06 
0.777777777778 -0.262626262626 0 0.8 1e-06 
0.833333333333 -0.262626262626 0 0.8 1e-06 
0.888888888889 -0.262626262626 0 0.8 1e-06 
0.944444444444 -0.262626262626 0 0.8 1e-06 
1.0 -0.262626262626 0 0.8 1e-06 
0.5 -0.222222222222 0 0.8 1e-06 
0.555555555556 -0.222222222222 0 0.8 1e-06 
0.611111111111 -0.222222222222 0 0.8 1e-06 
0.666666666667 -0.222222222222 0 0.8 1e-06 
0.722222222222 -0.222222222222 0 0.8 1e-06 
0.777777777778 -0.222222222222 0 0.8 1e-06 
0.833333333333 -0.222222222222 0 0.8 1e-06 
0.888888888889 -0.222222222222 0 0.8 1e-06 
0.944444444444 -0.222222222222 0 0.8 1e-06 
1.0 -0.222222222222 0 0.8 1e-06 
0.5 -0.181818181818 0 0.8 1e-06 
0.555555555556 -0.181818181818 0 0.8 1e-06 
0.611111111111 -0.181818181818 0 0.8 1e-06 
0.666666666667 -0.181818181818 0 0.8 1e-06 
0.722222222222 -0.181818181818 0 0.8 1e-06 
0.777777777778 -0.181818181818 0 0.8 1e-06 
0.833333333333 -0.181818181818 0 0.8 1e-06 
0.888888888889 -0.181818181818 0 0.8 1e-06 
0.944444444444 -0.181818181818 0 0.8 1e-06 
1.0 -0.181818181818 0 0.8 1e-06 
0.5 -0.141414141414 0 0.8 1e-06 
0.555555555556 -0.141414141414 0 0.8 1e-06 
0.611111111111 -0.141414141414 0 0.8 1e-06 
0.666666666667 -0.141414141414 0 0.8 1e-06 
0.722222222222 -0.141414141414 0 0.8 1e-06 
0.777777777778 -0.141414141414 0 0.8 1e-06 
0.833333333333 -0.141414141414 0 0.8 1e-06 
0.888888888889 -0.141414141414 0 0.8 1e-06 
0.944444444444 -0.141414141414 0 0.8 1e-06 
1.0 -0.141414141414 0 0.8 1e-06 
0.5 -0.10101010101 0 0.8 1e-06 
0.555555555556 -0.10101010101 0 0.8 1e-06 
0.611111111111 -0.10101010101 0 0.8 1e-06 
0.666666666667 -0.10101010101 0 0.8 1e-06 
0.722222222222 -0.10101010101 0 0.8 1e-06 
0.777777777778 -0.10101010101 0 0.8 1e-06 
0.833333333333 -0.10101010101 0 0.8 1e-06 
0.888888888889 -0.10101010101 0 0.8 1e-06 
0.944444444444 -0.10101010101 0 0.8 1e-06 
1.0 -0.10101010101 0 0.8 1e-06 
0.5 -0.0606060606061 0 0.8 1e-06 
0.555555555556 -0.0606060606061 0 0.8 1e-06 
0.611111111111 -0.0606060606061 0 0.8 1e-06 
0.666666666667 -0.0606060606061 0 0.8 1e-06 
0.722222222222 -0.0606060606061 0 0.8 1e-06 
0.777777777778 -0.0606060606061 0 0.8 1e-06 
0.833333333333 -0.0606060606061 0 0.8 1e-06 
0.888888888889 -0.0606060606061 0 0.8 1e-06 
0.944444444444 -0.0606060606061 0 0.8 1e-06 
1.0 -0.0606060606061 0 0.8 1e-06 
0.5 -0.020202020202 0 0.8 1e-06 
0.555555555556 -0.020202020202 0 0.8 1e-06 
0.611111111111 -0.020202020202 0 0.8 1e-06 
0.666666666667 -0.020202020202 0 0.8 1e-06 
0.722222222222 -0.020202020202 0 0.8 1e-06 
0.777777777778 -0.020202020202 0 0.8 1e-06 
0.833333333333 -0.020202020202 0 0.8 1e-06 
0.888888888889 -0.020202020202 0 0.8 1e-06 
0.944444444444 -0.020202020202 0 0.8 1e-06 
1.0 -0.020202020202 0 0.8 1e-06 
0.5 0.020202020202 0 0.8 1e-06 
0.555555555556 0.020202020202 0 0.8 1e-06 
0.611111111111 0.020202020202 0 0.8 1e-06 
0.666666666667 0.020202020202 0 0.8 1e-06 
0.722222222222 0.020202020202 0 0.8 1e-06 
0.777777777778 0.020202020202 0 0.8 1e-06 
0.833333333333 0.020202020202 0 0.8 1e-06 
0.888888888889 0.020202020202 0 0.8 1e-06 
0.944444444444 0.020202020202 0 0.8 1e-06 
1.0 0.020202020202 0 0.8 1e-06 
0.5 0.0606060606061 0 0.8 1e-06 
0.555555555556 0.0606060606061 0 0.8 1e-06 
0.611111111111 0.0606060606061 0 0.8 1e-06 
0.666666666667 0.0606060606061 0 0.8 1e-06 
0.722222222222 0.0606060606061 0 0.8 1e-06 
0.777777777778 0.0606060606061 0 0.8 1e-06 
0.833333333333 0.0606060606061 0 0.8 1e-06 
0.888888888889 0.0606060606061 0 0.8 1e-06 
0.944444444444 0.0606060606061 0 0.8 1e-06 
1.0 0.0606060606061 0 0.8 1e-06 
0.5 0.10101010101 0 0.8 1e-06 
0.555555555556 0.10101010101 0 0.8 1e-06 
0.611111111111 0.10101010101 0 0.8 1e-06 
0.666666666667 0.10101010101 0 0.8 1e-06 
0.722222222222 0.10101010101 0 0.8 1e-06 
0.777777777778 0.10101010101 0 0.8 1e-06 
0.833333333333 0.10101010101 0 0.8 1e-06 
0.888888888889 0.10101010101 0 0.8 1e-06 
0.944444444444 0.10101010101 0 0.8 1e-06 
1.0 0.10101010101 0 0.8 1e-06 
0.5 0.141414141414 0 0.8 1e-06 
0.555555555556 0.141414141414 0 0.8 1e-06 
0.611111111111 0.141414141414 0 0.8 1e-06 
0.666666666667 0.141414141414 0 0.8 1e-06 
0.722222222222 0.141414141414 0 0.8 1e-06 
0.777777777778 0.141414141414 0 0.8 1e-06 
0.833333333333 0.141414141414 0 0.8 1e-06 
0.888888888889 0.141414141414 0 0.8 1e-06 
0.944444444444 0.141414141414 0 0.8 1e-06 
1.0 0.141414141414 0 0.8 1e-06 
0.5 0.181818181818 0 0.8 1e-06 
0.555555555556 0.181818181818 0 0.8 1e-06 
0.611111111111 0.181818181818 0 0.8 1e-06 
0.666666666667 0.181818181818 0 0.8 1e-06 
0.722222222222 0.181818181818 0 0.8 1e-06 
0.777777777778 0.181818181818 0 0.8 1e-06 
0.833333333333 0.181818181818 0 0.8 1e-06 
0.888888888889 0.181818181818 0 0.8 1e-06 
0.944444444444 0.181818181818 0 0.8 1e-06 
1.0 0.181818181818 0 0.8 1e-06 
0.5 0.222222222222 0 0.8 1e-06 
0.555555555556 0.222222222222 0 0.8 1e-06 
0.611111111111 0.222222222222 0 0.8 1e-06 
0.666666666667 0.222222222222 0 0.8 1e-06 
0.722222222222 0.222222222222 0 0.8 1e-06 
0.777777777778 0.222222222222 0 0.8 1e-06 
0.833333333333 0.222222222222 0 0.8 1e-06 
0.888888888889 0.222222222222 0 0.8 1e-06 
0.944444444444 0.222222222222 0 0.8 1e-06 
1.0 0.222222222222 0 0.8 1e-06 
0.5 0.262626262626 0 0.8 1e-06 
0.555555555556 0.262626262626 0 0.8 1e-06 
0.611111111111 0.262626262626 0 0.8 1e-06 
0.666666666667 0.262626262626 0 0.8 1e-06 
0.722222222222 0.262626262626 0 0.8 1e-06 
0.777777777778 0.262626262626 0 0.8 1e-06 
0.833333333333 0.262626262626 0 0.8 1e-06 
0.888888888889 0.262626262626 0 0.8 1e-06 
0.944444444444 0.262626262626 0 0.8 1e-06 
1.0 0.262626262626 0 0.8 1e-06 
0.5 0.30303030303 0 0.8 1e-06 
0.555555555556 0.30303030303 0 0.8 1e-06 
0.611111111111 0.30303030303 0 0.8 1e-06 
0.666666666667 0.30303030303 0 0.8 1e-06 
0.722222222222 0.30303030303 0 0.8 1e-06 
0.777777777778 0.30303030303 0 0.8 1e-06 
0.833333333333 0.30303030303 0 0.8 1e-06 
0.888888888889 0.30303030303 0 0.8 1e-06 
0.944444444444 0.30303030303 0 0.8 1e-06 
1.0 0.30303030303 0 0.8 1e-06 
0.5 0.343434343434 0 0.8 1e-06 
0.555555555556 0.343434343434 0 0.8 1e-06 
0.611111111111 0.343434343434 0 0.8 1e-06 
0.666666666667 0.343434343434 0 0.8 1e-06 
0.722222222222 0.343434343434 0 0.8 1e-06 
0.777777777778 0.343434343434 0 0.8 1e-06 
0.833333333333 0.343434343434 0 0.8 1e-06 
0.888888888889 0.343434343434 0 0.8 1e-06 
0.944444444444 0.343434343434 0 0.8 1e-06 
1.0 0.343434343434 0 0.8 1e-06 
0.5 0.383838383838 0 0.8 1e-06 
0.555555555556 0.383838383838 0 0.8 1e-06 
0.611111111111 0.383838383838 0 0.8 1e-06 
0.666666666667 0.383838383838 0 0.8 1e-06 
0.722222222222 0.383838383838 0 0.8 1e-06 
0.777777777778 0.383838383838 0 0.8 1e-06 
0.833333333333 0.383838383838 0 0.8 1e-06 
0.888888888889 0.383838383838 0 0.8 1e-06 
0.944444444444 0.383838383838 0 0.8 1e-06 
1.0 0.383838383838 0 0.8 1e-06 
0.5 0.424242424242 0 0.8 1e-06 
0.555555555556 0.424242424242 0 0.8 1e-06 
0.611111111111 0.424242424242 0 0.8 1e-06 
0.666666666667 0.424242424242 0 0.8 1e-06 
0.722222222222 0.424242424242 0 0.8 1e-06 
0.777777777778 0.424242424242 0 0.8 1e-06 
0.833333333333 0.424242424242 0 0.8 1e-06 
0.888888888889 0.424242424242 0 0.8 1e-06 
0.944444444444 0.424242424242 0 0.8 1e-06 
1.0 0.424242424242 0 0.8 1e-06 
0.5 0.464646464646 0 0.8 1e-06 
0.555555555556 0.464646464646 0 0.8 1e-06 
0.611111111111 0.464646464646 0 0.8 1e-06 
0.666666666667 0.464646464646 0 0.8 1e-06 
0.722222222222 0.464646464646 0 0.8 1e-06 
0.777777777778 0.464646464646 0 0.8 1e-06 
0.833333333333 0.464646464646 0 0.8 1e-06 
0.888888888889 0.464646464646 0 0.8 1e-06 
0.944444444444 0.464646464646 0 0.8 1e-06 
1.0 0.464646464646 0 0.8 1e-06 
0.5 0.505050505051 0 0.8 1e-06 
0.555555555556 0.505050505051 0 0.8 1e-06 
0.611111111111 0.505050505051 0 0.8 1e-06 
0.666666666667 0.505050505051 0 0.8 1e-06 
0.722222222222 0.505050505051 0 0.8 1e-06 
0.777777777778 0.505050505051 0 0.8 1e-06 
0.833333333333 0.505050505051 0 0.8 1e-06 
0.888888888889 0.505050505051 0 0.8 1e-06 
0.944444444444 0.505050505051 0 0.8 1e-06 
1.0 0.505050505051 0 0.8 1e-06 
0.5 0.545454545455 0 0.8 1e-06 
0.555555555556 0.545454545455 0 0.8 1e-06 
0.611111111111 0.545454545455 0 0.8 1e-06 
0.666666666667 0.545454545455 0 0.8 1e-06 
0.722222222222 0.545454545455 0 0.8 1e-06 
0.777777777778 0.545454545455 0 0.8 1e-06 
0.833333333333 0.545454545455 0 0.8 1e-06 
0.888888888889 0.545454545455 0 0.8 1e-06 
0.944444444444 0.545454545455 0 0.8 1e-06 
1.0 0.545454545455 0 0.8 1e-06 
0.5 0.585858585859 0 0.8 1e-06 
0.555555555556 0.585858585859 0 0.8 1e-06 
0.611111111111 0.585858585859 0 0.8 1e-06 
0.666666666667 0.585858585859 0 0.8 1e-06 
0.722222222222 0.585858585859 0 0.8 1e-06 
0.777777777778 0.585858585859 0 0.8 1e-06 
0.833333333333 0.585858585859 0 0.8 1e-06 
0.888888888889 0.585858585859 0 0.8 1e-06 
0.944444444444 0.585858585859 0 0.8 1e-06 
1.0 0.585858585859 0 0.8 1e-06 
0.5 0.626262626263 0 0.8 1e-06 
0.555555555556 0.626262626263 0 0.8 1e-06 
0.611111111111 0.626262626263 0 0.8 1e-06 
0.666666666667 0.626262626263 0 0.8 1e-06 
0.722222222222 0.626262626263 0 0.8 1e-06 
0.777777777778 0.626262626263 0 0.8 1e-06 
0.833333333333 0.626262626263 0 0.8 1e-06 
0.888888888889 0.626262626263 0 0.8 1e-06 
0.944444444444 0.626262626263 0 0.8 1e-06 
1.0 0.626262626263 0 0.8 1e-06 
0.5 0.666666666667 0 0.8 1e-06 
0.555555555556 0.666666666667 0 0.8 1e-06 
0.611111111111 0.666666666667 0 0.8 1e-06 
0.666666666667 0.666666666667 0 0.8 1e-06 
0.722222222222 0.666666666667 0 0.8 1e-06 
0.777777777778 0.666666666667 0 0.8 1e-06 
0.833333333333 0.666666666667 0 0.8 1e-06 
0.888888888889 0.666666666667 0 0.8 1e-06 
0.944444444444 0.666666666667 0 0.8 1e-06 
1.0 0.666666666667 0 0.8 1e-06 
0.5 0.707070707071 0 0.8 1e-06 
0.555555555556 0.707070707071 0 0.8 1e-06 
0.611111111111 0.707070707071 0 0.8 1e-06 
0.666666666667 0.707070707071 0 0.8 1e-06 
0.722222222222 0.707070707071 0 0.8 1e-06 
0.777777777778 0.707070707071 0 0.8 1e-06 
0.833333333333 0.707070707071 0 0.8 1e-06 
0.888888888889 0.707070707071 0 0.8 1e-06 
0.944444444444 0.707070707071 0 0.8 1e-06 
1.0 0.707070707071 0 0.8 1e-06 
0.5 0.747474747475 0 0.8 1e-06 
0.555555555556 0.747474747475 0 0.8 1e-06 
0.611111111111 0.747474747475 0 0.8 1e-06 
0.666666666667 0.747474747475 0 0.8 1e-06 
0.722222222222 0.747474747475 0 0.8 1e-06 
0.777777777778 0.747474747475 0 0.8 1e-06 
0.833333333333 0.747474747475 0 0.8 1e-06 
0.888888888889 0.747474747475 0 0.8 1e-06 
0.944444444444 0.747474747475 0 0.8 1e-06 
1.0 0.747474747475 0 0.8 1e-06 
0.5 0.787878787879 0 0.8 1e-06 
0.555555555556 0.787878787879 0 0.8 1e-06 
0.611111111111 0.787878787879 0 0.8 1e-06 
0.666666666667 0.787878787879 0 0.8 1e-06 
0.722222222222 0.787878787879 0 0.8 1e-06 
0.777777777778 0.787878787879 0 0.8 1e-06 
0.833333333333 0.787878787879 0 0.8 1e-06 
0.888888888889 0.787878787879 0 0.8 1e-06 
0.944444444444 0.787878787879 0 0.8 1e-06 
1.0 0.787878787879 0 0.8 1e-06 
0.5 0.828282828283 0 0.8 1e-06 
0.555555555556 0.828282828283 0 0.8 1e-06 
0.611111111111 0.828282828283 0 0.8 1e-06 
0.666666666667 0.828282828283 0 0.8 1e-06 
0.722222222222 0.828282828283 0 0.8 1e-06 
0.777777777778 0.828282828283 0 0.8 1e-06 
0.833333333333 0.828282828283 0 0.8 1e-06 
0.888888888889 0.828282828283 0 0.8 1e-06 
0.944444444444 0.828282828283 0 0.8 1e-06 
1.0 0.828282828283 0 0.8 1e-06 
0.5 0.868686868687 0 0.8 1e-06 
0.555555555556 0.868686868687 0 0.8 1e-06 
0.611111111111 0.868686868687 0 0.8 1e-06 
0.666666666667 0.868686868687 0 0.8 1e-06 
0.722222222222 0.868686868687 0 0.8 1e-06 
0.777777777778 0.868686868687 0 0.8 1e-06 
0.833333333333 0.868686868687 0 0.8 1e-06 
0.888888888889 0.868686868687 0 0.8 1e-06 
0.944444444444 0.868686868687 0 0.8 1e-06 
1.0 0.868686868687 0 0.8 1e-06 
0.5 0.909090909091 0 0.8 1e-06 
0.555555555556 0.909090909091 0 0.8 1e-06 
0.611111111111 0.909090909091 0 0.8 1e-06 
0.666666666667 0.909090909091 0 0.8 1e-06 
0.722222222222 0.909090909091 0 0.8 1e-06 
0.777777777778 0.909090909091 0 0.8 1e-06 
0.833333333333 0.909090909091 0 0.8 1e-06 
0.888888888889 0.909090909091 0 0.8 1e-06 
0.944444444444 0.909090909091 0 0.8 1e-06 
1.0 0.909090909091 0 0.8 1e-06 
0.5 0.949494949495 0 0.8 1e-06 
0.555555555556 0.949494949495 0 0.8 1e-06 
0.611111111111 0.949494949495 0 0.8 1e-06 
0.666666666667 0.949494949495 0 0.8 1e-06 
0.722222222222 0.949494949495 0 0.8 1e-06 
0.777777777778 0.949494949495 0 0.8 1e-06 
0.833333333333 0.949494949495 0 0.8 1e-06 
0.888888888889 0.949494949495 0 0.8 1e-06 
0.944444444444 0.949494949495 0 0.8 1e-06 
1.0 0.949494949495 0 0.8 1e-06 
0.5 0.989898989899 0 0.8 1e-06 
0.555555555556 0.989898989899 0 0.8 1e-06 
0.611111111111 0.989898989899 0 0.8 1e-06 
0.666666666667 0.989898989899 0 0.8 1e-06 
0.722222222222 0.989898989899 0 0.8 1e-06 
0.777777777778 0.989898989899 0 0.8 1e-06 
0.833333333333 0.989898989899 0 0.8 1e-06 
0.888888888889 0.989898989899 0 0.8 1e-06 
0.944444444444 0.989898989899 0 0.8 1e-06 
1.0 0.989898989899 0 0.8 1e-06 
0.5 1.0303030303 0 0.8 1e-06 
0.555555555556 1.0303030303 0 0.8 1e-06 
0.611111111111 1.0303030303 0 0.8 1e-06 
0.666666666667 1.0303030303 0 0.8 1e-06 
0.722222222222 1.0303030303 0 0.8 1e-06 
0.777777777778 1.0303030303 0 0.8 1e-06 
0.833333333333 1.0303030303 0 0.8 1e-06 
0.888888888889 1.0303030303 0 0.8 1e-06 
0.944444444444 1.0303030303 0 0.8 1e-06 
1.0 1.0303030303 0 0.8 1e-06 
0.5 1.07070707071 0 0.8 1e-06 
0.555555555556 1.07070707071 0 0.8 1e-06 
0.611111111111 1.07070707071 0 0.8 1e-06 
0.666666666667 1.07070707071 0 0.8 1e-06 
0.722222222222 1.07070707071 0 0.8 1e-06 
0.777777777778 1.07070707071 0 0.8 1e-06 
0.833333333333 1.07070707071 0 0.8 1e-06 
0.888888888889 1.07070707071 0 0.8 1e-06 
0.944444444444 1.07070707071 0 0.8 1e-06 
1.0 1.07070707071 0 0.8 1e-06 
0.5 1.11111111111 0 0.8 1e-06 
0.555555555556 1.11111111111 0 0.8 1e-06 
0.611111111111 1.11111111111 0 0.8 1e-06 
0.666666666667 1.11111111111 0 0.8 1e-06 
0.722222222222 1.11111111111 0 0.8 1e-06 
0.777777777778 1.11111111111 0 0.8 1e-06 
0.833333333333 1.11111111111 0 0.8 1e-06 
0.888888888889 1.11111111111 0 0.8 1e-06 
0.944444444444 1.11111111111 0 0.8 1e-06 
1.0 1.11111111111 0 0.8 1e-06 
0.5 1.15151515152 0 0.8 1e-06 
0.555555555556 1.15151515152 0 0.8 1e-06 
0.611111111111 1.15151515152 0 0.8 1e-06 
0.666666666667 1.15151515152 0 0.8 1e-06 
0.722222222222 1.15151515152 0 0.8 1e-06 
0.777777777778 1.15151515152 0 0.8 1e-06 
0.833333333333 1.15151515152 0 0.8 1e-06 
0.888888888889 1.15151515152 0 0.8 1e-06 
0.944444444444 1.15151515152 0 0.8 1e-06 
1.0 1.15151515152 0 0.8 1e-06 
0.5 1.19191919192 0 0.8 1e-06 
0.555555555556 1.19191919192 0 0.8 1e-06 
0.611111111111 1.19191919192 0 0.8 1e-06 
0.666666666667 1.19191919192 0 0.8 1e-06 
0.722222222222 1.19191919192 0 0.8 1e-06 
0.777777777778 1.19191919192 0 0.8 1e-06 
0.833333333333 1.19191919192 0 0.8 1e-06 
0.888888888889 1.19191919192 0 0.8 1e-06 
0.944444444444 1.19191919192 0 0.8 1e-06 
1.0 1.19191919192 0 0.8 1e-06 
0.5 1.23232323232 0 0.8 1e-06 
0.555555555556 1.23232323232 0 0.8 1e-06 
0.611111111111 1.23232323232 0 0.8 1e-06 
0.666666666667 1.23232323232 0 0.8 1e-06 
0.722222222222 1.23232323232 0 0.8 1e-06 
0.777777777778 1.23232323232 0 0.8 1e-06 
0.833333333333 1.23232323232 0 0.8 1e-06 
0.888888888889 1.23232323232 0 0.8 1e-06 
0.944444444444 1.23232323232 0 0.8 1e-06 
1.0 1.23232323232 0 0.8 1e-06 
0.5 1.27272727273 0 0.8 1e-06 
0.555555555556 1.27272727273 0 0.8 1e-06 
0.611111111111 1.27272727273 0 0.8 1e-06 
0.666666666667 1.27272727273 0 0.8 1e-06 
0.722222222222 1.27272727273 0 0.8 1e-06 
0.777777777778 1.27272727273 0 0.8 1e-06 
0.833333333333 1.27272727273 0 0.8 1e-06 
0.888888888889 1.27272727273 0 0.8 1e-06 
0.944444444444 1.27272727273 0 0.8 1e-06 
1.0 1.27272727273 0 0.8 1e-06 
0.5 1.31313131313 0 0.8 1e-06 
0.555555555556 1.31313131313 0 0.8 1e-06 
0.611111111111 1.31313131313 0 0.8 1e-06 
0.666666666667 1.31313131313 0 0.8 1e-06 
0.722222222222 1.31313131313 0 0.8 1e-06 
0.777777777778 1.31313131313 0 0.8 1e-06 
0.833333333333 1.31313131313 0 0.8 1e-06 
0.888888888889 1.31313131313 0 0.8 1e-06 
0.944444444444 1.31313131313 0 0.8 1e-06 
1.0 1.31313131313 0 0.8 1e-06 
0.5 1.35353535354 0 0.8 1e-06 
0.555555555556 1.35353535354 0 0.8 1e-06 
0.611111111111 1.35353535354 0 0.8 1e-06 
0.666666666667 1.35353535354 0 0.8 1e-06 
0.722222222222 1.35353535354 0 0.8 1e-06 
0.777777777778 1.35353535354 0 0.8 1e-06 
0.833333333333 1.35353535354 0 0.8 1e-06 
0.888888888889 1.35353535354 0 0.8 1e-06 
0.944444444444 1.35353535354 0 0.8 1e-06 
1.0 1.35353535354 0 0.8 1e-06 
0.5 1.39393939394 0 0.8 1e-06 
0.555555555556 1.39393939394 0 0.8 1e-06 
0.611111111111 1.39393939394 0 0.8 1e-06 
0.666666666667 1.39393939394 0 0.8 1e-06 
0.722222222222 1.39393939394 0 0.8 1e-06 
0.777777777778 1.39393939394 0 0.8 1e-06 
0.833333333333 1.39393939394 0 0.8 1e-06 
0.888888888889 1.39393939394 0 0.8 1e-06 
0.944444444444 1.39393939394 0 0.8 1e-06 
1.0 1.39393939394 0 0.8 1e-06 
0.5 1.43434343434 0 0.8 1e-06 
0.555555555556 1.43434343434 0 0.8 1e-06 
0.611111111111 1.43434343434 0 0.8 1e-06 
0.666666666667 1.43434343434 0 0.8 1e-06 
0.722222222222 1.43434343434 0 0.8 1e-06 
0.777777777778 1.43434343434 0 0.8 1e-06 
0.833333333333 1.43434343434 0 0.8 1e-06 
0.888888888889 1.43434343434 0 0.8 1e-06 
0.944444444444 1.43434343434 0 0.8 1e-06 
1.0 1.43434343434 0 0.8 1e-06 
0.5 1.47474747475 0 0.8 1e-06 
0.555555555556 1.47474747475 0 0.8 1e-06 
0.611111111111 1.47474747475 0 0.8 1e-06 
0.666666666667 1.47474747475 0 0.8 1e-06 
0.722222222222 1.47474747475 0 0.8 1e-06 
0.777777777778 1.47474747475 0 0.8 1e-06 
0.833333333333 1.47474747475 0 0.8 1e-06 
0.888888888889 1.47474747475 0 0.8 1e-06 
0.944444444444 1.47474747475 0 0.8 1e-06 
1.0 1.47474747475 0 0.8 1e-06 
0.5 1.51515151515 0 0.8 1e-06 
0.555555555556 1.51515151515 0 0.8 1e-06 
0.611111111111 1.51515151515 0 0.8 1e-06 
0.666666666667 1.51515151515 0 0.8 1e-06 
0.722222222222 1.51515151515 0 0.8 1e-06 
0.777777777778 1.51515151515 0 0.8 1e-06 
0.833333333333 1.51515151515 0 0.8 1e-06 
0.888888888889 1.51515151515 0 0.8 1e-06 
0.944444444444 1.51515151515 0 0.8 1e-06 
1.0 1.51515151515 0 0.8 1e-06 
0.5 1.55555555556 0 0.8 1e-06 
0.555555555556 1.55555555556 0 0.8 1e-06 
0.611111111111 1.55555555556 0 0.8 1e-06 
0.666666666667 1.55555555556 0 0.8 1e-06 
0.722222222222 1.55555555556 0 0.8 1e-06 
0.777777777778 1.55555555556 0 0.8 1e-06 
0.833333333333 1.55555555556 0 0.8 1e-06 
0.888888888889 1.55555555556 0 0.8 1e-06 
0.944444444444 1.55555555556 0 0.8 1e-06 
1.0 1.55555555556 0 0.8 1e-06 
0.5 1.59595959596 0 0.8 1e-06 
0.555555555556 1.59595959596 0 0.8 1e-06 
0.611111111111 1.59595959596 0 0.8 1e-06 
0.666666666667 1.59595959596 0 0.8 1e-06 
0.722222222222 1.59595959596 0 0.8 1e-06 
0.777777777778 1.59595959596 0 0.8 1e-06 
0.833333333333 1.59595959596 0 0.8 1e-06 
0.888888888889 1.59595959596 0 0.8 1e-06 
0.944444444444 1.59595959596 0 0.8 1e-06 
1.0 1.59595959596 0 0.8 1e-06 
0.5 1.63636363636 0 0.8 1e-06 
0.555555555556 1.63636363636 0 0.8 1e-06 
0.611111111111 1.63636363636 0 0.8 1e-06 
0.666666666667 1.63636363636 0 0.8 1e-06 
0.722222222222 1.63636363636 0 0.8 1e-06 
0.777777777778 1.63636363636 0 0.8 1e-06 
0.833333333333 1.63636363636 0 0.8 1e-06 
0.888888888889 1.63636363636 0 0.8 1e-06 
0.944444444444 1.63636363636 0 0.8 1e-06 
1.0 1.63636363636 0 0.8 1e-06 
0.5 1.67676767677 0 0.8 1e-06 
0.555555555556 1.67676767677 0 0.8 1e-06 
0.611111111111 1.67676767677 0 0.8 1e-06 
0.666666666667 1.67676767677 0 0.8 1e-06 
0.722222222222 1.67676767677 0 0.8 1e-06 
0.777777777778 1.67676767677 0 0.8 1e-06 
0.833333333333 1.67676767677 0 0.8 1e-06 
0.888888888889 1.67676767677 0 0.8 1e-06 
0.944444444444 1.67676767677 0 0.8 1e-06 
1.0 1.67676767677 0 0.8 1e-06 
0.5 1.71717171717 0 0.8 1e-06 
0.555555555556 1.71717171717 0 0.8 1e-06 
0.611111111111 1.71717171717 0 0.8 1e-06 
0.666666666667 1.71717171717 0 0.8 1e-06 
0.722222222222 1.71717171717 0 0.8 1e-06 
0.777777777778 1.71717171717 0 0.8 1e-06 
0.833333333333 1.71717171717 0 0.8 1e-06 
0.888888888889 1.71717171717 0 0.8 1e-06 
0.944444444444 1.71717171717 0 0.8 1e-06 
1.0 1.71717171717 0 0.8 1e-06 
0.5 1.75757575758 0 0.8 1e-06 
0.555555555556 1.75757575758 0 0.8 1e-06 
0.611111111111 1.75757575758 0 0.8 1e-06 
0.666666666667 1.75757575758 0 0.8 1e-06 
0.722222222222 1.75757575758 0 0.8 1e-06 
0.777777777778 1.75757575758 0 0.8 1e-06 
0.833333333333 1.75757575758 0 0.8 1e-06 
0.888888888889 1.75757575758 0 0.8 1e-06 
0.944444444444 1.75757575758 0 0.8 1e-06 
1.0 1.75757575758 0 0.8 1e-06 
0.5 1.79797979798 0 0.8 1e-06 
0.555555555556 1.79797979798 0 0.8 1e-06 
0.611111111111 1.79797979798 0 0.8 1e-06 
0.666666666667 1.79797979798 0 0.8 1e-06 
0.722222222222 1.79797979798 0 0.8 1e-06 
0.777777777778 1.79797979798 0 0.8 1e-06 
0.833333333333 1.79797979798 0 0.8 1e-06 
0.888888888889 1.79797979798 0 0.8 1e-06 
0.944444444444 1.79797979798 0 0.8 1e-06 
1.0 1.79797979798 0 0.8 1e-06 
0.5 1.83838383838 0 0.8 1e-06 
0.555555555556 1.83838383838 0 0.8 1e-06 
0.611111111111 1.83838383838 0 0.8 1e-06 
0.666666666667 1.83838383838 0 0.8 1e-06 
0.722222222222 1.83838383838 0 0.8 1e-06 
0.777777777778 1.83838383838 0 0.8 1e-06 
0.833333333333 1.83838383838 0 0.8 1e-06 
0.888888888889 1.83838383838 0 0.8 1e-06 
0.944444444444 1.83838383838 0 0.8 1e-06 
1.0 1.83838383838 0 0.8 1e-06 
0.5 1.87878787879 0 0.8 1e-06 
0.555555555556 1.87878787879 0 0.8 1e-06 
0.611111111111 1.87878787879 0 0.8 1e-06 
0.666666666667 1.87878787879 0 0.8 1e-06 
0.722222222222 1.87878787879 0 0.8 1e-06 
0.777777777778 1.87878787879 0 0.8 1e-06 
0.833333333333 1.87878787879 0 0.8 1e-06 
0.888888888889 1.87878787879 0 0.8 1e-06 
0.944444444444 1.87878787879 0 0.8 1e-06 
1.0 1.87878787879 0 0.8 1e-06 
0.5 1.91919191919 0 0.8 1e-06 
0.555555555556 1.91919191919 0 0.8 1e-06 
0.611111111111 1.91919191919 0 0.8 1e-06 
0.666666666667 1.91919191919 0 0.8 1e-06 
0.722222222222 1.91919191919 0 0.8 1e-06 
0.777777777778 1.91919191919 0 0.8 1e-06 
0.833333333333 1.91919191919 0 0.8 1e-06 
0.888888888889 1.91919191919 0 0.8 1e-06 
0.944444444444 1.91919191919 0 0.8 1e-06 
1.0 1.91919191919 0 0.8 1e-06 
0.5 1.9595959596 0 0.8 1e-06 
0.555555555556 1.9595959596 0 0.8 1e-06 
0.611111111111 1.9595959596 0 0.8 1e-06 
0.666666666667 1.9595959596 0 0.8 1e-06 
0.722222222222 1.9595959596 0 0.8 1e-06 
0.777777777778 1.9595959596 0 0.8 1e-06 
0.833333333333 1.9595959596 0 0.8 1e-06 
0.888888888889 1.9595959596 0 0.8 1e-06 
0.944444444444 1.9595959596 0 0.8 1e-06 
1.0 1.9595959596 0 0.8 1e-06 
0.5 2.0 0 0.8 1e-06 
0.555555555556 2.0 0 0.8 1e-06 
0.611111111111 2.0 0 0.8 1e-06 
0.666666666667 2.0 0 0.8 1e-06 
0.722222222222 2.0 0 0.8 1e-06 
0.777777777778 2.0 0 0.8 1e-06 
0.833333333333 2.0 0 0.8 1e-06 
0.888888888889 2.0 0 0.8 1e-06 
0.944444444444 2.0 0 0.8 1e-06 
1.0 2.0 0 0.8 1e-06 
0.5 -2.0 0 1.2 1e-06 
0.555555555556 -2.0 0 1.2 1e-06 
0.611111111111 -2.0 0 1.2 1e-06 
0.666666666667 -2.0 0 1.2 1e-06 
0.722222222222 -2.0 0 1.2 1e-06 
0.777777777778 -2.0 0 1.2 1e-06 
0.833333333333 -2.0 0 1.2 1e-06 
0.888888888889 -2.0 0 1.2 1e-06 
0.944444444444 -2.0 0 1.2 1e-06 
1.0 -2.0 0 1.2 1e-06 
0.5 -1.9595959596 0 1.2 1e-06 
0.555555555556 -1.9595959596 0 1.2 1e-06 
0.611111111111 -1.9595959596 0 1.2 1e-06 
0.666666666667 -1.9595959596 0 1.2 1e-06 
0.722222222222 -1.9595959596 0 1.2 1e-06 
0.777777777778 -1.9595959596 0 1.2 1e-06 
0.833333333333 -1.9595959596 0 1.2 1e-06 
0.888888888889 -1.9595959596 0 1.2 1e-06 
0.944444444444 -1.9595959596 0 1.2 1e-06 
1.0 -1.9595959596 0 1.2 1e-06 
0.5 -1.91919191919 0 1.2 1e-06 
0.555555555556 -1.91919191919 0 1.2 1e-06 
0.611111111111 -1.91919191919 0 1.2 1e-06 
0.666666666667 -1.91919191919 0 1.2 1e-06 
0.722222222222 -1.91919191919 0 1.2 1e-06 
0.777777777778 -1.91919191919 0 1.2 1e-06 
0.833333333333 -1.91919191919 0 1.2 1e-06 
0.888888888889 -1.91919191919 0 1.2 1e-06 
0.944444444444 -1.91919191919 0 1.2 1e-06 
1.0 -1.91919191919 0 1.2 1e-06 
0.5 -1.87878787879 0 1.2 1e-06 
0.555555555556 -1.87878787879 0 1.2 1e-06 
0.611111111111 -1.87878787879 0 1.2 1e-06 
0.666666666667 -1.87878787879 0 1.2 1e-06 
0.722222222222 -1.87878787879 0 1.2 1e-06 
0.777777777778 -1.87878787879 0 1.2 1e-06 
0.833333333333 -1.87878787879 0 1.2 1e-06 
0.888888888889 -1.87878787879 0 1.2 1e-06 
0.944444444444 -1.87878787879 0 1.2 1e-06 
1.0 -1.87878787879 0 1.2 1e-06 
0.5 -1.83838383838 0 1.2 1e-06 
0.555555555556 -1.83838383838 0 1.2 1e-06 
0.611111111111 -1.83838383838 0 1.2 1e-06 
0.666666666667 -1.83838383838 0 1.2 1e-06 
0.722222222222 -1.83838383838 0 1.2 1e-06 
0.777777777778 -1.83838383838 0 1.2 1e-06 
0.833333333333 -1.83838383838 0 1.2 1e-06 
0.888888888889 -1.83838383838 0 1.2 1e-06 
0.944444444444 -1.83838383838 0 1.2 1e-06 
1.0 -1.83838383838 0 1.2 1e-06 
0.5 -1.79797979798 0 1.2 1e-06 
0.555555555556 -1.79797979798 0 1.2 1e-06 
0.611111111111 -1.79797979798 0 1.2 1e-06 
0.666666666667 -1.79797979798 0 1.2 1e-06 
0.722222222222 -1.79797979798 0 1.2 1e-06 
0.777777777778 -1.79797979798 0 1.2 1e-06 
0.833333333333 -1.79797979798 0 1.2 1e-06 
0.888888888889 -1.79797979798 0 1.2 1e-06 
0.944444444444 -1.79797979798 0 1.2 1e-06 
1.0 -1.79797979798 0 1.2 1e-06 
0.5 -1.75757575758 0 1.2 1e-06 
0.555555555556 -1.75757575758 0 1.2 1e-06 
0.611111111111 -1.75757575758 0 1.2 1e-06 
0.666666666667 -1.75757575758 0 1.2 1e-06 
0.722222222222 -1.75757575758 0 1.2 1e-06 
0.777777777778 -1.75757575758 0 1.2 1e-06 
0.833333333333 -1.75757575758 0 1.2 1e-06 
0.888888888889 -1.75757575758 0 1.2 1e-06 
0.944444444444 -1.75757575758 0 1.2 1e-06 
1.0 -1.75757575758 0 1.2 1e-06 
0.5 -1.71717171717 0 1.2 1e-06 
0.555555555556 -1.71717171717 0 1.2 1e-06 
0.611111111111 -1.71717171717 0 1.2 1e-06 
0.666666666667 -1.71717171717 0 1.2 1e-06 
0.722222222222 -1.71717171717 0 1.2 1e-06 
0.777777777778 -1.71717171717 0 1.2 1e-06 
0.833333333333 -1.71717171717 0 1.2 1e-06 
0.888888888889 -1.71717171717 0 1.2 1e-06 
0.944444444444 -1.71717171717 0 1.2 1e-06 
1.0 -1.71717171717 0 1.2 1e-06 
0.5 -1.67676767677 0 1.2 1e-06 
0.555555555556 -1.67676767677 0 1.2 1e-06 
0.611111111111 -1.67676767677 0 1.2 1e-06 
0.666666666667 -1.67676767677 0 1.2 1e-06 
0.722222222222 -1.67676767677 0 1.2 1e-06 
0.777777777778 -1.67676767677 0 1.2 1e-06 
0.833333333333 -1.67676767677 0 1.2 1e-06 
0.888888888889 -1.67676767677 0 1.2 1e-06 
0.944444444444 -1.67676767677 0 1.2 1e-06 
1.0 -1.67676767677 0 1.2 1e-06 
0.5 -1.63636363636 0 1.2 1e-06 
0.555555555556 -1.63636363636 0 1.2 1e-06 
0.611111111111 -1.63636363636 0 1.2 1e-06 
0.666666666667 -1.63636363636 0 1.2 1e-06 
0.722222222222 -1.63636363636 0 1.2 1e-06 
0.777777777778 -1.63636363636 0 1.2 1e-06 
0.833333333333 -1.63636363636 0 1.2 1e-06 
0.888888888889 -1.63636363636 0 1.2 1e-06 
0.944444444444 -1.63636363636 0 1.2 1e-06 
1.0 -1.63636363636 0 1.2 1e-06 
0.5 -1.59595959596 0 1.2 1e-06 
0.555555555556 -1.59595959596 0 1.2 1e-06 
0.611111111111 -1.59595959596 0 1.2 1e-06 
0.666666666667 -1.59595959596 0 1.2 1e-06 
0.722222222222 -1.59595959596 0 1.2 1e-06 
0.777777777778 -1.59595959596 0 1.2 1e-06 
0.833333333333 -1.59595959596 0 1.2 1e-06 
0.888888888889 -1.59595959596 0 1.2 1e-06 
0.944444444444 -1.59595959596 0 1.2 1e-06 
1.0 -1.59595959596 0 1.2 1e-06 
0.5 -1.55555555556 0 1.2 1e-06 
0.555555555556 -1.55555555556 0 1.2 1e-06 
0.611111111111 -1.55555555556 0 1.2 1e-06 
0.666666666667 -1.55555555556 0 1.2 1e-06 
0.722222222222 -1.55555555556 0 1.2 1e-06 
0.777777777778 -1.55555555556 0 1.2 1e-06 
0.833333333333 -1.55555555556 0 1.2 1e-06 
0.888888888889 -1.55555555556 0 1.2 1e-06 
0.944444444444 -1.55555555556 0 1.2 1e-06 
1.0 -1.55555555556 0 1.2 1e-06 
0.5 -1.51515151515 0 1.2 1e-06 
0.555555555556 -1.51515151515 0 1.2 1e-06 
0.611111111111 -1.51515151515 0 1.2 1e-06 
0.666666666667 -1.51515151515 0 1.2 1e-06 
0.722222222222 -1.51515151515 0 1.2 1e-06 
0.777777777778 -1.51515151515 0 1.2 1e-06 
0.833333333333 -1.51515151515 0 1.2 1e-06 
0.888888888889 -1.51515151515 0 1.2 1e-06 
0.944444444444 -1.51515151515 0 1.2 1e-06 
1.0 -1.51515151515 0 1.2 1e-06 
0.5 -1.47474747475 0 1.2 1e-06 
0.555555555556 -1.47474747475 0 1.2 1e-06 
0.611111111111 -1.47474747475 0 1.2 1e-06 
0.666666666667 -1.47474747475 0 1.2 1e-06 
0.722222222222 -1.47474747475 0 1.2 1e-06 
0.777777777778 -1.47474747475 0 1.2 1e-06 
0.833333333333 -1.47474747475 0 1.2 1e-06 
0.888888888889 -1.47474747475 0 1.2 1e-06 
0.944444444444 -1.47474747475 0 1.2 1e-06 
1.0 -1.47474747475 0 1.2 1e-06 
0.5 -1.43434343434 0 1.2 1e-06 
0.555555555556 -1.43434343434 0 1.2 1e-06 
0.611111111111 -1.43434343434 0 1.2 1e-06 
0.666666666667 -1.43434343434 0 1.2 1e-06 
0.722222222222 -1.43434343434 0 1.2 1e-06 
0.777777777778 -1.43434343434 0 1.2 1e-06 
0.833333333333 -1.43434343434 0 1.2 1e-06 
0.888888888889 -1.43434343434 0 1.2 1e-06 
0.944444444444 -1.43434343434 0 1.2 1e-06 
1.0 -1.43434343434 0 1.2 1e-06 
0.5 -1.39393939394 0 1.2 1e-06 
0.555555555556 -1.39393939394 0 1.2 1e-06 
0.611111111111 -1.39393939394 0 1.2 1e-06 
0.666666666667 -1.39393939394 0 1.2 1e-06 
0.722222222222 -1.39393939394 0 1.2 1e-06 
0.777777777778 -1.39393939394 0 1.2 1e-06 
0.833333333333 -1.39393939394 0 1.2 1e-06 
0.888888888889 -1.39393939394 0 1.2 1e-06 
0.944444444444 -1.39393939394 0 1.2 1e-06 
1.0 -1.39393939394 0 1.2 1e-06 
0.5 -1.35353535354 0 1.2 1e-06 
0.555555555556 -1.35353535354 0 1.2 1e-06 
0.611111111111 -1.35353535354 0 1.2 1e-06 
0.666666666667 -1.35353535354 0 1.2 1e-06 
0.722222222222 -1.35353535354 0 1.2 1e-06 
0.777777777778 -1.35353535354 0 1.2 1e-06 
0.833333333333 -1.35353535354 0 1.2 1e-06 
0.888888888889 -1.35353535354 0 1.2 1e-06 
0.944444444444 -1.35353535354 0 1.2 1e-06 
1.0 -1.35353535354 0 1.2 1e-06 
0.5 -1.31313131313 0 1.2 1e-06 
0.555555555556 -1.31313131313 0 1.2 1e-06 
0.611111111111 -1.31313131313 0 1.2 1e-06 
0.666666666667 -1.31313131313 0 1.2 1e-06 
0.722222222222 -1.31313131313 0 1.2 1e-06 
0.777777777778 -1.31313131313 0 1.2 1e-06 
0.833333333333 -1.31313131313 0 1.2 1e-06 
0.888888888889 -1.31313131313 0 1.2 1e-06 
0.944444444444 -1.31313131313 0 1.2 1e-06 
1.0 -1.31313131313 0 1.2 1e-06 
0.5 -1.27272727273 0 1.2 1e-06 
0.555555555556 -1.27272727273 0 1.2 1e-06 
0.611111111111 -1.27272727273 0 1.2 1e-06 
0.666666666667 -1.27272727273 0 1.2 1e-06 
0.722222222222 -1.27272727273 0 1.2 1e-06 
0.777777777778 -1.27272727273 0 1.2 1e-06 
0.833333333333 -1.27272727273 0 1.2 1e-06 
0.888888888889 -1.27272727273 0 1.2 1e-06 
0.944444444444 -1.27272727273 0 1.2 1e-06 
1.0 -1.27272727273 0 1.2 1e-06 
0.5 -1.23232323232 0 1.2 1e-06 
0.555555555556 -1.23232323232 0 1.2 1e-06 
0.611111111111 -1.23232323232 0 1.2 1e-06 
0.666666666667 -1.23232323232 0 1.2 1e-06 
0.722222222222 -1.23232323232 0 1.2 1e-06 
0.777777777778 -1.23232323232 0 1.2 1e-06 
0.833333333333 -1.23232323232 0 1.2 1e-06 
0.888888888889 -1.23232323232 0 1.2 1e-06 
0.944444444444 -1.23232323232 0 1.2 1e-06 
1.0 -1.23232323232 0 1.2 1e-06 
0.5 -1.19191919192 0 1.2 1e-06 
0.555555555556 -1.19191919192 0 1.2 1e-06 
0.611111111111 -1.19191919192 0 1.2 1e-06 
0.666666666667 -1.19191919192 0 1.2 1e-06 
0.722222222222 -1.19191919192 0 1.2 1e-06 
0.777777777778 -1.19191919192 0 1.2 1e-06 
0.833333333333 -1.19191919192 0 1.2 1e-06 
0.888888888889 -1.19191919192 0 1.2 1e-06 
0.944444444444 -1.19191919192 0 1.2 1e-06 
1.0 -1.19191919192 0 1.2 1e-06 
0.5 -1.15151515152 0 1.2 1e-06 
0.555555555556 -1.15151515152 0 1.2 1e-06 
0.611111111111 -1.15151515152 0 1.2 1e-06 
0.666666666667 -1.15151515152 0 1.2 1e-06 
0.722222222222 -1.15151515152 0 1.2 1e-06 
0.777777777778 -1.15151515152 0 1.2 1e-06 
0.833333333333 -1.15151515152 0 1.2 1e-06 
0.888888888889 -1.15151515152 0 1.2 1e-06 
0.944444444444 -1.15151515152 0 1.2 1e-06 
1.0 -1.15151515152 0 1.2 1e-06 
0.5 -1.11111111111 0 1.2 1e-06 
0.555555555556 -1.11111111111 0 1.2 1e-06 
0.611111111111 -1.11111111111 0 1.2 1e-06 
0.666666666667 -1.11111111111 0 1.2 1e-06 
0.722222222222 -1.11111111111 0 1.2 1e-06 
0.777777777778 -1.11111111111 0 1.2 1e-06 
0.833333333333 -1.11111111111 0 1.2 1e-06 
0.888888888889 -1.11111111111 0 1.2 1e-06 
0.944444444444 -1.11111111111 0 1.2 1e-06 
1.0 -1.11111111111 0 1.2 1e-06 
0.5 -1.07070707071 0 1.2 1e-06 
0.555555555556 -1.07070707071 0 1.2 1e-06 
0.611111111111 -1.07070707071 0 1.2 1e-06 
0.666666666667 -1.07070707071 0 1.2 1e-06 
0.722222222222 -1.07070707071 0 1.2 1e-06 
0.777777777778 -1.07070707071 0 1.2 1e-06 
0.833333333333 -1.07070707071 0 1.2 1e-06 
0.888888888889 -1.07070707071 0 1.2 1e-06 
0.944444444444 -1.07070707071 0 1.2 1e-06 
1.0 -1.07070707071 0 1.2 1e-06 
0.5 -1.0303030303 0 1.2 1e-06 
0.555555555556 -1.0303030303 0 1.2 1e-06 
0.611111111111 -1.0303030303 0 1.2 1e-06 
0.666666666667 -1.0303030303 0 1.2 1e-06 
0.722222222222 -1.0303030303 0 1.2 1e-06 
0.777777777778 -1.0303030303 0 1.2 1e-06 
0.833333333333 -1.0303030303 0 1.2 1e-06 
0.888888888889 -1.0303030303 0 1.2 1e-06 
0.944444444444 -1.0303030303 0 1.2 1e-06 
1.0 -1.0303030303 0 1.2 1e-06 
0.5 -0.989898989899 0 1.2 1e-06 
0.555555555556 -0.989898989899 0 1.2 1e-06 
0.611111111111 -0.989898989899 0 1.2 1e-06 
0.666666666667 -0.989898989899 0 1.2 1e-06 
0.722222222222 -0.989898989899 0 1.2 1e-06 
0.777777777778 -0.989898989899 0 1.2 1e-06 
0.833333333333 -0.989898989899 0 1.2 1e-06 
0.888888888889 -0.989898989899 0 1.2 1e-06 
0.944444444444 -0.989898989899 0 1.2 1e-06 
1.0 -0.989898989899 0 1.2 1e-06 
0.5 -0.949494949495 0 1.2 1e-06 
0.555555555556 -0.949494949495 0 1.2 1e-06 
0.611111111111 -0.949494949495 0 1.2 1e-06 
0.666666666667 -0.949494949495 0 1.2 1e-06 
0.722222222222 -0.949494949495 0 1.2 1e-06 
0.777777777778 -0.949494949495 0 1.2 1e-06 
0.833333333333 -0.949494949495 0 1.2 1e-06 
0.888888888889 -0.949494949495 0 1.2 1e-06 
0.944444444444 -0.949494949495 0 1.2 1e-06 
1.0 -0.949494949495 0 1.2 1e-06 
0.5 -0.909090909091 0 1.2 1e-06 
0.555555555556 -0.909090909091 0 1.2 1e-06 
0.611111111111 -0.909090909091 0 1.2 1e-06 
0.666666666667 -0.909090909091 0 1.2 1e-06 
0.722222222222 -0.909090909091 0 1.2 1e-06 
0.777777777778 -0.909090909091 0 1.2 1e-06 
0.833333333333 -0.909090909091 0 1.2 1e-06 
0.888888888889 -0.909090909091 0 1.2 1e-06 
0.944444444444 -0.909090909091 0 1.2 1e-06 
1.0 -0.909090909091 0 1.2 1e-06 
0.5 -0.868686868687 0 1.2 1e-06 
0.555555555556 -0.868686868687 0 1.2 1e-06 
0.611111111111 -0.868686868687 0 1.2 1e-06 
0.666666666667 -0.868686868687 0 1.2 1e-06 
0.722222222222 -0.868686868687 0 1.2 1e-06 
0.777777777778 -0.868686868687 0 1.2 1e-06 
0.833333333333 -0.868686868687 0 1.2 1e-06 
0.888888888889 -0.868686868687 0 1.2 1e-06 
0.944444444444 -0.868686868687 0 1.2 1e-06 
1.0 -0.868686868687 0 1.2 1e-06 
0.5 -0.828282828283 0 1.2 1e-06 
0.555555555556 -0.828282828283 0 1.2 1e-06 
0.611111111111 -0.828282828283 0 1.2 1e-06 
0.666666666667 -0.828282828283 0 1.2 1e-06 
0.722222222222 -0.828282828283 0 1.2 1e-06 
0.777777777778 -0.828282828283 0 1.2 1e-06 
0.833333333333 -0.828282828283 0 1.2 1e-06 
0.888888888889 -0.828282828283 0 1.2 1e-06 
0.944444444444 -0.828282828283 0 1.2 1e-06 
1.0 -0.828282828283 0 1.2 1e-06 
0.5 -0.787878787879 0 1.2 1e-06 
0.555555555556 -0.787878787879 0 1.2 1e-06 
0.611111111111 -0.787878787879 0 1.2 1e-06 
0.666666666667 -0.787878787879 0 1.2 1e-06 
0.722222222222 -0.787878787879 0 1.2 1e-06 
0.777777777778 -0.787878787879 0 1.2 1e-06 
0.833333333333 -0.787878787879 0 1.2 1e-06 
0.888888888889 -0.787878787879 0 1.2 1e-06 
0.944444444444 -0.787878787879 0 1.2 1e-06 
1.0 -0.787878787879 0 1.2 1e-06 
0.5 -0.747474747475 0 1.2 1e-06 
0.555555555556 -0.747474747475 0 1.2 1e-06 
0.611111111111 -0.747474747475 0 1.2 1e-06 
0.666666666667 -0.747474747475 0 1.2 1e-06 
0.722222222222 -0.747474747475 0 1.2 1e-06 
0.777777777778 -0.747474747475 0 1.2 1e-06 
0.833333333333 -0.747474747475 0 1.2 1e-06 
0.888888888889 -0.747474747475 0 1.2 1e-06 
0.944444444444 -0.747474747475 0 1.2 1e-06 
1.0 -0.747474747475 0 1.2 1e-06 
0.5 -0.707070707071 0 1.2 1e-06 
0.555555555556 -0.707070707071 0 1.2 1e-06 
0.611111111111 -0.707070707071 0 1.2 1e-06 
0.666666666667 -0.707070707071 0 1.2 1e-06 
0.722222222222 -0.707070707071 0 1.2 1e-06 
0.777777777778 -0.707070707071 0 1.2 1e-06 
0.833333333333 -0.707070707071 0 1.2 1e-06 
0.888888888889 -0.707070707071 0 1.2 1e-06 
0.944444444444 -0.707070707071 0 1.2 1e-06 
1.0 -0.707070707071 0 1.2 1e-06 
0.5 -0.666666666667 0 1.2 1e-06 
0.555555555556 -0.666666666667 0 1.2 1e-06 
0.611111111111 -0.666666666667 0 1.2 1e-06 
0.666666666667 -0.666666666667 0 1.2 1e-06 
0.722222222222 -0.666666666667 0 1.2 1e-06 
0.777777777778 -0.666666666667 0 1.2 1e-06 
0.833333333333 -0.666666666667 0 1.2 1e-06 
0.888888888889 -0.666666666667 0 1.2 1e-06 
0.944444444444 -0.666666666667 0 1.2 1e-06 
1.0 -0.666666666667 0 1.2 1e-06 
0.5 -0.626262626263 0 1.2 1e-06 
0.555555555556 -0.626262626263 0 1.2 1e-06 
0.611111111111 -0.626262626263 0 1.2 1e-06 
0.666666666667 -0.626262626263 0 1.2 1e-06 
0.722222222222 -0.626262626263 0 1.2 1e-06 
0.777777777778 -0.626262626263 0 1.2 1e-06 
0.833333333333 -0.626262626263 0 1.2 1e-06 
0.888888888889 -0.626262626263 0 1.2 1e-06 
0.944444444444 -0.626262626263 0 1.2 1e-06 
1.0 -0.626262626263 0 1.2 1e-06 
0.5 -0.585858585859 0 1.2 1e-06 
0.555555555556 -0.585858585859 0 1.2 1e-06 
0.611111111111 -0.585858585859 0 1.2 1e-06 
0.666666666667 -0.585858585859 0 1.2 1e-06 
0.722222222222 -0.585858585859 0 1.2 1e-06 
0.777777777778 -0.585858585859 0 1.2 1e-06 
0.833333333333 -0.585858585859 0 1.2 1e-06 
0.888888888889 -0.585858585859 0 1.2 1e-06 
0.944444444444 -0.585858585859 0 1.2 1e-06 
1.0 -0.585858585859 0 1.2 1e-06 
0.5 -0.545454545455 0 1.2 1e-06 
0.555555555556 -0.545454545455 0 1.2 1e-06 
0.611111111111 -0.545454545455 0 1.2 1e-06 
0.666666666667 -0.545454545455 0 1.2 1e-06 
0.722222222222 -0.545454545455 0 1.2 1e-06 
0.777777777778 -0.545454545455 0 1.2 1e-06 
0.833333333333 -0.545454545455 0 1.2 1e-06 
0.888888888889 -0.545454545455 0 1.2 1e-06 
0.944444444444 -0.545454545455 0 1.2 1e-06 
1.0 -0.545454545455 0 1.2 1e-06 
0.5 -0.505050505051 0 1.2 1e-06 
0.555555555556 -0.505050505051 0 1.2 1e-06 
0.611111111111 -0.505050505051 0 1.2 1e-06 
0.666666666667 -0.505050505051 0 1.2 1e-06 
0.722222222222 -0.505050505051 0 1.2 1e-06 
0.777777777778 -0.505050505051 0 1.2 1e-06 
0.833333333333 -0.505050505051 0 1.2 1e-06 
0.888888888889 -0.505050505051 0 1.2 1e-06 
0.944444444444 -0.505050505051 0 1.2 1e-06 
1.0 -0.505050505051 0 1.2 1e-06 
0.5 -0.464646464646 0 1.2 1e-06 
0.555555555556 -0.464646464646 0 1.2 1e-06 
0.611111111111 -0.464646464646 0 1.2 1e-06 
0.666666666667 -0.464646464646 0 1.2 1e-06 
0.722222222222 -0.464646464646 0 1.2 1e-06 
0.777777777778 -0.464646464646 0 1.2 1e-06 
0.833333333333 -0.464646464646 0 1.2 1e-06 
0.888888888889 -0.464646464646 0 1.2 1e-06 
0.944444444444 -0.464646464646 0 1.2 1e-06 
1.0 -0.464646464646 0 1.2 1e-06 
0.5 -0.424242424242 0 1.2 1e-06 
0.555555555556 -0.424242424242 0 1.2 1e-06 
0.611111111111 -0.424242424242 0 1.2 1e-06 
0.666666666667 -0.424242424242 0 1.2 1e-06 
0.722222222222 -0.424242424242 0 1.2 1e-06 
0.777777777778 -0.424242424242 0 1.2 1e-06 
0.833333333333 -0.424242424242 0 1.2 1e-06 
0.888888888889 -0.424242424242 0 1.2 1e-06 
0.944444444444 -0.424242424242 0 1.2 1e-06 
1.0 -0.424242424242 0 1.2 1e-06 
0.5 -0.383838383838 0 1.2 1e-06 
0.555555555556 -0.383838383838 0 1.2 1e-06 
0.611111111111 -0.383838383838 0 1.2 1e-06 
0.666666666667 -0.383838383838 0 1.2 1e-06 
0.722222222222 -0.383838383838 0 1.2 1e-06 
0.777777777778 -0.383838383838 0 1.2 1e-06 
0.833333333333 -0.383838383838 0 1.2 1e-06 
0.888888888889 -0.383838383838 0 1.2 1e-06 
0.944444444444 -0.383838383838 0 1.2 1e-06 
1.0 -0.383838383838 0 1.2 1e-06 
0.5 -0.343434343434 0 1.2 1e-06 
0.555555555556 -0.343434343434 0 1.2 1e-06 
0.611111111111 -0.343434343434 0 1.2 1e-06 
0.666666666667 -0.343434343434 0 1.2 1e-06 
0.722222222222 -0.343434343434 0 1.2 1e-06 
0.777777777778 -0.343434343434 0 1.2 1e-06 
0.833333333333 -0.343434343434 0 1.2 1e-06 
0.888888888889 -0.343434343434 0 1.2 1e-06 
0.944444444444 -0.343434343434 0 1.2 1e-06 
1.0 -0.343434343434 0 1.2 1e-06 
0.5 -0.30303030303 0 1.2 1e-06 
0.555555555556 -0.30303030303 0 1.2 1e-06 
0.611111111111 -0.30303030303 0 1.2 1e-06 
0.666666666667 -0.30303030303 0 1.2 1e-06 
0.722222222222 -0.30303030303 0 1.2 1e-06 
0.777777777778 -0.30303030303 0 1.2 1e-06 
0.833333333333 -0.30303030303 0 1.2 1e-06 
0.888888888889 -0.30303030303 0 1.2 1e-06 
0.944444444444 -0.30303030303 0 1.2 1e-06 
1.0 -0.30303030303 0 1.2 1e-06 
0.5 -0.262626262626 0 1.2 1e-06 
0.555555555556 -0.262626262626 0 1.2 1e-06 
0.611111111111 -0.262626262626 0 1.2 1e-06 
0.666666666667 -0.262626262626 0 1.2 1e-06 
0.722222222222 -0.262626262626 0 1.2 1e-06 
0.777777777778 -0.262626262626 0 1.2 1e-06 
0.833333333333 -0.262626262626 0 1.2 1e-06 
0.888888888889 -0.262626262626 0 1.2 1e-06 
0.944444444444 -0.262626262626 0 1.2 1e-06 
1.0 -0.262626262626 0 1.2 1e-06 
0.5 -0.222222222222 0 1.2 1e-06 
0.555555555556 -0.222222222222 0 1.2 1e-06 
0.611111111111 -0.222222222222 0 1.2 1e-06 
0.666666666667 -0.222222222222 0 1.2 1e-06 
0.722222222222 -0.222222222222 0 1.2 1e-06 
0.777777777778 -0.222222222222 0 1.2 1e-06 
0.833333333333 -0.222222222222 0 1.2 1e-06 
0.888888888889 -0.222222222222 0 1.2 1e-06 
0.944444444444 -0.222222222222 0 1.2 1e-06 
1.0 -0.222222222222 0 1.2 1e-06 
0.5 -0.181818181818 0 1.2 1e-06 
0.555555555556 -0.181818181818 0 1.2 1e-06 
0.611111111111 -0.181818181818 0 1.2 1e-06 
0.666666666667 -0.181818181818 0 1.2 1e-06 
0.722222222222 -0.181818181818 0 1.2 1e-06 
0.777777777778 -0.181818181818 0 1.2 1e-06 
0.833333333333 -0.181818181818 0 1.2 1e-06 
0.888888888889 -0.181818181818 0 1.2 1e-06 
0.944444444444 -0.181818181818 0 1.2 1e-06 
1.0 -0.181818181818 0 1.2 1e-06 
0.5 -0.141414141414 0 1.2 1e-06 
0.555555555556 -0.141414141414 0 1.2 1e-06 
0.611111111111 -0.141414141414 0 1.2 1e-06 
0.666666666667 -0.141414141414 0 1.2 1e-06 
0.722222222222 -0.141414141414 0 1.2 1e-06 
0.777777777778 -0.141414141414 0 1.2 1e-06 
0.833333333333 -0.141414141414 0 1.2 1e-06 
0.888888888889 -0.141414141414 0 1.2 1e-06 
0.944444444444 -0.141414141414 0 1.2 1e-06 
1.0 -0.141414141414 0 1.2 1e-06 
0.5 -0.10101010101 0 1.2 1e-06 
0.555555555556 -0.10101010101 0 1.2 1e-06 
0.611111111111 -0.10101010101 0 1.2 1e-06 
0.666666666667 -0.10101010101 0 1.2 1e-06 
0.722222222222 -0.10101010101 0 1.2 1e-06 
0.777777777778 -0.10101010101 0 1.2 1e-06 
0.833333333333 -0.10101010101 0 1.2 1e-06 
0.888888888889 -0.10101010101 0 1.2 1e-06 
0.944444444444 -0.10101010101 0 1.2 1e-06 
1.0 -0.10101010101 0 1.2 1e-06 
0.5 -0.0606060606061 0 1.2 1e-06 
0.555555555556 -0.0606060606061 0 1.2 1e-06 
0.611111111111 -0.0606060606061 0 1.2 1e-06 
0.666666666667 -0.0606060606061 0 1.2 1e-06 
0.722222222222 -0.0606060606061 0 1.2 1e-06 
0.777777777778 -0.0606060606061 0 1.2 1e-06 
0.833333333333 -0.0606060606061 0 1.2 1e-06 
0.888888888889 -0.0606060606061 0 1.2 1e-06 
0.944444444444 -0.0606060606061 0 1.2 1e-06 
1.0 -0.0606060606061 0 1.2 1e-06 
0.5 -0.020202020202 0 1.2 1e-06 
0.555555555556 -0.020202020202 0 1.2 1e-06 
0.611111111111 -0.020202020202 0 1.2 1e-06 
0.666666666667 -0.020202020202 0 1.2 1e-06 
0.722222222222 -0.020202020202 0 1.2 1e-06 
0.777777777778 -0.020202020202 0 1.2 1e-06 
0.833333333333 -0.020202020202 0 1.2 1e-06 
0.888888888889 -0.020202020202 0 1.2 1e-06 
0.944444444444 -0.020202020202 0 1.2 1e-06 
1.0 -0.020202020202 0 1.2 1e-06 
0.5 0.020202020202 0 1.2 1e-06 
0.555555555556 0.020202020202 0 1.2 1e-06 
0.611111111111 0.020202020202 0 1.2 1e-06 
0.666666666667 0.020202020202 0 1.2 1e-06 
0.722222222222 0.020202020202 0 1.2 1e-06 
0.777777777778 0.020202020202 0 1.2 1e-06 
0.833333333333 0.020202020202 0 1.2 1e-06 
0.888888888889 0.020202020202 0 1.2 1e-06 
0.944444444444 0.020202020202 0 1.2 1e-06 
1.0 0.020202020202 0 1.2 1e-06 
0.5 0.0606060606061 0 1.2 1e-06 
0.555555555556 0.0606060606061 0 1.2 1e-06 
0.611111111111 0.0606060606061 0 1.2 1e-06 
0.666666666667 0.0606060606061 0 1.2 1e-06 
0.722222222222 0.0606060606061 0 1.2 1e-06 
0.777777777778 0.0606060606061 0 1.2 1e-06 
0.833333333333 0.0606060606061 0 1.2 1e-06 
0.888888888889 0.0606060606061 0 1.2 1e-06 
0.944444444444 0.0606060606061 0 1.2 1e-06 
1.0 0.0606060606061 0 1.2 1e-06 
0.5 0.10101010101 0 1.2 1e-06 
0.555555555556 0.10101010101 0 1.2 1e-06 
0.611111111111 0.10101010101 0 1.2 1e-06 
0.666666666667 0.10101010101 0 1.2 1e-06 
0.722222222222 0.10101010101 0 1.2 1e-06 
0.777777777778 0.10101010101 0 1.2 1e-06 
0.833333333333 0.10101010101 0 1.2 1e-06 
0.888888888889 0.10101010101 0 1.2 1e-06 
0.944444444444 0.10101010101 0 1.2 1e-06 
1.0 0.10101010101 0 1.2 1e-06 
0.5 0.141414141414 0 1.2 1e-06 
0.555555555556 0.141414141414 0 1.2 1e-06 
0.611111111111 0.141414141414 0 1.2 1e-06 
0.666666666667 0.141414141414 0 1.2 1e-06 
0.722222222222 0.141414141414 0 1.2 1e-06 
0.777777777778 0.141414141414 0 1.2 1e-06 
0.833333333333 0.141414141414 0 1.2 1e-06 
0.888888888889 0.141414141414 0 1.2 1e-06 
0.944444444444 0.141414141414 0 1.2 1e-06 
1.0 0.141414141414 0 1.2 1e-06 
0.5 0.181818181818 0 1.2 1e-06 
0.555555555556 0.181818181818 0 1.2 1e-06 
0.611111111111 0.181818181818 0 1.2 1e-06 
0.666666666667 0.181818181818 0 1.2 1e-06 
0.722222222222 0.181818181818 0 1.2 1e-06 
0.777777777778 0.181818181818 0 1.2 1e-06 
0.833333333333 0.181818181818 0 1.2 1e-06 
0.888888888889 0.181818181818 0 1.2 1e-06 
0.944444444444 0.181818181818 0 1.2 1e-06 
1.0 0.181818181818 0 1.2 1e-06 
0.5 0.222222222222 0 1.2 1e-06 
0.555555555556 0.222222222222 0 1.2 1e-06 
0.611111111111 0.222222222222 0 1.2 1e-06 
0.666666666667 0.222222222222 0 1.2 1e-06 
0.722222222222 0.222222222222 0 1.2 1e-06 
0.777777777778 0.222222222222 0 1.2 1e-06 
0.833333333333 0.222222222222 0 1.2 1e-06 
0.888888888889 0.222222222222 0 1.2 1e-06 
0.944444444444 0.222222222222 0 1.2 1e-06 
1.0 0.222222222222 0 1.2 1e-06 
0.5 0.262626262626 0 1.2 1e-06 
0.555555555556 0.262626262626 0 1.2 1e-06 
0.611111111111 0.262626262626 0 1.2 1e-06 
0.666666666667 0.262626262626 0 1.2 1e-06 
0.722222222222 0.262626262626 0 1.2 1e-06 
0.777777777778 0.262626262626 0 1.2 1e-06 
0.833333333333 0.262626262626 0 1.2 1e-06 
0.888888888889 0.262626262626 0 1.2 1e-06 
0.944444444444 0.262626262626 0 1.2 1e-06 
1.0 0.262626262626 0 1.2 1e-06 
0.5 0.30303030303 0 1.2 1e-06 
0.555555555556 0.30303030303 0 1.2 1e-06 
0.611111111111 0.30303030303 0 1.2 1e-06 
0.666666666667 0.30303030303 0 1.2 1e-06 
0.722222222222 0.30303030303 0 1.2 1e-06 
0.777777777778 0.30303030303 0 1.2 1e-06 
0.833333333333 0.30303030303 0 1.2 1e-06 
0.888888888889 0.30303030303 0 1.2 1e-06 
0.944444444444 0.30303030303 0 1.2 1e-06 
1.0 0.30303030303 0 1.2 1e-06 
0.5 0.343434343434 0 1.2 1e-06 
0.555555555556 0.343434343434 0 1.2 1e-06 
0.611111111111 0.343434343434 0 1.2 1e-06 
0.666666666667 0.343434343434 0 1.2 1e-06 
0.722222222222 0.343434343434 0 1.2 1e-06 
0.777777777778 0.343434343434 0 1.2 1e-06 
0.833333333333 0.343434343434 0 1.2 1e-06 
0.888888888889 0.343434343434 0 1.2 1e-06 
0.944444444444 0.343434343434 0 1.2 1e-06 
1.0 0.343434343434 0 1.2 1e-06 
0.5 0.383838383838 0 1.2 1e-06 
0.555555555556 0.383838383838 0 1.2 1e-06 
0.611111111111 0.383838383838 0 1.2 1e-06 
0.666666666667 0.383838383838 0 1.2 1e-06 
0.722222222222 0.383838383838 0 1.2 1e-06 
0.777777777778 0.383838383838 0 1.2 1e-06 
0.833333333333 0.383838383838 0 1.2 1e-06 
0.888888888889 0.383838383838 0 1.2 1e-06 
0.944444444444 0.383838383838 0 1.2 1e-06 
1.0 0.383838383838 0 1.2 1e-06 
0.5 0.424242424242 0 1.2 1e-06 
0.555555555556 0.424242424242 0 1.2 1e-06 
0.611111111111 0.424242424242 0 1.2 1e-06 
0.666666666667 0.424242424242 0 1.2 1e-06 
0.722222222222 0.424242424242 0 1.2 1e-06 
0.777777777778 0.424242424242 0 1.2 1e-06 
0.833333333333 0.424242424242 0 1.2 1e-06 
0.888888888889 0.424242424242 0 1.2 1e-06 
0.944444444444 0.424242424242 0 1.2 1e-06 
1.0 0.424242424242 0 1.2 1e-06 
0.5 0.464646464646 0 1.2 1e-06 
0.555555555556 0.464646464646 0 1.2 1e-06 
0.611111111111 0.464646464646 0 1.2 1e-06 
0.666666666667 0.464646464646 0 1.2 1e-06 
0.722222222222 0.464646464646 0 1.2 1e-06 
0.777777777778 0.464646464646 0 1.2 1e-06 
0.833333333333 0.464646464646 0 1.2 1e-06 
0.888888888889 0.464646464646 0 1.2 1e-06 
0.944444444444 0.464646464646 0 1.2 1e-06 
1.0 0.464646464646 0 1.2 1e-06 
0.5 0.505050505051 0 1.2 1e-06 
0.555555555556 0.505050505051 0 1.2 1e-06 
0.611111111111 0.505050505051 0 1.2 1e-06 
0.666666666667 0.505050505051 0 1.2 1e-06 
0.722222222222 0.505050505051 0 1.2 1e-06 
0.777777777778 0.505050505051 0 1.2 1e-06 
0.833333333333 0.505050505051 0 1.2 1e-06 
0.888888888889 0.505050505051 0 1.2 1e-06 
0.944444444444 0.505050505051 0 1.2 1e-06 
1.0 0.505050505051 0 1.2 1e-06 
0.5 0.545454545455 0 1.2 1e-06 
0.555555555556 0.545454545455 0 1.2 1e-06 
0.611111111111 0.545454545455 0 1.2 1e-06 
0.666666666667 0.545454545455 0 1.2 1e-06 
0.722222222222 0.545454545455 0 1.2 1e-06 
0.777777777778 0.545454545455 0 1.2 1e-06 
0.833333333333 0.545454545455 0 1.2 1e-06 
0.888888888889 0.545454545455 0 1.2 1e-06 
0.944444444444 0.545454545455 0 1.2 1e-06 
1.0 0.545454545455 0 1.2 1e-06 
0.5 0.585858585859 0 1.2 1e-06 
0.555555555556 0.585858585859 0 1.2 1e-06 
0.611111111111 0.585858585859 0 1.2 1e-06 
0.666666666667 0.585858585859 0 1.2 1e-06 
0.722222222222 0.585858585859 0 1.2 1e-06 
0.777777777778 0.585858585859 0 1.2 1e-06 
0.833333333333 0.585858585859 0 1.2 1e-06 
0.888888888889 0.585858585859 0 1.2 1e-06 
0.944444444444 0.585858585859 0 1.2 1e-06 
1.0 0.585858585859 0 1.2 1e-06 
0.5 0.626262626263 0 1.2 1e-06 
0.555555555556 0.626262626263 0 1.2 1e-06 
0.611111111111 0.626262626263 0 1.2 1e-06 
0.666666666667 0.626262626263 0 1.2 1e-06 
0.722222222222 0.626262626263 0 1.2 1e-06 
0.777777777778 0.626262626263 0 1.2 1e-06 
0.833333333333 0.626262626263 0 1.2 1e-06 
0.888888888889 0.626262626263 0 1.2 1e-06 
0.944444444444 0.626262626263 0 1.2 1e-06 
1.0 0.626262626263 0 1.2 1e-06 
0.5 0.666666666667 0 1.2 1e-06 
0.555555555556 0.666666666667 0 1.2 1e-06 
0.611111111111 0.666666666667 0 1.2 1e-06 
0.666666666667 0.666666666667 0 1.2 1e-06 
0.722222222222 0.666666666667 0 1.2 1e-06 
0.777777777778 0.666666666667 0 1.2 1e-06 
0.833333333333 0.666666666667 0 1.2 1e-06 
0.888888888889 0.666666666667 0 1.2 1e-06 
0.944444444444 0.666666666667 0 1.2 1e-06 
1.0 0.666666666667 0 1.2 1e-06 
0.5 0.707070707071 0 1.2 1e-06 
0.555555555556 0.707070707071 0 1.2 1e-06 
0.611111111111 0.707070707071 0 1.2 1e-06 
0.666666666667 0.707070707071 0 1.2 1e-06 
0.722222222222 0.707070707071 0 1.2 1e-06 
0.777777777778 0.707070707071 0 1.2 1e-06 
0.833333333333 0.707070707071 0 1.2 1e-06 
0.888888888889 0.707070707071 0 1.2 1e-06 
0.944444444444 0.707070707071 0 1.2 1e-06 
1.0 0.707070707071 0 1.2 1e-06 
0.5 0.747474747475 0 1.2 1e-06 
0.555555555556 0.747474747475 0 1.2 1e-06 
0.611111111111 0.747474747475 0 1.2 1e-06 
0.666666666667 0.747474747475 0 1.2 1e-06 
0.722222222222 0.747474747475 0 1.2 1e-06 
0.777777777778 0.747474747475 0 1.2 1e-06 
0.833333333333 0.747474747475 0 1.2 1e-06 
0.888888888889 0.747474747475 0 1.2 1e-06 
0.944444444444 0.747474747475 0 1.2 1e-06 
1.0 0.747474747475 0 1.2 1e-06 
0.5 0.787878787879 0 1.2 1e-06 
0.555555555556 0.787878787879 0 1.2 1e-06 
0.611111111111 0.787878787879 0 1.2 1e-06 
0.666666666667 0.787878787879 0 1.2 1e-06 
0.722222222222 0.787878787879 0 1.2 1e-06 
0.777777777778 0.787878787879 0 1.2 1e-06 
0.833333333333 0.787878787879 0 1.2 1e-06 
0.888888888889 0.787878787879 0 1.2 1e-06 
0.944444444444 0.787878787879 0 1.2 1e-06 
1.0 0.787878787879 0 1.2 1e-06 
0.5 0.828282828283 0 1.2 1e-06 
0.555555555556 0.828282828283 0 1.2 1e-06 
0.611111111111 0.828282828283 0 1.2 1e-06 
0.666666666667 0.828282828283 0 1.2 1e-06 
0.722222222222 0.828282828283 0 1.2 1e-06 
0.777777777778 0.828282828283 0 1.2 1e-06 
0.833333333333 0.828282828283 0 1.2 1e-06 
0.888888888889 0.828282828283 0 1.2 1e-06 
0.944444444444 0.828282828283 0 1.2 1e-06 
1.0 0.828282828283 0 1.2 1e-06 
0.5 0.868686868687 0 1.2 1e-06 
0.555555555556 0.868686868687 0 1.2 1e-06 
0.611111111111 0.868686868687 0 1.2 1e-06 
0.666666666667 0.868686868687 0 1.2 1e-06 
0.722222222222 0.868686868687 0 1.2 1e-06 
0.777777777778 0.868686868687 0 1.2 1e-06 
0.833333333333 0.868686868687 0 1.2 1e-06 
0.888888888889 0.868686868687 0 1.2 1e-06 
0.944444444444 0.868686868687 0 1.2 1e-06 
1.0 0.868686868687 0 1.2 1e-06 
0.5 0.909090909091 0 1.2 1e-06 
0.555555555556 0.909090909091 0 1.2 1e-06 
0.611111111111 0.909090909091 0 1.2 1e-06 
0.666666666667 0.909090909091 0 1.2 1e-06 
0.722222222222 0.909090909091 0 1.2 1e-06 
0.777777777778 0.909090909091 0 1.2 1e-06 
0.833333333333 0.909090909091 0 1.2 1e-06 
0.888888888889 0.909090909091 0 1.2 1e-06 
0.944444444444 0.909090909091 0 1.2 1e-06 
1.0 0.909090909091 0 1.2 1e-06 
0.5 0.949494949495 0 1.2 1e-06 
0.555555555556 0.949494949495 0 1.2 1e-06 
0.611111111111 0.949494949495 0 1.2 1e-06 
0.666666666667 0.949494949495 0 1.2 1e-06 
0.722222222222 0.949494949495 0 1.2 1e-06 
0.777777777778 0.949494949495 0 1.2 1e-06 
0.833333333333 0.949494949495 0 1.2 1e-06 
0.888888888889 0.949494949495 0 1.2 1e-06 
0.944444444444 0.949494949495 0 1.2 1e-06 
1.0 0.949494949495 0 1.2 1e-06 
0.5 0.989898989899 0 1.2 1e-06 
0.555555555556 0.989898989899 0 1.2 1e-06 
0.611111111111 0.989898989899 0 1.2 1e-06 
0.666666666667 0.989898989899 0 1.2 1e-06 
0.722222222222 0.989898989899 0 1.2 1e-06 
0.777777777778 0.989898989899 0 1.2 1e-06 
0.833333333333 0.989898989899 0 1.2 1e-06 
0.888888888889 0.989898989899 0 1.2 1e-06 
0.944444444444 0.989898989899 0 1.2 1e-06 
1.0 0.989898989899 0 1.2 1e-06 
0.5 1.0303030303 0 1.2 1e-06 
0.555555555556 1.0303030303 0 1.2 1e-06 
0.611111111111 1.0303030303 0 1.2 1e-06 
0.666666666667 1.0303030303 0 1.2 1e-06 
0.722222222222 1.0303030303 0 1.2 1e-06 
0.777777777778 1.0303030303 0 1.2 1e-06 
0.833333333333 1.0303030303 0 1.2 1e-06 
0.888888888889 1.0303030303 0 1.2 1e-06 
0.944444444444 1.0303030303 0 1.2 1e-06 
1.0 1.0303030303 0 1.2 1e-06 
0.5 1.07070707071 0 1.2 1e-06 
0.555555555556 1.07070707071 0 1.2 1e-06 
0.611111111111 1.07070707071 0 1.2 1e-06 
0.666666666667 1.07070707071 0 1.2 1e-06 
0.722222222222 1.07070707071 0 1.2 1e-06 
0.777777777778 1.07070707071 0 1.2 1e-06 
0.833333333333 1.07070707071 0 1.2 1e-06 
0.888888888889 1.07070707071 0 1.2 1e-06 
0.944444444444 1.07070707071 0 1.2 1e-06 
1.0 1.07070707071 0 1.2 1e-06 
0.5 1.11111111111 0 1.2 1e-06 
0.555555555556 1.11111111111 0 1.2 1e-06 
0.611111111111 1.11111111111 0 1.2 1e-06 
0.666666666667 1.11111111111 0 1.2 1e-06 
0.722222222222 1.11111111111 0 1.2 1e-06 
0.777777777778 1.11111111111 0 1.2 1e-06 
0.833333333333 1.11111111111 0 1.2 1e-06 
0.888888888889 1.11111111111 0 1.2 1e-06 
0.944444444444 1.11111111111 0 1.2 1e-06 
1.0 1.11111111111 0 1.2 1e-06 
0.5 1.15151515152 0 1.2 1e-06 
0.555555555556 1.15151515152 0 1.2 1e-06 
0.611111111111 1.15151515152 0 1.2 1e-06 
0.666666666667 1.15151515152 0 1.2 1e-06 
0.722222222222 1.15151515152 0 1.2 1e-06 
0.777777777778 1.15151515152 0 1.2 1e-06 
0.833333333333 1.15151515152 0 1.2 1e-06 
0.888888888889 1.15151515152 0 1.2 1e-06 
0.944444444444 1.15151515152 0 1.2 1e-06 
1.0 1.15151515152 0 1.2 1e-06 
0.5 1.19191919192 0 1.2 1e-06 
0.555555555556 1.19191919192 0 1.2 1e-06 
0.611111111111 1.19191919192 0 1.2 1e-06 
0.666666666667 1.19191919192 0 1.2 1e-06 
0.722222222222 1.19191919192 0 1.2 1e-06 
0.777777777778 1.19191919192 0 1.2 1e-06 
0.833333333333 1.19191919192 0 1.2 1e-06 
0.888888888889 1.19191919192 0 1.2 1e-06 
0.944444444444 1.19191919192 0 1.2 1e-06 
1.0 1.19191919192 0 1.2 1e-06 
0.5 1.23232323232 0 1.2 1e-06 
0.555555555556 1.23232323232 0 1.2 1e-06 
0.611111111111 1.23232323232 0 1.2 1e-06 
0.666666666667 1.23232323232 0 1.2 1e-06 
0.722222222222 1.23232323232 0 1.2 1e-06 
0.777777777778 1.23232323232 0 1.2 1e-06 
0.833333333333 1.23232323232 0 1.2 1e-06 
0.888888888889 1.23232323232 0 1.2 1e-06 
0.944444444444 1.23232323232 0 1.2 1e-06 
1.0 1.23232323232 0 1.2 1e-06 
0.5 1.27272727273 0 1.2 1e-06 
0.555555555556 1.27272727273 0 1.2 1e-06 
0.611111111111 1.27272727273 0 1.2 1e-06 
0.666666666667 1.27272727273 0 1.2 1e-06 
0.722222222222 1.27272727273 0 1.2 1e-06 
0.777777777778 1.27272727273 0 1.2 1e-06 
0.833333333333 1.27272727273 0 1.2 1e-06 
0.888888888889 1.27272727273 0 1.2 1e-06 
0.944444444444 1.27272727273 0 1.2 1e-06 
1.0 1.27272727273 0 1.2 1e-06 
0.5 1.31313131313 0 1.2 1e-06 
0.555555555556 1.31313131313 0 1.2 1e-06 
0.611111111111 1.31313131313 0 1.2 1e-06 
0.666666666667 1.31313131313 0 1.2 1e-06 
0.722222222222 1.31313131313 0 1.2 1e-06 
0.777777777778 1.31313131313 0 1.2 1e-06 
0.833333333333 1.31313131313 0 1.2 1e-06 
0.888888888889 1.31313131313 0 1.2 1e-06 
0.944444444444 1.31313131313 0 1.2 1e-06 
1.0 1.31313131313 0 1.2 1e-06 
0.5 1.35353535354 0 1.2 1e-06 
0.555555555556 1.35353535354 0 1.2 1e-06 
0.611111111111 1.35353535354 0 1.2 1e-06 
0.666666666667 1.35353535354 0 1.2 1e-06 
0.722222222222 1.35353535354 0 1.2 1e-06 
0.777777777778 1.35353535354 0 1.2 1e-06 
0.833333333333 1.35353535354 0 1.2 1e-06 
0.888888888889 1.35353535354 0 1.2 1e-06 
0.944444444444 1.35353535354 0 1.2 1e-06 
1.0 1.35353535354 0 1.2 1e-06 
0.5 1.39393939394 0 1.2 1e-06 
0.555555555556 1.39393939394 0 1.2 1e-06 
0.611111111111 1.39393939394 0 1.2 1e-06 
0.666666666667 1.39393939394 0 1.2 1e-06 
0.722222222222 1.39393939394 0 1.2 1e-06 
0.777777777778 1.39393939394 0 1.2 1e-06 
0.833333333333 1.39393939394 0 1.2 1e-06 
0.888888888889 1.39393939394 0 1.2 1e-06 
0.944444444444 1.39393939394 0 1.2 1e-06 
1.0 1.39393939394 0 1.2 1e-06 
0.5 1.43434343434 0 1.2 1e-06 
0.555555555556 1.43434343434 0 1.2 1e-06 
0.611111111111 1.43434343434 0 1.2 1e-06 
0.666666666667 1.43434343434 0 1.2 1e-06 
0.722222222222 1.43434343434 0 1.2 1e-06 
0.777777777778 1.43434343434 0 1.2 1e-06 
0.833333333333 1.43434343434 0 1.2 1e-06 
0.888888888889 1.43434343434 0 1.2 1e-06 
0.944444444444 1.43434343434 0 1.2 1e-06 
1.0 1.43434343434 0 1.2 1e-06 
0.5 1.47474747475 0 1.2 1e-06 
0.555555555556 1.47474747475 0 1.2 1e-06 
0.611111111111 1.47474747475 0 1.2 1e-06 
0.666666666667 1.47474747475 0 1.2 1e-06 
0.722222222222 1.47474747475 0 1.2 1e-06 
0.777777777778 1.47474747475 0 1.2 1e-06 
0.833333333333 1.47474747475 0 1.2 1e-06 
0.888888888889 1.47474747475 0 1.2 1e-06 
0.944444444444 1.47474747475 0 1.2 1e-06 
1.0 1.47474747475 0 1.2 1e-06 
0.5 1.51515151515 0 1.2 1e-06 
0.555555555556 1.51515151515 0 1.2 1e-06 
0.611111111111 1.51515151515 0 1.2 1e-06 
0.666666666667 1.51515151515 0 1.2 1e-06 
0.722222222222 1.51515151515 0 1.2 1e-06 
0.777777777778 1.51515151515 0 1.2 1e-06 
0.833333333333 1.51515151515 0 1.2 1e-06 
0.888888888889 1.51515151515 0 1.2 1e-06 
0.944444444444 1.51515151515 0 1.2 1e-06 
1.0 1.51515151515 0 1.2 1e-06 
0.5 1.55555555556 0 1.2 1e-06 
0.555555555556 1.55555555556 0 1.2 1e-06 
0.611111111111 1.55555555556 0 1.2 1e-06 
0.666666666667 1.55555555556 0 1.2 1e-06 
0.722222222222 1.55555555556 0 1.2 1e-06 
0.777777777778 1.55555555556 0 1.2 1e-06 
0.833333333333 1.55555555556 0 1.2 1e-06 
0.888888888889 1.55555555556 0 1.2 1e-06 
0.944444444444 1.55555555556 0 1.2 1e-06 
1.0 1.55555555556 0 1.2 1e-06 
0.5 1.59595959596 0 1.2 1e-06 
0.555555555556 1.59595959596 0 1.2 1e-06 
0.611111111111 1.59595959596 0 1.2 1e-06 
0.666666666667 1.59595959596 0 1.2 1e-06 
0.722222222222 1.59595959596 0 1.2 1e-06 
0.777777777778 1.59595959596 0 1.2 1e-06 
0.833333333333 1.59595959596 0 1.2 1e-06 
0.888888888889 1.59595959596 0 1.2 1e-06 
0.944444444444 1.59595959596 0 1.2 1e-06 
1.0 1.59595959596 0 1.2 1e-06 
0.5 1.63636363636 0 1.2 1e-06 
0.555555555556 1.63636363636 0 1.2 1e-06 
0.611111111111 1.63636363636 0 1.2 1e-06 
0.666666666667 1.63636363636 0 1.2 1e-06 
0.722222222222 1.63636363636 0 1.2 1e-06 
0.777777777778 1.63636363636 0 1.2 1e-06 
0.833333333333 1.63636363636 0 1.2 1e-06 
0.888888888889 1.63636363636 0 1.2 1e-06 
0.944444444444 1.63636363636 0 1.2 1e-06 
1.0 1.63636363636 0 1.2 1e-06 
0.5 1.67676767677 0 1.2 1e-06 
0.555555555556 1.67676767677 0 1.2 1e-06 
0.611111111111 1.67676767677 0 1.2 1e-06 
0.666666666667 1.67676767677 0 1.2 1e-06 
0.722222222222 1.67676767677 0 1.2 1e-06 
0.777777777778 1.67676767677 0 1.2 1e-06 
0.833333333333 1.67676767677 0 1.2 1e-06 
0.888888888889 1.67676767677 0 1.2 1e-06 
0.944444444444 1.67676767677 0 1.2 1e-06 
1.0 1.67676767677 0 1.2 1e-06 
0.5 1.71717171717 0 1.2 1e-06 
0.555555555556 1.71717171717 0 1.2 1e-06 
0.611111111111 1.71717171717 0 1.2 1e-06 
0.666666666667 1.71717171717 0 1.2 1e-06 
0.722222222222 1.71717171717 0 1.2 1e-06 
0.777777777778 1.71717171717 0 1.2 1e-06 
0.833333333333 1.71717171717 0 1.2 1e-06 
0.888888888889 1.71717171717 0 1.2 1e-06 
0.944444444444 1.71717171717 0 1.2 1e-06 
1.0 1.71717171717 0 1.2 1e-06 
0.5 1.75757575758 0 1.2 1e-06 
0.555555555556 1.75757575758 0 1.2 1e-06 
0.611111111111 1.75757575758 0 1.2 1e-06 
0.666666666667 1.75757575758 0 1.2 1e-06 
0.722222222222 1.75757575758 0 1.2 1e-06 
0.777777777778 1.75757575758 0 1.2 1e-06 
0.833333333333 1.75757575758 0 1.2 1e-06 
0.888888888889 1.75757575758 0 1.2 1e-06 
0.944444444444 1.75757575758 0 1.2 1e-06 
1.0 1.75757575758 0 1.2 1e-06 
0.5 1.79797979798 0 1.2 1e-06 
0.555555555556 1.79797979798 0 1.2 1e-06 
0.611111111111 1.79797979798 0 1.2 1e-06 
0.666666666667 1.79797979798 0 1.2 1e-06 
0.722222222222 1.79797979798 0 1.2 1e-06 
0.777777777778 1.79797979798 0 1.2 1e-06 
0.833333333333 1.79797979798 0 1.2 1e-06 
0.888888888889 1.79797979798 0 1.2 1e-06 
0.944444444444 1.79797979798 0 1.2 1e-06 
1.0 1.79797979798 0 1.2 1e-06 
0.5 1.83838383838 0 1.2 1e-06 
0.555555555556 1.83838383838 0 1.2 1e-06 
0.611111111111 1.83838383838 0 1.2 1e-06 
0.666666666667 1.83838383838 0 1.2 1e-06 
0.722222222222 1.83838383838 0 1.2 1e-06 
0.777777777778 1.83838383838 0 1.2 1e-06 
0.833333333333 1.83838383838 0 1.2 1e-06 
0.888888888889 1.83838383838 0 1.2 1e-06 
0.944444444444 1.83838383838 0 1.2 1e-06 
1.0 1.83838383838 0 1.2 1e-06 
0.5 1.87878787879 0 1.2 1e-06 
0.555555555556 1.87878787879 0 1.2 1e-06 
0.611111111111 1.87878787879 0 1.2 1e-06 
0.666666666667 1.87878787879 0 1.2 1e-06 
0.722222222222 1.87878787879 0 1.2 1e-06 
0.777777777778 1.87878787879 0 1.2 1e-06 
0.833333333333 1.87878787879 0 1.2 1e-06 
0.888888888889 1.87878787879 0 1.2 1e-06 
0.944444444444 1.87878787879 0 1.2 1e-06 
1.0 1.87878787879 0 1.2 1e-06 
0.5 1.91919191919 0 1.2 1e-06 
0.555555555556 1.91919191919 0 1.2 1e-06 
0.611111111111 1.91919191919 0 1.2 1e-06 
0.666666666667 1.91919191919 0 1.2 1e-06 
0.722222222222 1.91919191919 0 1.2 1e-06 
0.777777777778 1.91919191919 0 1.2 1e-06 
0.833333333333 1.91919191919 0 1.2 1e-06 
0.888888888889 1.91919191919 0 1.2 1e-06 
0.944444444444 1.91919191919 0 1.2 1e-06 
1.0 1.91919191919 0 1.2 1e-06 
0.5 1.9595959596 0 1.2 1e-06 
0.555555555556 1.9595959596 0 1.2 1e-06 
0.611111111111 1.9595959596 0 1.2 1e-06 
0.666666666667 1.9595959596 0 1.2 1e-06 
0.722222222222 1.9595959596 0 1.2 1e-06 
0.777777777778 1.9595959596 0 1.2 1e-06 
0.833333333333 1.9595959596 0 1.2 1e-06 
0.888888888889 1.9595959596 0 1.2 1e-06 
0.944444444444 1.9595959596 0 1.2 1e-06 
1.0 1.9595959596 0 1.2 1e-06 
0.5 2.0 0 1.2 1e-06 
0.555555555556 2.0 0 1.2 1e-06 
0.611111111111 2.0 0 1.2 1e-06 
0.666666666667 2.0 0 1.2 1e-06 
0.722222222222 2.0 0 1.2 1e-06 
0.777777777778 2.0 0 1.2 1e-06 
0.833333333333 2.0 0 1.2 1e-06 
0.888888888889 2.0 0 1.2 1e-06 
0.944444444444 2.0 0 1.2 1e-06 
1.0 2.0 0 1.2 1e-06 
0.5 -2.0 0 1.6 1e-06 
0.555555555556 -2.0 0 1.6 1e-06 
0.611111111111 -2.0 0 1.6 1e-06 
0.666666666667 -2.0 0 1.6 1e-06 
0.722222222222 -2.0 0 1.6 1e-06 
0.777777777778 -2.0 0 1.6 1e-06 
0.833333333333 -2.0 0 1.6 1e-06 
0.888888888889 -2.0 0 1.6 1e-06 
0.944444444444 -2.0 0 1.6 1e-06 
1.0 -2.0 0 1.6 1e-06 
0.5 -1.9595959596 0 1.6 1e-06 
0.555555555556 -1.9595959596 0 1.6 1e-06 
0.611111111111 -1.9595959596 0 1.6 1e-06 
0.666666666667 -1.9595959596 0 1.6 1e-06 
0.722222222222 -1.9595959596 0 1.6 1e-06 
0.777777777778 -1.9595959596 0 1.6 1e-06 
0.833333333333 -1.9595959596 0 1.6 1e-06 
0.888888888889 -1.9595959596 0 1.6 1e-06 
0.944444444444 -1.9595959596 0 1.6 1e-06 
1.0 -1.9595959596 0 1.6 1e-06 
0.5 -1.91919191919 0 1.6 1e-06 
0.555555555556 -1.91919191919 0 1.6 1e-06 
0.611111111111 -1.91919191919 0 1.6 1e-06 
0.666666666667 -1.91919191919 0 1.6 1e-06 
0.722222222222 -1.91919191919 0 1.6 1e-06 
0.777777777778 -1.91919191919 0 1.6 1e-06 
0.833333333333 -1.91919191919 0 1.6 1e-06 
0.888888888889 -1.91919191919 0 1.6 1e-06 
0.944444444444 -1.91919191919 0 1.6 1e-06 
1.0 -1.91919191919 0 1.6 1e-06 
0.5 -1.87878787879 0 1.6 1e-06 
0.555555555556 -1.87878787879 0 1.6 1e-06 
0.611111111111 -1.87878787879 0 1.6 1e-06 
0.666666666667 -1.87878787879 0 1.6 1e-06 
0.722222222222 -1.87878787879 0 1.6 1e-06 
0.777777777778 -1.87878787879 0 1.6 1e-06 
0.833333333333 -1.87878787879 0 1.6 1e-06 
0.888888888889 -1.87878787879 0 1.6 1e-06 
0.944444444444 -1.87878787879 0 1.6 1e-06 
1.0 -1.87878787879 0 1.6 1e-06 
0.5 -1.83838383838 0 1.6 1e-06 
0.555555555556 -1.83838383838 0 1.6 1e-06 
0.611111111111 -1.83838383838 0 1.6 1e-06 
0.666666666667 -1.83838383838 0 1.6 1e-06 
0.722222222222 -1.83838383838 0 1.6 1e-06 
0.777777777778 -1.83838383838 0 1.6 1e-06 
0.833333333333 -1.83838383838 0 1.6 1e-06 
0.888888888889 -1.83838383838 0 1.6 1e-06 
0.944444444444 -1.83838383838 0 1.6 1e-06 
1.0 -1.83838383838 0 1.6 1e-06 
0.5 -1.79797979798 0 1.6 1e-06 
0.555555555556 -1.79797979798 0 1.6 1e-06 
0.611111111111 -1.79797979798 0 1.6 1e-06 
0.666666666667 -1.79797979798 0 1.6 1e-06 
0.722222222222 -1.79797979798 0 1.6 1e-06 
0.777777777778 -1.79797979798 0 1.6 1e-06 
0.833333333333 -1.79797979798 0 1.6 1e-06 
0.888888888889 -1.79797979798 0 1.6 1e-06 
0.944444444444 -1.79797979798 0 1.6 1e-06 
1.0 -1.79797979798 0 1.6 1e-06 
0.5 -1.75757575758 0 1.6 1e-06 
0.555555555556 -1.75757575758 0 1.6 1e-06 
0.611111111111 -1.75757575758 0 1.6 1e-06 
0.666666666667 -1.75757575758 0 1.6 1e-06 
0.722222222222 -1.75757575758 0 1.6 1e-06 
0.777777777778 -1.75757575758 0 1.6 1e-06 
0.833333333333 -1.75757575758 0 1.6 1e-06 
0.888888888889 -1.75757575758 0 1.6 1e-06 
0.944444444444 -1.75757575758 0 1.6 1e-06 
1.0 -1.75757575758 0 1.6 1e-06 
0.5 -1.71717171717 0 1.6 1e-06 
0.555555555556 -1.71717171717 0 1.6 1e-06 
0.611111111111 -1.71717171717 0 1.6 1e-06 
0.666666666667 -1.71717171717 0 1.6 1e-06 
0.722222222222 -1.71717171717 0 1.6 1e-06 
0.777777777778 -1.71717171717 0 1.6 1e-06 
0.833333333333 -1.71717171717 0 1.6 1e-06 
0.888888888889 -1.71717171717 0 1.6 1e-06 
0.944444444444 -1.71717171717 0 1.6 1e-06 
1.0 -1.71717171717 0 1.6 1e-06 
0.5 -1.67676767677 0 1.6 1e-06 
0.555555555556 -1.67676767677 0 1.6 1e-06 
0.611111111111 -1.67676767677 0 1.6 1e-06 
0.666666666667 -1.67676767677 0 1.6 1e-06 
0.722222222222 -1.67676767677 0 1.6 1e-06 
0.777777777778 -1.67676767677 0 1.6 1e-06 
0.833333333333 -1.67676767677 0 1.6 1e-06 
0.888888888889 -1.67676767677 0 1.6 1e-06 
0.944444444444 -1.67676767677 0 1.6 1e-06 
1.0 -1.67676767677 0 1.6 1e-06 
0.5 -1.63636363636 0 1.6 1e-06 
0.555555555556 -1.63636363636 0 1.6 1e-06 
0.611111111111 -1.63636363636 0 1.6 1e-06 
0.666666666667 -1.63636363636 0 1.6 1e-06 
0.722222222222 -1.63636363636 0 1.6 1e-06 
0.777777777778 -1.63636363636 0 1.6 1e-06 
0.833333333333 -1.63636363636 0 1.6 1e-06 
0.888888888889 -1.63636363636 0 1.6 1e-06 
0.944444444444 -1.63636363636 0 1.6 1e-06 
1.0 -1.63636363636 0 1.6 1e-06 
0.5 -1.59595959596 0 1.6 1e-06 
0.555555555556 -1.59595959596 0 1.6 1e-06 
0.611111111111 -1.59595959596 0 1.6 1e-06 
0.666666666667 -1.59595959596 0 1.6 1e-06 
0.722222222222 -1.59595959596 0 1.6 1e-06 
0.777777777778 -1.59595959596 0 1.6 1e-06 
0.833333333333 -1.59595959596 0 1.6 1e-06 
0.888888888889 -1.59595959596 0 1.6 1e-06 
0.944444444444 -1.59595959596 0 1.6 1e-06 
1.0 -1.59595959596 0 1.6 1e-06 
0.5 -1.55555555556 0 1.6 1e-06 
0.555555555556 -1.55555555556 0 1.6 1e-06 
0.611111111111 -1.55555555556 0 1.6 1e-06 
0.666666666667 -1.55555555556 0 1.6 1e-06 
0.722222222222 -1.55555555556 0 1.6 1e-06 
0.777777777778 -1.55555555556 0 1.6 1e-06 
0.833333333333 -1.55555555556 0 1.6 1e-06 
0.888888888889 -1.55555555556 0 1.6 1e-06 
0.944444444444 -1.55555555556 0 1.6 1e-06 
1.0 -1.55555555556 0 1.6 1e-06 
0.5 -1.51515151515 0 1.6 1e-06 
0.555555555556 -1.51515151515 0 1.6 1e-06 
0.611111111111 -1.51515151515 0 1.6 1e-06 
0.666666666667 -1.51515151515 0 1.6 1e-06 
0.722222222222 -1.51515151515 0 1.6 1e-06 
0.777777777778 -1.51515151515 0 1.6 1e-06 
0.833333333333 -1.51515151515 0 1.6 1e-06 
0.888888888889 -1.51515151515 0 1.6 1e-06 
0.944444444444 -1.51515151515 0 1.6 1e-06 
1.0 -1.51515151515 0 1.6 1e-06 
0.5 -1.47474747475 0 1.6 1e-06 
0.555555555556 -1.47474747475 0 1.6 1e-06 
0.611111111111 -1.47474747475 0 1.6 1e-06 
0.666666666667 -1.47474747475 0 1.6 1e-06 
0.722222222222 -1.47474747475 0 1.6 1e-06 
0.777777777778 -1.47474747475 0 1.6 1e-06 
0.833333333333 -1.47474747475 0 1.6 1e-06 
0.888888888889 -1.47474747475 0 1.6 1e-06 
0.944444444444 -1.47474747475 0 1.6 1e-06 
1.0 -1.47474747475 0 1.6 1e-06 
0.5 -1.43434343434 0 1.6 1e-06 
0.555555555556 -1.43434343434 0 1.6 1e-06 
0.611111111111 -1.43434343434 0 1.6 1e-06 
0.666666666667 -1.43434343434 0 1.6 1e-06 
0.722222222222 -1.43434343434 0 1.6 1e-06 
0.777777777778 -1.43434343434 0 1.6 1e-06 
0.833333333333 -1.43434343434 0 1.6 1e-06 
0.888888888889 -1.43434343434 0 1.6 1e-06 
0.944444444444 -1.43434343434 0 1.6 1e-06 
1.0 -1.43434343434 0 1.6 1e-06 
0.5 -1.39393939394 0 1.6 1e-06 
0.555555555556 -1.39393939394 0 1.6 1e-06 
0.611111111111 -1.39393939394 0 1.6 1e-06 
0.666666666667 -1.39393939394 0 1.6 1e-06 
0.722222222222 -1.39393939394 0 1.6 1e-06 
0.777777777778 -1.39393939394 0 1.6 1e-06 
0.833333333333 -1.39393939394 0 1.6 1e-06 
0.888888888889 -1.39393939394 0 1.6 1e-06 
0.944444444444 -1.39393939394 0 1.6 1e-06 
1.0 -1.39393939394 0 1.6 1e-06 
0.5 -1.35353535354 0 1.6 1e-06 
0.555555555556 -1.35353535354 0 1.6 1e-06 
0.611111111111 -1.35353535354 0 1.6 1e-06 
0.666666666667 -1.35353535354 0 1.6 1e-06 
0.722222222222 -1.35353535354 0 1.6 1e-06 
0.777777777778 -1.35353535354 0 1.6 1e-06 
0.833333333333 -1.35353535354 0 1.6 1e-06 
0.888888888889 -1.35353535354 0 1.6 1e-06 
0.944444444444 -1.35353535354 0 1.6 1e-06 
1.0 -1.35353535354 0 1.6 1e-06 
0.5 -1.31313131313 0 1.6 1e-06 
0.555555555556 -1.31313131313 0 1.6 1e-06 
0.611111111111 -1.31313131313 0 1.6 1e-06 
0.666666666667 -1.31313131313 0 1.6 1e-06 
0.722222222222 -1.31313131313 0 1.6 1e-06 
0.777777777778 -1.31313131313 0 1.6 1e-06 
0.833333333333 -1.31313131313 0 1.6 1e-06 
0.888888888889 -1.31313131313 0 1.6 1e-06 
0.944444444444 -1.31313131313 0 1.6 1e-06 
1.0 -1.31313131313 0 1.6 1e-06 
0.5 -1.27272727273 0 1.6 1e-06 
0.555555555556 -1.27272727273 0 1.6 1e-06 
0.611111111111 -1.27272727273 0 1.6 1e-06 
0.666666666667 -1.27272727273 0 1.6 1e-06 
0.722222222222 -1.27272727273 0 1.6 1e-06 
0.777777777778 -1.27272727273 0 1.6 1e-06 
0.833333333333 -1.27272727273 0 1.6 1e-06 
0.888888888889 -1.27272727273 0 1.6 1e-06 
0.944444444444 -1.27272727273 0 1.6 1e-06 
1.0 -1.27272727273 0 1.6 1e-06 
0.5 -1.23232323232 0 1.6 1e-06 
0.555555555556 -1.23232323232 0 1.6 1e-06 
0.611111111111 -1.23232323232 0 1.6 1e-06 
0.666666666667 -1.23232323232 0 1.6 1e-06 
0.722222222222 -1.23232323232 0 1.6 1e-06 
0.777777777778 -1.23232323232 0 1.6 1e-06 
0.833333333333 -1.23232323232 0 1.6 1e-06 
0.888888888889 -1.23232323232 0 1.6 1e-06 
0.944444444444 -1.23232323232 0 1.6 1e-06 
1.0 -1.23232323232 0 1.6 1e-06 
0.5 -1.19191919192 0 1.6 1e-06 
0.555555555556 -1.19191919192 0 1.6 1e-06 
0.611111111111 -1.19191919192 0 1.6 1e-06 
0.666666666667 -1.19191919192 0 1.6 1e-06 
0.722222222222 -1.19191919192 0 1.6 1e-06 
0.777777777778 -1.19191919192 0 1.6 1e-06 
0.833333333333 -1.19191919192 0 1.6 1e-06 
0.888888888889 -1.19191919192 0 1.6 1e-06 
0.944444444444 -1.19191919192 0 1.6 1e-06 
1.0 -1.19191919192 0 1.6 1e-06 
0.5 -1.15151515152 0 1.6 1e-06 
0.555555555556 -1.15151515152 0 1.6 1e-06 
0.611111111111 -1.15151515152 0 1.6 1e-06 
0.666666666667 -1.15151515152 0 1.6 1e-06 
0.722222222222 -1.15151515152 0 1.6 1e-06 
0.777777777778 -1.15151515152 0 1.6 1e-06 
0.833333333333 -1.15151515152 0 1.6 1e-06 
0.888888888889 -1.15151515152 0 1.6 1e-06 
0.944444444444 -1.15151515152 0 1.6 1e-06 
1.0 -1.15151515152 0 1.6 1e-06 
0.5 -1.11111111111 0 1.6 1e-06 
0.555555555556 -1.11111111111 0 1.6 1e-06 
0.611111111111 -1.11111111111 0 1.6 1e-06 
0.666666666667 -1.11111111111 0 1.6 1e-06 
0.722222222222 -1.11111111111 0 1.6 1e-06 
0.777777777778 -1.11111111111 0 1.6 1e-06 
0.833333333333 -1.11111111111 0 1.6 1e-06 
0.888888888889 -1.11111111111 0 1.6 1e-06 
0.944444444444 -1.11111111111 0 1.6 1e-06 
1.0 -1.11111111111 0 1.6 1e-06 
0.5 -1.07070707071 0 1.6 1e-06 
0.555555555556 -1.07070707071 0 1.6 1e-06 
0.611111111111 -1.07070707071 0 1.6 1e-06 
0.666666666667 -1.07070707071 0 1.6 1e-06 
0.722222222222 -1.07070707071 0 1.6 1e-06 
0.777777777778 -1.07070707071 0 1.6 1e-06 
0.833333333333 -1.07070707071 0 1.6 1e-06 
0.888888888889 -1.07070707071 0 1.6 1e-06 
0.944444444444 -1.07070707071 0 1.6 1e-06 
1.0 -1.07070707071 0 1.6 1e-06 
0.5 -1.0303030303 0 1.6 1e-06 
0.555555555556 -1.0303030303 0 1.6 1e-06 
0.611111111111 -1.0303030303 0 1.6 1e-06 
0.666666666667 -1.0303030303 0 1.6 1e-06 
0.722222222222 -1.0303030303 0 1.6 1e-06 
0.777777777778 -1.0303030303 0 1.6 1e-06 
0.833333333333 -1.0303030303 0 1.6 1e-06 
0.888888888889 -1.0303030303 0 1.6 1e-06 
0.944444444444 -1.0303030303 0 1.6 1e-06 
1.0 -1.0303030303 0 1.6 1e-06 
0.5 -0.989898989899 0 1.6 1e-06 
0.555555555556 -0.989898989899 0 1.6 1e-06 
0.611111111111 -0.989898989899 0 1.6 1e-06 
0.666666666667 -0.989898989899 0 1.6 1e-06 
0.722222222222 -0.989898989899 0 1.6 1e-06 
0.777777777778 -0.989898989899 0 1.6 1e-06 
0.833333333333 -0.989898989899 0 1.6 1e-06 
0.888888888889 -0.989898989899 0 1.6 1e-06 
0.944444444444 -0.989898989899 0 1.6 1e-06 
1.0 -0.989898989899 0 1.6 1e-06 
0.5 -0.949494949495 0 1.6 1e-06 
0.555555555556 -0.949494949495 0 1.6 1e-06 
0.611111111111 -0.949494949495 0 1.6 1e-06 
0.666666666667 -0.949494949495 0 1.6 1e-06 
0.722222222222 -0.949494949495 0 1.6 1e-06 
0.777777777778 -0.949494949495 0 1.6 1e-06 
0.833333333333 -0.949494949495 0 1.6 1e-06 
0.888888888889 -0.949494949495 0 1.6 1e-06 
0.944444444444 -0.949494949495 0 1.6 1e-06 
1.0 -0.949494949495 0 1.6 1e-06 
0.5 -0.909090909091 0 1.6 1e-06 
0.555555555556 -0.909090909091 0 1.6 1e-06 
0.611111111111 -0.909090909091 0 1.6 1e-06 
0.666666666667 -0.909090909091 0 1.6 1e-06 
0.722222222222 -0.909090909091 0 1.6 1e-06 
0.777777777778 -0.909090909091 0 1.6 1e-06 
0.833333333333 -0.909090909091 0 1.6 1e-06 
0.888888888889 -0.909090909091 0 1.6 1e-06 
0.944444444444 -0.909090909091 0 1.6 1e-06 
1.0 -0.909090909091 0 1.6 1e-06 
0.5 -0.868686868687 0 1.6 1e-06 
0.555555555556 -0.868686868687 0 1.6 1e-06 
0.611111111111 -0.868686868687 0 1.6 1e-06 
0.666666666667 -0.868686868687 0 1.6 1e-06 
0.722222222222 -0.868686868687 0 1.6 1e-06 
0.777777777778 -0.868686868687 0 1.6 1e-06 
0.833333333333 -0.868686868687 0 1.6 1e-06 
0.888888888889 -0.868686868687 0 1.6 1e-06 
0.944444444444 -0.868686868687 0 1.6 1e-06 
1.0 -0.868686868687 0 1.6 1e-06 
0.5 -0.828282828283 0 1.6 1e-06 
0.555555555556 -0.828282828283 0 1.6 1e-06 
0.611111111111 -0.828282828283 0 1.6 1e-06 
0.666666666667 -0.828282828283 0 1.6 1e-06 
0.722222222222 -0.828282828283 0 1.6 1e-06 
0.777777777778 -0.828282828283 0 1.6 1e-06 
0.833333333333 -0.828282828283 0 1.6 1e-06 
0.888888888889 -0.828282828283 0 1.6 1e-06 
0.944444444444 -0.828282828283 0 1.6 1e-06 
1.0 -0.828282828283 0 1.6 1e-06 
0.5 -0.787878787879 0 1.6 1e-06 
0.555555555556 -0.787878787879 0 1.6 1e-06 
0.611111111111 -0.787878787879 0 1.6 1e-06 
0.666666666667 -0.787878787879 0 1.6 1e-06 
0.722222222222 -0.787878787879 0 1.6 1e-06 
0.777777777778 -0.787878787879 0 1.6 1e-06 
0.833333333333 -0.787878787879 0 1.6 1e-06 
0.888888888889 -0.787878787879 0 1.6 1e-06 
0.944444444444 -0.787878787879 0 1.6 1e-06 
1.0 -0.787878787879 0 1.6 1e-06 
0.5 -0.747474747475 0 1.6 1e-06 
0.555555555556 -0.747474747475 0 1.6 1e-06 
0.611111111111 -0.747474747475 0 1.6 1e-06 
0.666666666667 -0.747474747475 0 1.6 1e-06 
0.722222222222 -0.747474747475 0 1.6 1e-06 
0.777777777778 -0.747474747475 0 1.6 1e-06 
0.833333333333 -0.747474747475 0 1.6 1e-06 
0.888888888889 -0.747474747475 0 1.6 1e-06 
0.944444444444 -0.747474747475 0 1.6 1e-06 
1.0 -0.747474747475 0 1.6 1e-06 
0.5 -0.707070707071 0 1.6 1e-06 
0.555555555556 -0.707070707071 0 1.6 1e-06 
0.611111111111 -0.707070707071 0 1.6 1e-06 
0.666666666667 -0.707070707071 0 1.6 1e-06 
0.722222222222 -0.707070707071 0 1.6 1e-06 
0.777777777778 -0.707070707071 0 1.6 1e-06 
0.833333333333 -0.707070707071 0 1.6 1e-06 
0.888888888889 -0.707070707071 0 1.6 1e-06 
0.944444444444 -0.707070707071 0 1.6 1e-06 
1.0 -0.707070707071 0 1.6 1e-06 
0.5 -0.666666666667 0 1.6 1e-06 
0.555555555556 -0.666666666667 0 1.6 1e-06 
0.611111111111 -0.666666666667 0 1.6 1e-06 
0.666666666667 -0.666666666667 0 1.6 1e-06 
0.722222222222 -0.666666666667 0 1.6 1e-06 
0.777777777778 -0.666666666667 0 1.6 1e-06 
0.833333333333 -0.666666666667 0 1.6 1e-06 
0.888888888889 -0.666666666667 0 1.6 1e-06 
0.944444444444 -0.666666666667 0 1.6 1e-06 
1.0 -0.666666666667 0 1.6 1e-06 
0.5 -0.626262626263 0 1.6 1e-06 
0.555555555556 -0.626262626263 0 1.6 1e-06 
0.611111111111 -0.626262626263 0 1.6 1e-06 
0.666666666667 -0.626262626263 0 1.6 1e-06 
0.722222222222 -0.626262626263 0 1.6 1e-06 
0.777777777778 -0.626262626263 0 1.6 1e-06 
0.833333333333 -0.626262626263 0 1.6 1e-06 
0.888888888889 -0.626262626263 0 1.6 1e-06 
0.944444444444 -0.626262626263 0 1.6 1e-06 
1.0 -0.626262626263 0 1.6 1e-06 
0.5 -0.585858585859 0 1.6 1e-06 
0.555555555556 -0.585858585859 0 1.6 1e-06 
0.611111111111 -0.585858585859 0 1.6 1e-06 
0.666666666667 -0.585858585859 0 1.6 1e-06 
0.722222222222 -0.585858585859 0 1.6 1e-06 
0.777777777778 -0.585858585859 0 1.6 1e-06 
0.833333333333 -0.585858585859 0 1.6 1e-06 
0.888888888889 -0.585858585859 0 1.6 1e-06 
0.944444444444 -0.585858585859 0 1.6 1e-06 
1.0 -0.585858585859 0 1.6 1e-06 
0.5 -0.545454545455 0 1.6 1e-06 
0.555555555556 -0.545454545455 0 1.6 1e-06 
0.611111111111 -0.545454545455 0 1.6 1e-06 
0.666666666667 -0.545454545455 0 1.6 1e-06 
0.722222222222 -0.545454545455 0 1.6 1e-06 
0.777777777778 -0.545454545455 0 1.6 1e-06 
0.833333333333 -0.545454545455 0 1.6 1e-06 
0.888888888889 -0.545454545455 0 1.6 1e-06 
0.944444444444 -0.545454545455 0 1.6 1e-06 
1.0 -0.545454545455 0 1.6 1e-06 
0.5 -0.505050505051 0 1.6 1e-06 
0.555555555556 -0.505050505051 0 1.6 1e-06 
0.611111111111 -0.505050505051 0 1.6 1e-06 
0.666666666667 -0.505050505051 0 1.6 1e-06 
0.722222222222 -0.505050505051 0 1.6 1e-06 
0.777777777778 -0.505050505051 0 1.6 1e-06 
0.833333333333 -0.505050505051 0 1.6 1e-06 
0.888888888889 -0.505050505051 0 1.6 1e-06 
0.944444444444 -0.505050505051 0 1.6 1e-06 
1.0 -0.505050505051 0 1.6 1e-06 
0.5 -0.464646464646 0 1.6 1e-06 
0.555555555556 -0.464646464646 0 1.6 1e-06 
0.611111111111 -0.464646464646 0 1.6 1e-06 
0.666666666667 -0.464646464646 0 1.6 1e-06 
0.722222222222 -0.464646464646 0 1.6 1e-06 
0.777777777778 -0.464646464646 0 1.6 1e-06 
0.833333333333 -0.464646464646 0 1.6 1e-06 
0.888888888889 -0.464646464646 0 1.6 1e-06 
0.944444444444 -0.464646464646 0 1.6 1e-06 
1.0 -0.464646464646 0 1.6 1e-06 
0.5 -0.424242424242 0 1.6 1e-06 
0.555555555556 -0.424242424242 0 1.6 1e-06 
0.611111111111 -0.424242424242 0 1.6 1e-06 
0.666666666667 -0.424242424242 0 1.6 1e-06 
0.722222222222 -0.424242424242 0 1.6 1e-06 
0.777777777778 -0.424242424242 0 1.6 1e-06 
0.833333333333 -0.424242424242 0 1.6 1e-06 
0.888888888889 -0.424242424242 0 1.6 1e-06 
0.944444444444 -0.424242424242 0 1.6 1e-06 
1.0 -0.424242424242 0 1.6 1e-06 
0.5 -0.383838383838 0 1.6 1e-06 
0.555555555556 -0.383838383838 0 1.6 1e-06 
0.611111111111 -0.383838383838 0 1.6 1e-06 
0.666666666667 -0.383838383838 0 1.6 1e-06 
0.722222222222 -0.383838383838 0 1.6 1e-06 
0.777777777778 -0.383838383838 0 1.6 1e-06 
0.833333333333 -0.383838383838 0 1.6 1e-06 
0.888888888889 -0.383838383838 0 1.6 1e-06 
0.944444444444 -0.383838383838 0 1.6 1e-06 
1.0 -0.383838383838 0 1.6 1e-06 
0.5 -0.343434343434 0 1.6 1e-06 
0.555555555556 -0.343434343434 0 1.6 1e-06 
0.611111111111 -0.343434343434 0 1.6 1e-06 
0.666666666667 -0.343434343434 0 1.6 1e-06 
0.722222222222 -0.343434343434 0 1.6 1e-06 
0.777777777778 -0.343434343434 0 1.6 1e-06 
0.833333333333 -0.343434343434 0 1.6 1e-06 
0.888888888889 -0.343434343434 0 1.6 1e-06 
0.944444444444 -0.343434343434 0 1.6 1e-06 
1.0 -0.343434343434 0 1.6 1e-06 
0.5 -0.30303030303 0 1.6 1e-06 
0.555555555556 -0.30303030303 0 1.6 1e-06 
0.611111111111 -0.30303030303 0 1.6 1e-06 
0.666666666667 -0.30303030303 0 1.6 1e-06 
0.722222222222 -0.30303030303 0 1.6 1e-06 
0.777777777778 -0.30303030303 0 1.6 1e-06 
0.833333333333 -0.30303030303 0 1.6 1e-06 
0.888888888889 -0.30303030303 0 1.6 1e-06 
0.944444444444 -0.30303030303 0 1.6 1e-06 
1.0 -0.30303030303 0 1.6 1e-06 
0.5 -0.262626262626 0 1.6 1e-06 
0.555555555556 -0.262626262626 0 1.6 1e-06 
0.611111111111 -0.262626262626 0 1.6 1e-06 
0.666666666667 -0.262626262626 0 1.6 1e-06 
0.722222222222 -0.262626262626 0 1.6 1e-06 
0.777777777778 -0.262626262626 0 1.6 1e-06 
0.833333333333 -0.262626262626 0 1.6 1e-06 
0.888888888889 -0.262626262626 0 1.6 1e-06 
0.944444444444 -0.262626262626 0 1.6 1e-06 
1.0 -0.262626262626 0 1.6 1e-06 
0.5 -0.222222222222 0 1.6 1e-06 
0.555555555556 -0.222222222222 0 1.6 1e-06 
0.611111111111 -0.222222222222 0 1.6 1e-06 
0.666666666667 -0.222222222222 0 1.6 1e-06 
0.722222222222 -0.222222222222 0 1.6 1e-06 
0.777777777778 -0.222222222222 0 1.6 1e-06 
0.833333333333 -0.222222222222 0 1.6 1e-06 
0.888888888889 -0.222222222222 0 1.6 1e-06 
0.944444444444 -0.222222222222 0 1.6 1e-06 
1.0 -0.222222222222 0 1.6 1e-06 
0.5 -0.181818181818 0 1.6 1e-06 
0.555555555556 -0.181818181818 0 1.6 1e-06 
0.611111111111 -0.181818181818 0 1.6 1e-06 
0.666666666667 -0.181818181818 0 1.6 1e-06 
0.722222222222 -0.181818181818 0 1.6 1e-06 
0.777777777778 -0.181818181818 0 1.6 1e-06 
0.833333333333 -0.181818181818 0 1.6 1e-06 
0.888888888889 -0.181818181818 0 1.6 1e-06 
0.944444444444 -0.181818181818 0 1.6 1e-06 
1.0 -0.181818181818 0 1.6 1e-06 
0.5 -0.141414141414 0 1.6 1e-06 
0.555555555556 -0.141414141414 0 1.6 1e-06 
0.611111111111 -0.141414141414 0 1.6 1e-06 
0.666666666667 -0.141414141414 0 1.6 1e-06 
0.722222222222 -0.141414141414 0 1.6 1e-06 
0.777777777778 -0.141414141414 0 1.6 1e-06 
0.833333333333 -0.141414141414 0 1.6 1e-06 
0.888888888889 -0.141414141414 0 1.6 1e-06 
0.944444444444 -0.141414141414 0 1.6 1e-06 
1.0 -0.141414141414 0 1.6 1e-06 
0.5 -0.10101010101 0 1.6 1e-06 
0.555555555556 -0.10101010101 0 1.6 1e-06 
0.611111111111 -0.10101010101 0 1.6 1e-06 
0.666666666667 -0.10101010101 0 1.6 1e-06 
0.722222222222 -0.10101010101 0 1.6 1e-06 
0.777777777778 -0.10101010101 0 1.6 1e-06 
0.833333333333 -0.10101010101 0 1.6 1e-06 
0.888888888889 -0.10101010101 0 1.6 1e-06 
0.944444444444 -0.10101010101 0 1.6 1e-06 
1.0 -0.10101010101 0 1.6 1e-06 
0.5 -0.0606060606061 0 1.6 1e-06 
0.555555555556 -0.0606060606061 0 1.6 1e-06 
0.611111111111 -0.0606060606061 0 1.6 1e-06 
0.666666666667 -0.0606060606061 0 1.6 1e-06 
0.722222222222 -0.0606060606061 0 1.6 1e-06 
0.777777777778 -0.0606060606061 0 1.6 1e-06 
0.833333333333 -0.0606060606061 0 1.6 1e-06 
0.888888888889 -0.0606060606061 0 1.6 1e-06 
0.944444444444 -0.0606060606061 0 1.6 1e-06 
1.0 -0.0606060606061 0 1.6 1e-06 
0.5 -0.020202020202 0 1.6 1e-06 
0.555555555556 -0.020202020202 0 1.6 1e-06 
0.611111111111 -0.020202020202 0 1.6 1e-06 
0.666666666667 -0.020202020202 0 1.6 1e-06 
0.722222222222 -0.020202020202 0 1.6 1e-06 
0.777777777778 -0.020202020202 0 1.6 1e-06 
0.833333333333 -0.020202020202 0 1.6 1e-06 
0.888888888889 -0.020202020202 0 1.6 1e-06 
0.944444444444 -0.020202020202 0 1.6 1e-06 
1.0 -0.020202020202 0 1.6 1e-06 
0.5 0.020202020202 0 1.6 1e-06 
0.555555555556 0.020202020202 0 1.6 1e-06 
0.611111111111 0.020202020202 0 1.6 1e-06 
0.666666666667 0.020202020202 0 1.6 1e-06 
0.722222222222 0.020202020202 0 1.6 1e-06 
0.777777777778 0.020202020202 0 1.6 1e-06 
0.833333333333 0.020202020202 0 1.6 1e-06 
0.888888888889 0.020202020202 0 1.6 1e-06 
0.944444444444 0.020202020202 0 1.6 1e-06 
1.0 0.020202020202 0 1.6 1e-06 
0.5 0.0606060606061 0 1.6 1e-06 
0.555555555556 0.0606060606061 0 1.6 1e-06 
0.611111111111 0.0606060606061 0 1.6 1e-06 
0.666666666667 0.0606060606061 0 1.6 1e-06 
0.722222222222 0.0606060606061 0 1.6 1e-06 
0.777777777778 0.0606060606061 0 1.6 1e-06 
0.833333333333 0.0606060606061 0 1.6 1e-06 
0.888888888889 0.0606060606061 0 1.6 1e-06 
0.944444444444 0.0606060606061 0 1.6 1e-06 
1.0 0.0606060606061 0 1.6 1e-06 
0.5 0.10101010101 0 1.6 1e-06 
0.555555555556 0.10101010101 0 1.6 1e-06 
0.611111111111 0.10101010101 0 1.6 1e-06 
0.666666666667 0.10101010101 0 1.6 1e-06 
0.722222222222 0.10101010101 0 1.6 1e-06 
0.777777777778 0.10101010101 0 1.6 1e-06 
0.833333333333 0.10101010101 0 1.6 1e-06 
0.888888888889 0.10101010101 0 1.6 1e-06 
0.944444444444 0.10101010101 0 1.6 1e-06 
1.0 0.10101010101 0 1.6 1e-06 
0.5 0.141414141414 0 1.6 1e-06 
0.555555555556 0.141414141414 0 1.6 1e-06 
0.611111111111 0.141414141414 0 1.6 1e-06 
0.666666666667 0.141414141414 0 1.6 1e-06 
0.722222222222 0.141414141414 0 1.6 1e-06 
0.777777777778 0.141414141414 0 1.6 1e-06 
0.833333333333 0.141414141414 0 1.6 1e-06 
0.888888888889 0.141414141414 0 1.6 1e-06 
0.944444444444 0.141414141414 0 1.6 1e-06 
1.0 0.141414141414 0 1.6 1e-06 
0.5 0.181818181818 0 1.6 1e-06 
0.555555555556 0.181818181818 0 1.6 1e-06 
0.611111111111 0.181818181818 0 1.6 1e-06 
0.666666666667 0.181818181818 0 1.6 1e-06 
0.722222222222 0.181818181818 0 1.6 1e-06 
0.777777777778 0.181818181818 0 1.6 1e-06 
0.833333333333 0.181818181818 0 1.6 1e-06 
0.888888888889 0.181818181818 0 1.6 1e-06 
0.944444444444 0.181818181818 0 1.6 1e-06 
1.0 0.181818181818 0 1.6 1e-06 
0.5 0.222222222222 0 1.6 1e-06 
0.555555555556 0.222222222222 0 1.6 1e-06 
0.611111111111 0.222222222222 0 1.6 1e-06 
0.666666666667 0.222222222222 0 1.6 1e-06 
0.722222222222 0.222222222222 0 1.6 1e-06 
0.777777777778 0.222222222222 0 1.6 1e-06 
0.833333333333 0.222222222222 0 1.6 1e-06 
0.888888888889 0.222222222222 0 1.6 1e-06 
0.944444444444 0.222222222222 0 1.6 1e-06 
1.0 0.222222222222 0 1.6 1e-06 
0.5 0.262626262626 0 1.6 1e-06 
0.555555555556 0.262626262626 0 1.6 1e-06 
0.611111111111 0.262626262626 0 1.6 1e-06 
0.666666666667 0.262626262626 0 1.6 1e-06 
0.722222222222 0.262626262626 0 1.6 1e-06 
0.777777777778 0.262626262626 0 1.6 1e-06 
0.833333333333 0.262626262626 0 1.6 1e-06 
0.888888888889 0.262626262626 0 1.6 1e-06 
0.944444444444 0.262626262626 0 1.6 1e-06 
1.0 0.262626262626 0 1.6 1e-06 
0.5 0.30303030303 0 1.6 1e-06 
0.555555555556 0.30303030303 0 1.6 1e-06 
0.611111111111 0.30303030303 0 1.6 1e-06 
0.666666666667 0.30303030303 0 1.6 1e-06 
0.722222222222 0.30303030303 0 1.6 1e-06 
0.777777777778 0.30303030303 0 1.6 1e-06 
0.833333333333 0.30303030303 0 1.6 1e-06 
0.888888888889 0.30303030303 0 1.6 1e-06 
0.944444444444 0.30303030303 0 1.6 1e-06 
1.0 0.30303030303 0 1.6 1e-06 
0.5 0.343434343434 0 1.6 1e-06 
0.555555555556 0.343434343434 0 1.6 1e-06 
0.611111111111 0.343434343434 0 1.6 1e-06 
0.666666666667 0.343434343434 0 1.6 1e-06 
0.722222222222 0.343434343434 0 1.6 1e-06 
0.777777777778 0.343434343434 0 1.6 1e-06 
0.833333333333 0.343434343434 0 1.6 1e-06 
0.888888888889 0.343434343434 0 1.6 1e-06 
0.944444444444 0.343434343434 0 1.6 1e-06 
1.0 0.343434343434 0 1.6 1e-06 
0.5 0.383838383838 0 1.6 1e-06 
0.555555555556 0.383838383838 0 1.6 1e-06 
0.611111111111 0.383838383838 0 1.6 1e-06 
0.666666666667 0.383838383838 0 1.6 1e-06 
0.722222222222 0.383838383838 0 1.6 1e-06 
0.777777777778 0.383838383838 0 1.6 1e-06 
0.833333333333 0.383838383838 0 1.6 1e-06 
0.888888888889 0.383838383838 0 1.6 1e-06 
0.944444444444 0.383838383838 0 1.6 1e-06 
1.0 0.383838383838 0 1.6 1e-06 
0.5 0.424242424242 0 1.6 1e-06 
0.555555555556 0.424242424242 0 1.6 1e-06 
0.611111111111 0.424242424242 0 1.6 1e-06 
0.666666666667 0.424242424242 0 1.6 1e-06 
0.722222222222 0.424242424242 0 1.6 1e-06 
0.777777777778 0.424242424242 0 1.6 1e-06 
0.833333333333 0.424242424242 0 1.6 1e-06 
0.888888888889 0.424242424242 0 1.6 1e-06 
0.944444444444 0.424242424242 0 1.6 1e-06 
1.0 0.424242424242 0 1.6 1e-06 
0.5 0.464646464646 0 1.6 1e-06 
0.555555555556 0.464646464646 0 1.6 1e-06 
0.611111111111 0.464646464646 0 1.6 1e-06 
0.666666666667 0.464646464646 0 1.6 1e-06 
0.722222222222 0.464646464646 0 1.6 1e-06 
0.777777777778 0.464646464646 0 1.6 1e-06 
0.833333333333 0.464646464646 0 1.6 1e-06 
0.888888888889 0.464646464646 0 1.6 1e-06 
0.944444444444 0.464646464646 0 1.6 1e-06 
1.0 0.464646464646 0 1.6 1e-06 
0.5 0.505050505051 0 1.6 1e-06 
0.555555555556 0.505050505051 0 1.6 1e-06 
0.611111111111 0.505050505051 0 1.6 1e-06 
0.666666666667 0.505050505051 0 1.6 1e-06 
0.722222222222 0.505050505051 0 1.6 1e-06 
0.777777777778 0.505050505051 0 1.6 1e-06 
0.833333333333 0.505050505051 0 1.6 1e-06 
0.888888888889 0.505050505051 0 1.6 1e-06 
0.944444444444 0.505050505051 0 1.6 1e-06 
1.0 0.505050505051 0 1.6 1e-06 
0.5 0.545454545455 0 1.6 1e-06 
0.555555555556 0.545454545455 0 1.6 1e-06 
0.611111111111 0.545454545455 0 1.6 1e-06 
0.666666666667 0.545454545455 0 1.6 1e-06 
0.722222222222 0.545454545455 0 1.6 1e-06 
0.777777777778 0.545454545455 0 1.6 1e-06 
0.833333333333 0.545454545455 0 1.6 1e-06 
0.888888888889 0.545454545455 0 1.6 1e-06 
0.944444444444 0.545454545455 0 1.6 1e-06 
1.0 0.545454545455 0 1.6 1e-06 
0.5 0.585858585859 0 1.6 1e-06 
0.555555555556 0.585858585859 0 1.6 1e-06 
0.611111111111 0.585858585859 0 1.6 1e-06 
0.666666666667 0.585858585859 0 1.6 1e-06 
0.722222222222 0.585858585859 0 1.6 1e-06 
0.777777777778 0.585858585859 0 1.6 1e-06 
0.833333333333 0.585858585859 0 1.6 1e-06 
0.888888888889 0.585858585859 0 1.6 1e-06 
0.944444444444 0.585858585859 0 1.6 1e-06 
1.0 0.585858585859 0 1.6 1e-06 
0.5 0.626262626263 0 1.6 1e-06 
0.555555555556 0.626262626263 0 1.6 1e-06 
0.611111111111 0.626262626263 0 1.6 1e-06 
0.666666666667 0.626262626263 0 1.6 1e-06 
0.722222222222 0.626262626263 0 1.6 1e-06 
0.777777777778 0.626262626263 0 1.6 1e-06 
0.833333333333 0.626262626263 0 1.6 1e-06 
0.888888888889 0.626262626263 0 1.6 1e-06 
0.944444444444 0.626262626263 0 1.6 1e-06 
1.0 0.626262626263 0 1.6 1e-06 
0.5 0.666666666667 0 1.6 1e-06 
0.555555555556 0.666666666667 0 1.6 1e-06 
0.611111111111 0.666666666667 0 1.6 1e-06 
0.666666666667 0.666666666667 0 1.6 1e-06 
0.722222222222 0.666666666667 0 1.6 1e-06 
0.777777777778 0.666666666667 0 1.6 1e-06 
0.833333333333 0.666666666667 0 1.6 1e-06 
0.888888888889 0.666666666667 0 1.6 1e-06 
0.944444444444 0.666666666667 0 1.6 1e-06 
1.0 0.666666666667 0 1.6 1e-06 
0.5 0.707070707071 0 1.6 1e-06 
0.555555555556 0.707070707071 0 1.6 1e-06 
0.611111111111 0.707070707071 0 1.6 1e-06 
0.666666666667 0.707070707071 0 1.6 1e-06 
0.722222222222 0.707070707071 0 1.6 1e-06 
0.777777777778 0.707070707071 0 1.6 1e-06 
0.833333333333 0.707070707071 0 1.6 1e-06 
0.888888888889 0.707070707071 0 1.6 1e-06 
0.944444444444 0.707070707071 0 1.6 1e-06 
1.0 0.707070707071 0 1.6 1e-06 
0.5 0.747474747475 0 1.6 1e-06 
0.555555555556 0.747474747475 0 1.6 1e-06 
0.611111111111 0.747474747475 0 1.6 1e-06 
0.666666666667 0.747474747475 0 1.6 1e-06 
0.722222222222 0.747474747475 0 1.6 1e-06 
0.777777777778 0.747474747475 0 1.6 1e-06 
0.833333333333 0.747474747475 0 1.6 1e-06 
0.888888888889 0.747474747475 0 1.6 1e-06 
0.944444444444 0.747474747475 0 1.6 1e-06 
1.0 0.747474747475 0 1.6 1e-06 
0.5 0.787878787879 0 1.6 1e-06 
0.555555555556 0.787878787879 0 1.6 1e-06 
0.611111111111 0.787878787879 0 1.6 1e-06 
0.666666666667 0.787878787879 0 1.6 1e-06 
0.722222222222 0.787878787879 0 1.6 1e-06 
0.777777777778 0.787878787879 0 1.6 1e-06 
0.833333333333 0.787878787879 0 1.6 1e-06 
0.888888888889 0.787878787879 0 1.6 1e-06 
0.944444444444 0.787878787879 0 1.6 1e-06 
1.0 0.787878787879 0 1.6 1e-06 
0.5 0.828282828283 0 1.6 1e-06 
0.555555555556 0.828282828283 0 1.6 1e-06 
0.611111111111 0.828282828283 0 1.6 1e-06 
0.666666666667 0.828282828283 0 1.6 1e-06 
0.722222222222 0.828282828283 0 1.6 1e-06 
0.777777777778 0.828282828283 0 1.6 1e-06 
0.833333333333 0.828282828283 0 1.6 1e-06 
0.888888888889 0.828282828283 0 1.6 1e-06 
0.944444444444 0.828282828283 0 1.6 1e-06 
1.0 0.828282828283 0 1.6 1e-06 
0.5 0.868686868687 0 1.6 1e-06 
0.555555555556 0.868686868687 0 1.6 1e-06 
0.611111111111 0.868686868687 0 1.6 1e-06 
0.666666666667 0.868686868687 0 1.6 1e-06 
0.722222222222 0.868686868687 0 1.6 1e-06 
0.777777777778 0.868686868687 0 1.6 1e-06 
0.833333333333 0.868686868687 0 1.6 1e-06 
0.888888888889 0.868686868687 0 1.6 1e-06 
0.944444444444 0.868686868687 0 1.6 1e-06 
1.0 0.868686868687 0 1.6 1e-06 
0.5 0.909090909091 0 1.6 1e-06 
0.555555555556 0.909090909091 0 1.6 1e-06 
0.611111111111 0.909090909091 0 1.6 1e-06 
0.666666666667 0.909090909091 0 1.6 1e-06 
0.722222222222 0.909090909091 0 1.6 1e-06 
0.777777777778 0.909090909091 0 1.6 1e-06 
0.833333333333 0.909090909091 0 1.6 1e-06 
0.888888888889 0.909090909091 0 1.6 1e-06 
0.944444444444 0.909090909091 0 1.6 1e-06 
1.0 0.909090909091 0 1.6 1e-06 
0.5 0.949494949495 0 1.6 1e-06 
0.555555555556 0.949494949495 0 1.6 1e-06 
0.611111111111 0.949494949495 0 1.6 1e-06 
0.666666666667 0.949494949495 0 1.6 1e-06 
0.722222222222 0.949494949495 0 1.6 1e-06 
0.777777777778 0.949494949495 0 1.6 1e-06 
0.833333333333 0.949494949495 0 1.6 1e-06 
0.888888888889 0.949494949495 0 1.6 1e-06 
0.944444444444 0.949494949495 0 1.6 1e-06 
1.0 0.949494949495 0 1.6 1e-06 
0.5 0.989898989899 0 1.6 1e-06 
0.555555555556 0.989898989899 0 1.6 1e-06 
0.611111111111 0.989898989899 0 1.6 1e-06 
0.666666666667 0.989898989899 0 1.6 1e-06 
0.722222222222 0.989898989899 0 1.6 1e-06 
0.777777777778 0.989898989899 0 1.6 1e-06 
0.833333333333 0.989898989899 0 1.6 1e-06 
0.888888888889 0.989898989899 0 1.6 1e-06 
0.944444444444 0.989898989899 0 1.6 1e-06 
1.0 0.989898989899 0 1.6 1e-06 
0.5 1.0303030303 0 1.6 1e-06 
0.555555555556 1.0303030303 0 1.6 1e-06 
0.611111111111 1.0303030303 0 1.6 1e-06 
0.666666666667 1.0303030303 0 1.6 1e-06 
0.722222222222 1.0303030303 0 1.6 1e-06 
0.777777777778 1.0303030303 0 1.6 1e-06 
0.833333333333 1.0303030303 0 1.6 1e-06 
0.888888888889 1.0303030303 0 1.6 1e-06 
0.944444444444 1.0303030303 0 1.6 1e-06 
1.0 1.0303030303 0 1.6 1e-06 
0.5 1.07070707071 0 1.6 1e-06 
0.555555555556 1.07070707071 0 1.6 1e-06 
0.611111111111 1.07070707071 0 1.6 1e-06 
0.666666666667 1.07070707071 0 1.6 1e-06 
0.722222222222 1.07070707071 0 1.6 1e-06 
0.777777777778 1.07070707071 0 1.6 1e-06 
0.833333333333 1.07070707071 0 1.6 1e-06 
0.888888888889 1.07070707071 0 1.6 1e-06 
0.944444444444 1.07070707071 0 1.6 1e-06 
1.0 1.07070707071 0 1.6 1e-06 
0.5 1.11111111111 0 1.6 1e-06 
0.555555555556 1.11111111111 0 1.6 1e-06 
0.611111111111 1.11111111111 0 1.6 1e-06 
0.666666666667 1.11111111111 0 1.6 1e-06 
0.722222222222 1.11111111111 0 1.6 1e-06 
0.777777777778 1.11111111111 0 1.6 1e-06 
0.833333333333 1.11111111111 0 1.6 1e-06 
0.888888888889 1.11111111111 0 1.6 1e-06 
0.944444444444 1.11111111111 0 1.6 1e-06 
1.0 1.11111111111 0 1.6 1e-06 
0.5 1.15151515152 0 1.6 1e-06 
0.555555555556 1.15151515152 0 1.6 1e-06 
0.611111111111 1.15151515152 0 1.6 1e-06 
0.666666666667 1.15151515152 0 1.6 1e-06 
0.722222222222 1.15151515152 0 1.6 1e-06 
0.777777777778 1.15151515152 0 1.6 1e-06 
0.833333333333 1.15151515152 0 1.6 1e-06 
0.888888888889 1.15151515152 0 1.6 1e-06 
0.944444444444 1.15151515152 0 1.6 1e-06 
1.0 1.15151515152 0 1.6 1e-06 
0.5 1.19191919192 0 1.6 1e-06 
0.555555555556 1.19191919192 0 1.6 1e-06 
0.611111111111 1.19191919192 0 1.6 1e-06 
0.666666666667 1.19191919192 0 1.6 1e-06 
0.722222222222 1.19191919192 0 1.6 1e-06 
0.777777777778 1.19191919192 0 1.6 1e-06 
0.833333333333 1.19191919192 0 1.6 1e-06 
0.888888888889 1.19191919192 0 1.6 1e-06 
0.944444444444 1.19191919192 0 1.6 1e-06 
1.0 1.19191919192 0 1.6 1e-06 
0.5 1.23232323232 0 1.6 1e-06 
0.555555555556 1.23232323232 0 1.6 1e-06 
0.611111111111 1.23232323232 0 1.6 1e-06 
0.666666666667 1.23232323232 0 1.6 1e-06 
0.722222222222 1.23232323232 0 1.6 1e-06 
0.777777777778 1.23232323232 0 1.6 1e-06 
0.833333333333 1.23232323232 0 1.6 1e-06 
0.888888888889 1.23232323232 0 1.6 1e-06 
0.944444444444 1.23232323232 0 1.6 1e-06 
1.0 1.23232323232 0 1.6 1e-06 
0.5 1.27272727273 0 1.6 1e-06 
0.555555555556 1.27272727273 0 1.6 1e-06 
0.611111111111 1.27272727273 0 1.6 1e-06 
0.666666666667 1.27272727273 0 1.6 1e-06 
0.722222222222 1.27272727273 0 1.6 1e-06 
0.777777777778 1.27272727273 0 1.6 1e-06 
0.833333333333 1.27272727273 0 1.6 1e-06 
0.888888888889 1.27272727273 0 1.6 1e-06 
0.944444444444 1.27272727273 0 1.6 1e-06 
1.0 1.27272727273 0 1.6 1e-06 
0.5 1.31313131313 0 1.6 1e-06 
0.555555555556 1.31313131313 0 1.6 1e-06 
0.611111111111 1.31313131313 0 1.6 1e-06 
0.666666666667 1.31313131313 0 1.6 1e-06 
0.722222222222 1.31313131313 0 1.6 1e-06 
0.777777777778 1.31313131313 0 1.6 1e-06 
0.833333333333 1.31313131313 0 1.6 1e-06 
0.888888888889 1.31313131313 0 1.6 1e-06 
0.944444444444 1.31313131313 0 1.6 1e-06 
1.0 1.31313131313 0 1.6 1e-06 
0.5 1.35353535354 0 1.6 1e-06 
0.555555555556 1.35353535354 0 1.6 1e-06 
0.611111111111 1.35353535354 0 1.6 1e-06 
0.666666666667 1.35353535354 0 1.6 1e-06 
0.722222222222 1.35353535354 0 1.6 1e-06 
0.777777777778 1.35353535354 0 1.6 1e-06 
0.833333333333 1.35353535354 0 1.6 1e-06 
0.888888888889 1.35353535354 0 1.6 1e-06 
0.944444444444 1.35353535354 0 1.6 1e-06 
1.0 1.35353535354 0 1.6 1e-06 
0.5 1.39393939394 0 1.6 1e-06 
0.555555555556 1.39393939394 0 1.6 1e-06 
0.611111111111 1.39393939394 0 1.6 1e-06 
0.666666666667 1.39393939394 0 1.6 1e-06 
0.722222222222 1.39393939394 0 1.6 1e-06 
0.777777777778 1.39393939394 0 1.6 1e-06 
0.833333333333 1.39393939394 0 1.6 1e-06 
0.888888888889 1.39393939394 0 1.6 1e-06 
0.944444444444 1.39393939394 0 1.6 1e-06 
1.0 1.39393939394 0 1.6 1e-06 
0.5 1.43434343434 0 1.6 1e-06 
0.555555555556 1.43434343434 0 1.6 1e-06 
0.611111111111 1.43434343434 0 1.6 1e-06 
0.666666666667 1.43434343434 0 1.6 1e-06 
0.722222222222 1.43434343434 0 1.6 1e-06 
0.777777777778 1.43434343434 0 1.6 1e-06 
0.833333333333 1.43434343434 0 1.6 1e-06 
0.888888888889 1.43434343434 0 1.6 1e-06 
0.944444444444 1.43434343434 0 1.6 1e-06 
1.0 1.43434343434 0 1.6 1e-06 
0.5 1.47474747475 0 1.6 1e-06 
0.555555555556 1.47474747475 0 1.6 1e-06 
0.611111111111 1.47474747475 0 1.6 1e-06 
0.666666666667 1.47474747475 0 1.6 1e-06 
0.722222222222 1.47474747475 0 1.6 1e-06 
0.777777777778 1.47474747475 0 1.6 1e-06 
0.833333333333 1.47474747475 0 1.6 1e-06 
0.888888888889 1.47474747475 0 1.6 1e-06 
0.944444444444 1.47474747475 0 1.6 1e-06 
1.0 1.47474747475 0 1.6 1e-06 
0.5 1.51515151515 0 1.6 1e-06 
0.555555555556 1.51515151515 0 1.6 1e-06 
0.611111111111 1.51515151515 0 1.6 1e-06 
0.666666666667 1.51515151515 0 1.6 1e-06 
0.722222222222 1.51515151515 0 1.6 1e-06 
0.777777777778 1.51515151515 0 1.6 1e-06 
0.833333333333 1.51515151515 0 1.6 1e-06 
0.888888888889 1.51515151515 0 1.6 1e-06 
0.944444444444 1.51515151515 0 1.6 1e-06 
1.0 1.51515151515 0 1.6 1e-06 
0.5 1.55555555556 0 1.6 1e-06 
0.555555555556 1.55555555556 0 1.6 1e-06 
0.611111111111 1.55555555556 0 1.6 1e-06 
0.666666666667 1.55555555556 0 1.6 1e-06 
0.722222222222 1.55555555556 0 1.6 1e-06 
0.777777777778 1.55555555556 0 1.6 1e-06 
0.833333333333 1.55555555556 0 1.6 1e-06 
0.888888888889 1.55555555556 0 1.6 1e-06 
0.944444444444 1.55555555556 0 1.6 1e-06 
1.0 1.55555555556 0 1.6 1e-06 
0.5 1.59595959596 0 1.6 1e-06 
0.555555555556 1.59595959596 0 1.6 1e-06 
0.611111111111 1.59595959596 0 1.6 1e-06 
0.666666666667 1.59595959596 0 1.6 1e-06 
0.722222222222 1.59595959596 0 1.6 1e-06 
0.777777777778 1.59595959596 0 1.6 1e-06 
0.833333333333 1.59595959596 0 1.6 1e-06 
0.888888888889 1.59595959596 0 1.6 1e-06 
0.944444444444 1.59595959596 0 1.6 1e-06 
1.0 1.59595959596 0 1.6 1e-06 
0.5 1.63636363636 0 1.6 1e-06 
0.555555555556 1.63636363636 0 1.6 1e-06 
0.611111111111 1.63636363636 0 1.6 1e-06 
0.666666666667 1.63636363636 0 1.6 1e-06 
0.722222222222 1.63636363636 0 1.6 1e-06 
0.777777777778 1.63636363636 0 1.6 1e-06 
0.833333333333 1.63636363636 0 1.6 1e-06 
0.888888888889 1.63636363636 0 1.6 1e-06 
0.944444444444 1.63636363636 0 1.6 1e-06 
1.0 1.63636363636 0 1.6 1e-06 
0.5 1.67676767677 0 1.6 1e-06 
0.555555555556 1.67676767677 0 1.6 1e-06 
0.611111111111 1.67676767677 0 1.6 1e-06 
0.666666666667 1.67676767677 0 1.6 1e-06 
0.722222222222 1.67676767677 0 1.6 1e-06 
0.777777777778 1.67676767677 0 1.6 1e-06 
0.833333333333 1.67676767677 0 1.6 1e-06 
0.888888888889 1.67676767677 0 1.6 1e-06 
0.944444444444 1.67676767677 0 1.6 1e-06 
1.0 1.67676767677 0 1.6 1e-06 
0.5 1.71717171717 0 1.6 1e-06 
0.555555555556 1.71717171717 0 1.6 1e-06 
0.611111111111 1.71717171717 0 1.6 1e-06 
0.666666666667 1.71717171717 0 1.6 1e-06 
0.722222222222 1.71717171717 0 1.6 1e-06 
0.777777777778 1.71717171717 0 1.6 1e-06 
0.833333333333 1.71717171717 0 1.6 1e-06 
0.888888888889 1.71717171717 0 1.6 1e-06 
0.944444444444 1.71717171717 0 1.6 1e-06 
1.0 1.71717171717 0 1.6 1e-06 
0.5 1.75757575758 0 1.6 1e-06 
0.555555555556 1.75757575758 0 1.6 1e-06 
0.611111111111 1.75757575758 0 1.6 1e-06 
0.666666666667 1.75757575758 0 1.6 1e-06 
0.722222222222 1.75757575758 0 1.6 1e-06 
0.777777777778 1.75757575758 0 1.6 1e-06 
0.833333333333 1.75757575758 0 1.6 1e-06 
0.888888888889 1.75757575758 0 1.6 1e-06 
0.944444444444 1.75757575758 0 1.6 1e-06 
1.0 1.75757575758 0 1.6 1e-06 
0.5 1.79797979798 0 1.6 1e-06 
0.555555555556 1.79797979798 0 1.6 1e-06 
0.611111111111 1.79797979798 0 1.6 1e-06 
0.666666666667 1.79797979798 0 1.6 1e-06 
0.722222222222 1.79797979798 0 1.6 1e-06 
0.777777777778 1.79797979798 0 1.6 1e-06 
0.833333333333 1.79797979798 0 1.6 1e-06 
0.888888888889 1.79797979798 0 1.6 1e-06 
0.944444444444 1.79797979798 0 1.6 1e-06 
1.0 1.79797979798 0 1.6 1e-06 
0.5 1.83838383838 0 1.6 1e-06 
0.555555555556 1.83838383838 0 1.6 1e-06 
0.611111111111 1.83838383838 0 1.6 1e-06 
0.666666666667 1.83838383838 0 1.6 1e-06 
0.722222222222 1.83838383838 0 1.6 1e-06 
0.777777777778 1.83838383838 0 1.6 1e-06 
0.833333333333 1.83838383838 0 1.6 1e-06 
0.888888888889 1.83838383838 0 1.6 1e-06 
0.944444444444 1.83838383838 0 1.6 1e-06 
1.0 1.83838383838 0 1.6 1e-06 
0.5 1.87878787879 0 1.6 1e-06 
0.555555555556 1.87878787879 0 1.6 1e-06 
0.611111111111 1.87878787879 0 1.6 1e-06 
0.666666666667 1.87878787879 0 1.6 1e-06 
0.722222222222 1.87878787879 0 1.6 1e-06 
0.777777777778 1.87878787879 0 1.6 1e-06 
0.833333333333 1.87878787879 0 1.6 1e-06 
0.888888888889 1.87878787879 0 1.6 1e-06 
0.944444444444 1.87878787879 0 1.6 1e-06 
1.0 1.87878787879 0 1.6 1e-06 
0.5 1.91919191919 0 1.6 1e-06 
0.555555555556 1.91919191919 0 1.6 1e-06 
0.611111111111 1.91919191919 0 1.6 1e-06 
0.666666666667 1.91919191919 0 1.6 1e-06 
0.722222222222 1.91919191919 0 1.6 1e-06 
0.777777777778 1.91919191919 0 1.6 1e-06 
0.833333333333 1.91919191919 0 1.6 1e-06 
0.888888888889 1.91919191919 0 1.6 1e-06 
0.944444444444 1.91919191919 0 1.6 1e-06 
1.0 1.91919191919 0 1.6 1e-06 
0.5 1.9595959596 0 1.6 1e-06 
0.555555555556 1.9595959596 0 1.6 1e-06 
0.611111111111 1.9595959596 0 1.6 1e-06 
0.666666666667 1.9595959596 0 1.6 1e-06 
0.722222222222 1.9595959596 0 1.6 1e-06 
0.777777777778 1.9595959596 0 1.6 1e-06 
0.833333333333 1.9595959596 0 1.6 1e-06 
0.888888888889 1.9595959596 0 1.6 1e-06 
0.944444444444 1.9595959596 0 1.6 1e-06 
1.0 1.9595959596 0 1.6 1e-06 
0.5 2.0 0 1.6 1e-06 
0.555555555556 2.0 0 1.6 1e-06 
0.611111111111 2.0 0 1.6 1e-06 
0.666666666667 2.0 0 1.6 1e-06 
0.722222222222 2.0 0 1.6 1e-06 
0.777777777778 2.0 0 1.6 1e-06 
0.833333333333 2.0 0 1.6 1e-06 
0.888888888889 2.0 0 1.6 1e-06 
0.944444444444 2.0 0 1.6 1e-06 
1.0 2.0 0 1.6 1e-06 
0.5 -2.0 0 2.0 1e-06 
0.555555555556 -2.0 0 2.0 1e-06 
0.611111111111 -2.0 0 2.0 1e-06 
0.666666666667 -2.0 0 2.0 1e-06 
0.722222222222 -2.0 0 2.0 1e-06 
0.777777777778 -2.0 0 2.0 1e-06 
0.833333333333 -2.0 0 2.0 1e-06 
0.888888888889 -2.0 0 2.0 1e-06 
0.944444444444 -2.0 0 2.0 1e-06 
1.0 -2.0 0 2.0 1e-06 
0.5 -1.9595959596 0 2.0 1e-06 
0.555555555556 -1.9595959596 0 2.0 1e-06 
0.611111111111 -1.9595959596 0 2.0 1e-06 
0.666666666667 -1.9595959596 0 2.0 1e-06 
0.722222222222 -1.9595959596 0 2.0 1e-06 
0.777777777778 -1.9595959596 0 2.0 1e-06 
0.833333333333 -1.9595959596 0 2.0 1e-06 
0.888888888889 -1.9595959596 0 2.0 1e-06 
0.944444444444 -1.9595959596 0 2.0 1e-06 
1.0 -1.9595959596 0 2.0 1e-06 
0.5 -1.91919191919 0 2.0 1e-06 
0.555555555556 -1.91919191919 0 2.0 1e-06 
0.611111111111 -1.91919191919 0 2.0 1e-06 
0.666666666667 -1.91919191919 0 2.0 1e-06 
0.722222222222 -1.91919191919 0 2.0 1e-06 
0.777777777778 -1.91919191919 0 2.0 1e-06 
0.833333333333 -1.91919191919 0 2.0 1e-06 
0.888888888889 -1.91919191919 0 2.0 1e-06 
0.944444444444 -1.91919191919 0 2.0 1e-06 
1.0 -1.91919191919 0 2.0 1e-06 
0.5 -1.87878787879 0 2.0 1e-06 
0.555555555556 -1.87878787879 0 2.0 1e-06 
0.611111111111 -1.87878787879 0 2.0 1e-06 
0.666666666667 -1.87878787879 0 2.0 1e-06 
0.722222222222 -1.87878787879 0 2.0 1e-06 
0.777777777778 -1.87878787879 0 2.0 1e-06 
0.833333333333 -1.87878787879 0 2.0 1e-06 
0.888888888889 -1.87878787879 0 2.0 1e-06 
0.944444444444 -1.87878787879 0 2.0 1e-06 
1.0 -1.87878787879 0 2.0 1e-06 
0.5 -1.83838383838 0 2.0 1e-06 
0.555555555556 -1.83838383838 0 2.0 1e-06 
0.611111111111 -1.83838383838 0 2.0 1e-06 
0.666666666667 -1.83838383838 0 2.0 1e-06 
0.722222222222 -1.83838383838 0 2.0 1e-06 
0.777777777778 -1.83838383838 0 2.0 1e-06 
0.833333333333 -1.83838383838 0 2.0 1e-06 
0.888888888889 -1.83838383838 0 2.0 1e-06 
0.944444444444 -1.83838383838 0 2.0 1e-06 
1.0 -1.83838383838 0 2.0 1e-06 
0.5 -1.79797979798 0 2.0 1e-06 
0.555555555556 -1.79797979798 0 2.0 1e-06 
0.611111111111 -1.79797979798 0 2.0 1e-06 
0.666666666667 -1.79797979798 0 2.0 1e-06 
0.722222222222 -1.79797979798 0 2.0 1e-06 
0.777777777778 -1.79797979798 0 2.0 1e-06 
0.833333333333 -1.79797979798 0 2.0 1e-06 
0.888888888889 -1.79797979798 0 2.0 1e-06 
0.944444444444 -1.79797979798 0 2.0 1e-06 
1.0 -1.79797979798 0 2.0 1e-06 
0.5 -1.75757575758 0 2.0 1e-06 
0.555555555556 -1.75757575758 0 2.0 1e-06 
0.611111111111 -1.75757575758 0 2.0 1e-06 
0.666666666667 -1.75757575758 0 2.0 1e-06 
0.722222222222 -1.75757575758 0 2.0 1e-06 
0.777777777778 -1.75757575758 0 2.0 1e-06 
0.833333333333 -1.75757575758 0 2.0 1e-06 
0.888888888889 -1.75757575758 0 2.0 1e-06 
0.944444444444 -1.75757575758 0 2.0 1e-06 
1.0 -1.75757575758 0 2.0 1e-06 
0.5 -1.71717171717 0 2.0 1e-06 
0.555555555556 -1.71717171717 0 2.0 1e-06 
0.611111111111 -1.71717171717 0 2.0 1e-06 
0.666666666667 -1.71717171717 0 2.0 1e-06 
0.722222222222 -1.71717171717 0 2.0 1e-06 
0.777777777778 -1.71717171717 0 2.0 1e-06 
0.833333333333 -1.71717171717 0 2.0 1e-06 
0.888888888889 -1.71717171717 0 2.0 1e-06 
0.944444444444 -1.71717171717 0 2.0 1e-06 
1.0 -1.71717171717 0 2.0 1e-06 
0.5 -1.67676767677 0 2.0 1e-06 
0.555555555556 -1.67676767677 0 2.0 1e-06 
0.611111111111 -1.67676767677 0 2.0 1e-06 
0.666666666667 -1.67676767677 0 2.0 1e-06 
0.722222222222 -1.67676767677 0 2.0 1e-06 
0.777777777778 -1.67676767677 0 2.0 1e-06 
0.833333333333 -1.67676767677 0 2.0 1e-06 
0.888888888889 -1.67676767677 0 2.0 1e-06 
0.944444444444 -1.67676767677 0 2.0 1e-06 
1.0 -1.67676767677 0 2.0 1e-06 
0.5 -1.63636363636 0 2.0 1e-06 
0.555555555556 -1.63636363636 0 2.0 1e-06 
0.611111111111 -1.63636363636 0 2.0 1e-06 
0.666666666667 -1.63636363636 0 2.0 1e-06 
0.722222222222 -1.63636363636 0 2.0 1e-06 
0.777777777778 -1.63636363636 0 2.0 1e-06 
0.833333333333 -1.63636363636 0 2.0 1e-06 
0.888888888889 -1.63636363636 0 2.0 1e-06 
0.944444444444 -1.63636363636 0 2.0 1e-06 
1.0 -1.63636363636 0 2.0 1e-06 
0.5 -1.59595959596 0 2.0 1e-06 
0.555555555556 -1.59595959596 0 2.0 1e-06 
0.611111111111 -1.59595959596 0 2.0 1e-06 
0.666666666667 -1.59595959596 0 2.0 1e-06 
0.722222222222 -1.59595959596 0 2.0 1e-06 
0.777777777778 -1.59595959596 0 2.0 1e-06 
0.833333333333 -1.59595959596 0 2.0 1e-06 
0.888888888889 -1.59595959596 0 2.0 1e-06 
0.944444444444 -1.59595959596 0 2.0 1e-06 
1.0 -1.59595959596 0 2.0 1e-06 
0.5 -1.55555555556 0 2.0 1e-06 
0.555555555556 -1.55555555556 0 2.0 1e-06 
0.611111111111 -1.55555555556 0 2.0 1e-06 
0.666666666667 -1.55555555556 0 2.0 1e-06 
0.722222222222 -1.55555555556 0 2.0 1e-06 
0.777777777778 -1.55555555556 0 2.0 1e-06 
0.833333333333 -1.55555555556 0 2.0 1e-06 
0.888888888889 -1.55555555556 0 2.0 1e-06 
0.944444444444 -1.55555555556 0 2.0 1e-06 
1.0 -1.55555555556 0 2.0 1e-06 
0.5 -1.51515151515 0 2.0 1e-06 
0.555555555556 -1.51515151515 0 2.0 1e-06 
0.611111111111 -1.51515151515 0 2.0 1e-06 
0.666666666667 -1.51515151515 0 2.0 1e-06 
0.722222222222 -1.51515151515 0 2.0 1e-06 
0.777777777778 -1.51515151515 0 2.0 1e-06 
0.833333333333 -1.51515151515 0 2.0 1e-06 
0.888888888889 -1.51515151515 0 2.0 1e-06 
0.944444444444 -1.51515151515 0 2.0 1e-06 
1.0 -1.51515151515 0 2.0 1e-06 
0.5 -1.47474747475 0 2.0 1e-06 
0.555555555556 -1.47474747475 0 2.0 1e-06 
0.611111111111 -1.47474747475 0 2.0 1e-06 
0.666666666667 -1.47474747475 0 2.0 1e-06 
0.722222222222 -1.47474747475 0 2.0 1e-06 
0.777777777778 -1.47474747475 0 2.0 1e-06 
0.833333333333 -1.47474747475 0 2.0 1e-06 
0.888888888889 -1.47474747475 0 2.0 1e-06 
0.944444444444 -1.47474747475 0 2.0 1e-06 
1.0 -1.47474747475 0 2.0 1e-06 
0.5 -1.43434343434 0 2.0 1e-06 
0.555555555556 -1.43434343434 0 2.0 1e-06 
0.611111111111 -1.43434343434 0 2.0 1e-06 
0.666666666667 -1.43434343434 0 2.0 1e-06 
0.722222222222 -1.43434343434 0 2.0 1e-06 
0.777777777778 -1.43434343434 0 2.0 1e-06 
0.833333333333 -1.43434343434 0 2.0 1e-06 
0.888888888889 -1.43434343434 0 2.0 1e-06 
0.944444444444 -1.43434343434 0 2.0 1e-06 
1.0 -1.43434343434 0 2.0 1e-06 
0.5 -1.39393939394 0 2.0 1e-06 
0.555555555556 -1.39393939394 0 2.0 1e-06 
0.611111111111 -1.39393939394 0 2.0 1e-06 
0.666666666667 -1.39393939394 0 2.0 1e-06 
0.722222222222 -1.39393939394 0 2.0 1e-06 
0.777777777778 -1.39393939394 0 2.0 1e-06 
0.833333333333 -1.39393939394 0 2.0 1e-06 
0.888888888889 -1.39393939394 0 2.0 1e-06 
0.944444444444 -1.39393939394 0 2.0 1e-06 
1.0 -1.39393939394 0 2.0 1e-06 
0.5 -1.35353535354 0 2.0 1e-06 
0.555555555556 -1.35353535354 0 2.0 1e-06 
0.611111111111 -1.35353535354 0 2.0 1e-06 
0.666666666667 -1.35353535354 0 2.0 1e-06 
0.722222222222 -1.35353535354 0 2.0 1e-06 
0.777777777778 -1.35353535354 0 2.0 1e-06 
0.833333333333 -1.35353535354 0 2.0 1e-06 
0.888888888889 -1.35353535354 0 2.0 1e-06 
0.944444444444 -1.35353535354 0 2.0 1e-06 
1.0 -1.35353535354 0 2.0 1e-06 
0.5 -1.31313131313 0 2.0 1e-06 
0.555555555556 -1.31313131313 0 2.0 1e-06 
0.611111111111 -1.31313131313 0 2.0 1e-06 
0.666666666667 -1.31313131313 0 2.0 1e-06 
0.722222222222 -1.31313131313 0 2.0 1e-06 
0.777777777778 -1.31313131313 0 2.0 1e-06 
0.833333333333 -1.31313131313 0 2.0 1e-06 
0.888888888889 -1.31313131313 0 2.0 1e-06 
0.944444444444 -1.31313131313 0 2.0 1e-06 
1.0 -1.31313131313 0 2.0 1e-06 
0.5 -1.27272727273 0 2.0 1e-06 
0.555555555556 -1.27272727273 0 2.0 1e-06 
0.611111111111 -1.27272727273 0 2.0 1e-06 
0.666666666667 -1.27272727273 0 2.0 1e-06 
0.722222222222 -1.27272727273 0 2.0 1e-06 
0.777777777778 -1.27272727273 0 2.0 1e-06 
0.833333333333 -1.27272727273 0 2.0 1e-06 
0.888888888889 -1.27272727273 0 2.0 1e-06 
0.944444444444 -1.27272727273 0 2.0 1e-06 
1.0 -1.27272727273 0 2.0 1e-06 
0.5 -1.23232323232 0 2.0 1e-06 
0.555555555556 -1.23232323232 0 2.0 1e-06 
0.611111111111 -1.23232323232 0 2.0 1e-06 
0.666666666667 -1.23232323232 0 2.0 1e-06 
0.722222222222 -1.23232323232 0 2.0 1e-06 
0.777777777778 -1.23232323232 0 2.0 1e-06 
0.833333333333 -1.23232323232 0 2.0 1e-06 
0.888888888889 -1.23232323232 0 2.0 1e-06 
0.944444444444 -1.23232323232 0 2.0 1e-06 
1.0 -1.23232323232 0 2.0 1e-06 
0.5 -1.19191919192 0 2.0 1e-06 
0.555555555556 -1.19191919192 0 2.0 1e-06 
0.611111111111 -1.19191919192 0 2.0 1e-06 
0.666666666667 -1.19191919192 0 2.0 1e-06 
0.722222222222 -1.19191919192 0 2.0 1e-06 
0.777777777778 -1.19191919192 0 2.0 1e-06 
0.833333333333 -1.19191919192 0 2.0 1e-06 
0.888888888889 -1.19191919192 0 2.0 1e-06 
0.944444444444 -1.19191919192 0 2.0 1e-06 
1.0 -1.19191919192 0 2.0 1e-06 
0.5 -1.15151515152 0 2.0 1e-06 
0.555555555556 -1.15151515152 0 2.0 1e-06 
0.611111111111 -1.15151515152 0 2.0 1e-06 
0.666666666667 -1.15151515152 0 2.0 1e-06 
0.722222222222 -1.15151515152 0 2.0 1e-06 
0.777777777778 -1.15151515152 0 2.0 1e-06 
0.833333333333 -1.15151515152 0 2.0 1e-06 
0.888888888889 -1.15151515152 0 2.0 1e-06 
0.944444444444 -1.15151515152 0 2.0 1e-06 
1.0 -1.15151515152 0 2.0 1e-06 
0.5 -1.11111111111 0 2.0 1e-06 
0.555555555556 -1.11111111111 0 2.0 1e-06 
0.611111111111 -1.11111111111 0 2.0 1e-06 
0.666666666667 -1.11111111111 0 2.0 1e-06 
0.722222222222 -1.11111111111 0 2.0 1e-06 
0.777777777778 -1.11111111111 0 2.0 1e-06 
0.833333333333 -1.11111111111 0 2.0 1e-06 
0.888888888889 -1.11111111111 0 2.0 1e-06 
0.944444444444 -1.11111111111 0 2.0 1e-06 
1.0 -1.11111111111 0 2.0 1e-06 
0.5 -1.07070707071 0 2.0 1e-06 
0.555555555556 -1.07070707071 0 2.0 1e-06 
0.611111111111 -1.07070707071 0 2.0 1e-06 
0.666666666667 -1.07070707071 0 2.0 1e-06 
0.722222222222 -1.07070707071 0 2.0 1e-06 
0.777777777778 -1.07070707071 0 2.0 1e-06 
0.833333333333 -1.07070707071 0 2.0 1e-06 
0.888888888889 -1.07070707071 0 2.0 1e-06 
0.944444444444 -1.07070707071 0 2.0 1e-06 
1.0 -1.07070707071 0 2.0 1e-06 
0.5 -1.0303030303 0 2.0 1e-06 
0.555555555556 -1.0303030303 0 2.0 1e-06 
0.611111111111 -1.0303030303 0 2.0 1e-06 
0.666666666667 -1.0303030303 0 2.0 1e-06 
0.722222222222 -1.0303030303 0 2.0 1e-06 
0.777777777778 -1.0303030303 0 2.0 1e-06 
0.833333333333 -1.0303030303 0 2.0 1e-06 
0.888888888889 -1.0303030303 0 2.0 1e-06 
0.944444444444 -1.0303030303 0 2.0 1e-06 
1.0 -1.0303030303 0 2.0 1e-06 
0.5 -0.989898989899 0 2.0 1e-06 
0.555555555556 -0.989898989899 0 2.0 1e-06 
0.611111111111 -0.989898989899 0 2.0 1e-06 
0.666666666667 -0.989898989899 0 2.0 1e-06 
0.722222222222 -0.989898989899 0 2.0 1e-06 
0.777777777778 -0.989898989899 0 2.0 1e-06 
0.833333333333 -0.989898989899 0 2.0 1e-06 
0.888888888889 -0.989898989899 0 2.0 1e-06 
0.944444444444 -0.989898989899 0 2.0 1e-06 
1.0 -0.989898989899 0 2.0 1e-06 
0.5 -0.949494949495 0 2.0 1e-06 
0.555555555556 -0.949494949495 0 2.0 1e-06 
0.611111111111 -0.949494949495 0 2.0 1e-06 
0.666666666667 -0.949494949495 0 2.0 1e-06 
0.722222222222 -0.949494949495 0 2.0 1e-06 
0.777777777778 -0.949494949495 0 2.0 1e-06 
0.833333333333 -0.949494949495 0 2.0 1e-06 
0.888888888889 -0.949494949495 0 2.0 1e-06 
0.944444444444 -0.949494949495 0 2.0 1e-06 
1.0 -0.949494949495 0 2.0 1e-06 
0.5 -0.909090909091 0 2.0 1e-06 
0.555555555556 -0.909090909091 0 2.0 1e-06 
0.611111111111 -0.909090909091 0 2.0 1e-06 
0.666666666667 -0.909090909091 0 2.0 1e-06 
0.722222222222 -0.909090909091 0 2.0 1e-06 
0.777777777778 -0.909090909091 0 2.0 1e-06 
0.833333333333 -0.909090909091 0 2.0 1e-06 
0.888888888889 -0.909090909091 0 2.0 1e-06 
0.944444444444 -0.909090909091 0 2.0 1e-06 
1.0 -0.909090909091 0 2.0 1e-06 
0.5 -0.868686868687 0 2.0 1e-06 
0.555555555556 -0.868686868687 0 2.0 1e-06 
0.611111111111 -0.868686868687 0 2.0 1e-06 
0.666666666667 -0.868686868687 0 2.0 1e-06 
0.722222222222 -0.868686868687 0 2.0 1e-06 
0.777777777778 -0.868686868687 0 2.0 1e-06 
0.833333333333 -0.868686868687 0 2.0 1e-06 
0.888888888889 -0.868686868687 0 2.0 1e-06 
0.944444444444 -0.868686868687 0 2.0 1e-06 
1.0 -0.868686868687 0 2.0 1e-06 
0.5 -0.828282828283 0 2.0 1e-06 
0.555555555556 -0.828282828283 0 2.0 1e-06 
0.611111111111 -0.828282828283 0 2.0 1e-06 
0.666666666667 -0.828282828283 0 2.0 1e-06 
0.722222222222 -0.828282828283 0 2.0 1e-06 
0.777777777778 -0.828282828283 0 2.0 1e-06 
0.833333333333 -0.828282828283 0 2.0 1e-06 
0.888888888889 -0.828282828283 0 2.0 1e-06 
0.944444444444 -0.828282828283 0 2.0 1e-06 
1.0 -0.828282828283 0 2.0 1e-06 
0.5 -0.787878787879 0 2.0 1e-06 
0.555555555556 -0.787878787879 0 2.0 1e-06 
0.611111111111 -0.787878787879 0 2.0 1e-06 
0.666666666667 -0.787878787879 0 2.0 1e-06 
0.722222222222 -0.787878787879 0 2.0 1e-06 
0.777777777778 -0.787878787879 0 2.0 1e-06 
0.833333333333 -0.787878787879 0 2.0 1e-06 
0.888888888889 -0.787878787879 0 2.0 1e-06 
0.944444444444 -0.787878787879 0 2.0 1e-06 
1.0 -0.787878787879 0 2.0 1e-06 
0.5 -0.747474747475 0 2.0 1e-06 
0.555555555556 -0.747474747475 0 2.0 1e-06 
0.611111111111 -0.747474747475 0 2.0 1e-06 
0.666666666667 -0.747474747475 0 2.0 1e-06 
0.722222222222 -0.747474747475 0 2.0 1e-06 
0.777777777778 -0.747474747475 0 2.0 1e-06 
0.833333333333 -0.747474747475 0 2.0 1e-06 
0.888888888889 -0.747474747475 0 2.0 1e-06 
0.944444444444 -0.747474747475 0 2.0 1e-06 
1.0 -0.747474747475 0 2.0 1e-06 
0.5 -0.707070707071 0 2.0 1e-06 
0.555555555556 -0.707070707071 0 2.0 1e-06 
0.611111111111 -0.707070707071 0 2.0 1e-06 
0.666666666667 -0.707070707071 0 2.0 1e-06 
0.722222222222 -0.707070707071 0 2.0 1e-06 
0.777777777778 -0.707070707071 0 2.0 1e-06 
0.833333333333 -0.707070707071 0 2.0 1e-06 
0.888888888889 -0.707070707071 0 2.0 1e-06 
0.944444444444 -0.707070707071 0 2.0 1e-06 
1.0 -0.707070707071 0 2.0 1e-06 
0.5 -0.666666666667 0 2.0 1e-06 
0.555555555556 -0.666666666667 0 2.0 1e-06 
0.611111111111 -0.666666666667 0 2.0 1e-06 
0.666666666667 -0.666666666667 0 2.0 1e-06 
0.722222222222 -0.666666666667 0 2.0 1e-06 
0.777777777778 -0.666666666667 0 2.0 1e-06 
0.833333333333 -0.666666666667 0 2.0 1e-06 
0.888888888889 -0.666666666667 0 2.0 1e-06 
0.944444444444 -0.666666666667 0 2.0 1e-06 
1.0 -0.666666666667 0 2.0 1e-06 
0.5 -0.626262626263 0 2.0 1e-06 
0.555555555556 -0.626262626263 0 2.0 1e-06 
0.611111111111 -0.626262626263 0 2.0 1e-06 
0.666666666667 -0.626262626263 0 2.0 1e-06 
0.722222222222 -0.626262626263 0 2.0 1e-06 
0.777777777778 -0.626262626263 0 2.0 1e-06 
0.833333333333 -0.626262626263 0 2.0 1e-06 
0.888888888889 -0.626262626263 0 2.0 1e-06 
0.944444444444 -0.626262626263 0 2.0 1e-06 
1.0 -0.626262626263 0 2.0 1e-06 
0.5 -0.585858585859 0 2.0 1e-06 
0.555555555556 -0.585858585859 0 2.0 1e-06 
0.611111111111 -0.585858585859 0 2.0 1e-06 
0.666666666667 -0.585858585859 0 2.0 1e-06 
0.722222222222 -0.585858585859 0 2.0 1e-06 
0.777777777778 -0.585858585859 0 2.0 1e-06 
0.833333333333 -0.585858585859 0 2.0 1e-06 
0.888888888889 -0.585858585859 0 2.0 1e-06 
0.944444444444 -0.585858585859 0 2.0 1e-06 
1.0 -0.585858585859 0 2.0 1e-06 
0.5 -0.545454545455 0 2.0 1e-06 
0.555555555556 -0.545454545455 0 2.0 1e-06 
0.611111111111 -0.545454545455 0 2.0 1e-06 
0.666666666667 -0.545454545455 0 2.0 1e-06 
0.722222222222 -0.545454545455 0 2.0 1e-06 
0.777777777778 -0.545454545455 0 2.0 1e-06 
0.833333333333 -0.545454545455 0 2.0 1e-06 
0.888888888889 -0.545454545455 0 2.0 1e-06 
0.944444444444 -0.545454545455 0 2.0 1e-06 
1.0 -0.545454545455 0 2.0 1e-06 
0.5 -0.505050505051 0 2.0 1e-06 
0.555555555556 -0.505050505051 0 2.0 1e-06 
0.611111111111 -0.505050505051 0 2.0 1e-06 
0.666666666667 -0.505050505051 0 2.0 1e-06 
0.722222222222 -0.505050505051 0 2.0 1e-06 
0.777777777778 -0.505050505051 0 2.0 1e-06 
0.833333333333 -0.505050505051 0 2.0 1e-06 
0.888888888889 -0.505050505051 0 2.0 1e-06 
0.944444444444 -0.505050505051 0 2.0 1e-06 
1.0 -0.505050505051 0 2.0 1e-06 
0.5 -0.464646464646 0 2.0 1e-06 
0.555555555556 -0.464646464646 0 2.0 1e-06 
0.611111111111 -0.464646464646 0 2.0 1e-06 
0.666666666667 -0.464646464646 0 2.0 1e-06 
0.722222222222 -0.464646464646 0 2.0 1e-06 
0.777777777778 -0.464646464646 0 2.0 1e-06 
0.833333333333 -0.464646464646 0 2.0 1e-06 
0.888888888889 -0.464646464646 0 2.0 1e-06 
0.944444444444 -0.464646464646 0 2.0 1e-06 
1.0 -0.464646464646 0 2.0 1e-06 
0.5 -0.424242424242 0 2.0 1e-06 
0.555555555556 -0.424242424242 0 2.0 1e-06 
0.611111111111 -0.424242424242 0 2.0 1e-06 
0.666666666667 -0.424242424242 0 2.0 1e-06 
0.722222222222 -0.424242424242 0 2.0 1e-06 
0.777777777778 -0.424242424242 0 2.0 1e-06 
0.833333333333 -0.424242424242 0 2.0 1e-06 
0.888888888889 -0.424242424242 0 2.0 1e-06 
0.944444444444 -0.424242424242 0 2.0 1e-06 
1.0 -0.424242424242 0 2.0 1e-06 
0.5 -0.383838383838 0 2.0 1e-06 
0.555555555556 -0.383838383838 0 2.0 1e-06 
0.611111111111 -0.383838383838 0 2.0 1e-06 
0.666666666667 -0.383838383838 0 2.0 1e-06 
0.722222222222 -0.383838383838 0 2.0 1e-06 
0.777777777778 -0.383838383838 0 2.0 1e-06 
0.833333333333 -0.383838383838 0 2.0 1e-06 
0.888888888889 -0.383838383838 0 2.0 1e-06 
0.944444444444 -0.383838383838 0 2.0 1e-06 
1.0 -0.383838383838 0 2.0 1e-06 
0.5 -0.343434343434 0 2.0 1e-06 
0.555555555556 -0.343434343434 0 2.0 1e-06 
0.611111111111 -0.343434343434 0 2.0 1e-06 
0.666666666667 -0.343434343434 0 2.0 1e-06 
0.722222222222 -0.343434343434 0 2.0 1e-06 
0.777777777778 -0.343434343434 0 2.0 1e-06 
0.833333333333 -0.343434343434 0 2.0 1e-06 
0.888888888889 -0.343434343434 0 2.0 1e-06 
0.944444444444 -0.343434343434 0 2.0 1e-06 
1.0 -0.343434343434 0 2.0 1e-06 
0.5 -0.30303030303 0 2.0 1e-06 
0.555555555556 -0.30303030303 0 2.0 1e-06 
0.611111111111 -0.30303030303 0 2.0 1e-06 
0.666666666667 -0.30303030303 0 2.0 1e-06 
0.722222222222 -0.30303030303 0 2.0 1e-06 
0.777777777778 -0.30303030303 0 2.0 1e-06 
0.833333333333 -0.30303030303 0 2.0 1e-06 
0.888888888889 -0.30303030303 0 2.0 1e-06 
0.944444444444 -0.30303030303 0 2.0 1e-06 
1.0 -0.30303030303 0 2.0 1e-06 
0.5 -0.262626262626 0 2.0 1e-06 
0.555555555556 -0.262626262626 0 2.0 1e-06 
0.611111111111 -0.262626262626 0 2.0 1e-06 
0.666666666667 -0.262626262626 0 2.0 1e-06 
0.722222222222 -0.262626262626 0 2.0 1e-06 
0.777777777778 -0.262626262626 0 2.0 1e-06 
0.833333333333 -0.262626262626 0 2.0 1e-06 
0.888888888889 -0.262626262626 0 2.0 1e-06 
0.944444444444 -0.262626262626 0 2.0 1e-06 
1.0 -0.262626262626 0 2.0 1e-06 
0.5 -0.222222222222 0 2.0 1e-06 
0.555555555556 -0.222222222222 0 2.0 1e-06 
0.611111111111 -0.222222222222 0 2.0 1e-06 
0.666666666667 -0.222222222222 0 2.0 1e-06 
0.722222222222 -0.222222222222 0 2.0 1e-06 
0.777777777778 -0.222222222222 0 2.0 1e-06 
0.833333333333 -0.222222222222 0 2.0 1e-06 
0.888888888889 -0.222222222222 0 2.0 1e-06 
0.944444444444 -0.222222222222 0 2.0 1e-06 
1.0 -0.222222222222 0 2.0 1e-06 
0.5 -0.181818181818 0 2.0 1e-06 
0.555555555556 -0.181818181818 0 2.0 1e-06 
0.611111111111 -0.181818181818 0 2.0 1e-06 
0.666666666667 -0.181818181818 0 2.0 1e-06 
0.722222222222 -0.181818181818 0 2.0 1e-06 
0.777777777778 -0.181818181818 0 2.0 1e-06 
0.833333333333 -0.181818181818 0 2.0 1e-06 
0.888888888889 -0.181818181818 0 2.0 1e-06 
0.944444444444 -0.181818181818 0 2.0 1e-06 
1.0 -0.181818181818 0 2.0 1e-06 
0.5 -0.141414141414 0 2.0 1e-06 
0.555555555556 -0.141414141414 0 2.0 1e-06 
0.611111111111 -0.141414141414 0 2.0 1e-06 
0.666666666667 -0.141414141414 0 2.0 1e-06 
0.722222222222 -0.141414141414 0 2.0 1e-06 
0.777777777778 -0.141414141414 0 2.0 1e-06 
0.833333333333 -0.141414141414 0 2.0 1e-06 
0.888888888889 -0.141414141414 0 2.0 1e-06 
0.944444444444 -0.141414141414 0 2.0 1e-06 
1.0 -0.141414141414 0 2.0 1e-06 
0.5 -0.10101010101 0 2.0 1e-06 
0.555555555556 -0.10101010101 0 2.0 1e-06 
0.611111111111 -0.10101010101 0 2.0 1e-06 
0.666666666667 -0.10101010101 0 2.0 1e-06 
0.722222222222 -0.10101010101 0 2.0 1e-06 
0.777777777778 -0.10101010101 0 2.0 1e-06 
0.833333333333 -0.10101010101 0 2.0 1e-06 
0.888888888889 -0.10101010101 0 2.0 1e-06 
0.944444444444 -0.10101010101 0 2.0 1e-06 
1.0 -0.10101010101 0 2.0 1e-06 
0.5 -0.0606060606061 0 2.0 1e-06 
0.555555555556 -0.0606060606061 0 2.0 1e-06 
0.611111111111 -0.0606060606061 0 2.0 1e-06 
0.666666666667 -0.0606060606061 0 2.0 1e-06 
0.722222222222 -0.0606060606061 0 2.0 1e-06 
0.777777777778 -0.0606060606061 0 2.0 1e-06 
0.833333333333 -0.0606060606061 0 2.0 1e-06 
0.888888888889 -0.0606060606061 0 2.0 1e-06 
0.944444444444 -0.0606060606061 0 2.0 1e-06 
1.0 -0.0606060606061 0 2.0 1e-06 
0.5 -0.020202020202 0 2.0 1e-06 
0.555555555556 -0.020202020202 0 2.0 1e-06 
0.611111111111 -0.020202020202 0 2.0 1e-06 
0.666666666667 -0.020202020202 0 2.0 1e-06 
0.722222222222 -0.020202020202 0 2.0 1e-06 
0.777777777778 -0.020202020202 0 2.0 1e-06 
0.833333333333 -0.020202020202 0 2.0 1e-06 
0.888888888889 -0.020202020202 0 2.0 1e-06 
0.944444444444 -0.020202020202 0 2.0 1e-06 
1.0 -0.020202020202 0 2.0 1e-06 
0.5 0.020202020202 0 2.0 1e-06 
0.555555555556 0.020202020202 0 2.0 1e-06 
0.611111111111 0.020202020202 0 2.0 1e-06 
0.666666666667 0.020202020202 0 2.0 1e-06 
0.722222222222 0.020202020202 0 2.0 1e-06 
0.777777777778 0.020202020202 0 2.0 1e-06 
0.833333333333 0.020202020202 0 2.0 1e-06 
0.888888888889 0.020202020202 0 2.0 1e-06 
0.944444444444 0.020202020202 0 2.0 1e-06 
1.0 0.020202020202 0 2.0 1e-06 
0.5 0.0606060606061 0 2.0 1e-06 
0.555555555556 0.0606060606061 0 2.0 1e-06 
0.611111111111 0.0606060606061 0 2.0 1e-06 
0.666666666667 0.0606060606061 0 2.0 1e-06 
0.722222222222 0.0606060606061 0 2.0 1e-06 
0.777777777778 0.0606060606061 0 2.0 1e-06 
0.833333333333 0.0606060606061 0 2.0 1e-06 
0.888888888889 0.0606060606061 0 2.0 1e-06 
0.944444444444 0.0606060606061 0 2.0 1e-06 
1.0 0.0606060606061 0 2.0 1e-06 
0.5 0.10101010101 0 2.0 1e-06 
0.555555555556 0.10101010101 0 2.0 1e-06 
0.611111111111 0.10101010101 0 2.0 1e-06 
0.666666666667 0.10101010101 0 2.0 1e-06 
0.722222222222 0.10101010101 0 2.0 1e-06 
0.777777777778 0.10101010101 0 2.0 1e-06 
0.833333333333 0.10101010101 0 2.0 1e-06 
0.888888888889 0.10101010101 0 2.0 1e-06 
0.944444444444 0.10101010101 0 2.0 1e-06 
1.0 0.10101010101 0 2.0 1e-06 
0.5 0.141414141414 0 2.0 1e-06 
0.555555555556 0.141414141414 0 2.0 1e-06 
0.611111111111 0.141414141414 0 2.0 1e-06 
0.666666666667 0.141414141414 0 2.0 1e-06 
0.722222222222 0.141414141414 0 2.0 1e-06 
0.777777777778 0.141414141414 0 2.0 1e-06 
0.833333333333 0.141414141414 0 2.0 1e-06 
0.888888888889 0.141414141414 0 2.0 1e-06 
0.944444444444 0.141414141414 0 2.0 1e-06 
1.0 0.141414141414 0 2.0 1e-06 
0.5 0.181818181818 0 2.0 1e-06 
0.555555555556 0.181818181818 0 2.0 1e-06 
0.611111111111 0.181818181818 0 2.0 1e-06 
0.666666666667 0.181818181818 0 2.0 1e-06 
0.722222222222 0.181818181818 0 2.0 1e-06 
0.777777777778 0.181818181818 0 2.0 1e-06 
0.833333333333 0.181818181818 0 2.0 1e-06 
0.888888888889 0.181818181818 0 2.0 1e-06 
0.944444444444 0.181818181818 0 2.0 1e-06 
1.0 0.181818181818 0 2.0 1e-06 
0.5 0.222222222222 0 2.0 1e-06 
0.555555555556 0.222222222222 0 2.0 1e-06 
0.611111111111 0.222222222222 0 2.0 1e-06 
0.666666666667 0.222222222222 0 2.0 1e-06 
0.722222222222 0.222222222222 0 2.0 1e-06 
0.777777777778 0.222222222222 0 2.0 1e-06 
0.833333333333 0.222222222222 0 2.0 1e-06 
0.888888888889 0.222222222222 0 2.0 1e-06 
0.944444444444 0.222222222222 0 2.0 1e-06 
1.0 0.222222222222 0 2.0 1e-06 
0.5 0.262626262626 0 2.0 1e-06 
0.555555555556 0.262626262626 0 2.0 1e-06 
0.611111111111 0.262626262626 0 2.0 1e-06 
0.666666666667 0.262626262626 0 2.0 1e-06 
0.722222222222 0.262626262626 0 2.0 1e-06 
0.777777777778 0.262626262626 0 2.0 1e-06 
0.833333333333 0.262626262626 0 2.0 1e-06 
0.888888888889 0.262626262626 0 2.0 1e-06 
0.944444444444 0.262626262626 0 2.0 1e-06 
1.0 0.262626262626 0 2.0 1e-06 
0.5 0.30303030303 0 2.0 1e-06 
0.555555555556 0.30303030303 0 2.0 1e-06 
0.611111111111 0.30303030303 0 2.0 1e-06 
0.666666666667 0.30303030303 0 2.0 1e-06 
0.722222222222 0.30303030303 0 2.0 1e-06 
0.777777777778 0.30303030303 0 2.0 1e-06 
0.833333333333 0.30303030303 0 2.0 1e-06 
0.888888888889 0.30303030303 0 2.0 1e-06 
0.944444444444 0.30303030303 0 2.0 1e-06 
1.0 0.30303030303 0 2.0 1e-06 
0.5 0.343434343434 0 2.0 1e-06 
0.555555555556 0.343434343434 0 2.0 1e-06 
0.611111111111 0.343434343434 0 2.0 1e-06 
0.666666666667 0.343434343434 0 2.0 1e-06 
0.722222222222 0.343434343434 0 2.0 1e-06 
0.777777777778 0.343434343434 0 2.0 1e-06 
0.833333333333 0.343434343434 0 2.0 1e-06 
0.888888888889 0.343434343434 0 2.0 1e-06 
0.944444444444 0.343434343434 0 2.0 1e-06 
1.0 0.343434343434 0 2.0 1e-06 
0.5 0.383838383838 0 2.0 1e-06 
0.555555555556 0.383838383838 0 2.0 1e-06 
0.611111111111 0.383838383838 0 2.0 1e-06 
0.666666666667 0.383838383838 0 2.0 1e-06 
0.722222222222 0.383838383838 0 2.0 1e-06 
0.777777777778 0.383838383838 0 2.0 1e-06 
0.833333333333 0.383838383838 0 2.0 1e-06 
0.888888888889 0.383838383838 0 2.0 1e-06 
0.944444444444 0.383838383838 0 2.0 1e-06 
1.0 0.383838383838 0 2.0 1e-06 
0.5 0.424242424242 0 2.0 1e-06 
0.555555555556 0.424242424242 0 2.0 1e-06 
0.611111111111 0.424242424242 0 2.0 1e-06 
0.666666666667 0.424242424242 0 2.0 1e-06 
0.722222222222 0.424242424242 0 2.0 1e-06 
0.777777777778 0.424242424242 0 2.0 1e-06 
0.833333333333 0.424242424242 0 2.0 1e-06 
0.888888888889 0.424242424242 0 2.0 1e-06 
0.944444444444 0.424242424242 0 2.0 1e-06 
1.0 0.424242424242 0 2.0 1e-06 
0.5 0.464646464646 0 2.0 1e-06 
0.555555555556 0.464646464646 0 2.0 1e-06 
0.611111111111 0.464646464646 0 2.0 1e-06 
0.666666666667 0.464646464646 0 2.0 1e-06 
0.722222222222 0.464646464646 0 2.0 1e-06 
0.777777777778 0.464646464646 0 2.0 1e-06 
0.833333333333 0.464646464646 0 2.0 1e-06 
0.888888888889 0.464646464646 0 2.0 1e-06 
0.944444444444 0.464646464646 0 2.0 1e-06 
1.0 0.464646464646 0 2.0 1e-06 
0.5 0.505050505051 0 2.0 1e-06 
0.555555555556 0.505050505051 0 2.0 1e-06 
0.611111111111 0.505050505051 0 2.0 1e-06 
0.666666666667 0.505050505051 0 2.0 1e-06 
0.722222222222 0.505050505051 0 2.0 1e-06 
0.777777777778 0.505050505051 0 2.0 1e-06 
0.833333333333 0.505050505051 0 2.0 1e-06 
0.888888888889 0.505050505051 0 2.0 1e-06 
0.944444444444 0.505050505051 0 2.0 1e-06 
1.0 0.505050505051 0 2.0 1e-06 
0.5 0.545454545455 0 2.0 1e-06 
0.555555555556 0.545454545455 0 2.0 1e-06 
0.611111111111 0.545454545455 0 2.0 1e-06 
0.666666666667 0.545454545455 0 2.0 1e-06 
0.722222222222 0.545454545455 0 2.0 1e-06 
0.777777777778 0.545454545455 0 2.0 1e-06 
0.833333333333 0.545454545455 0 2.0 1e-06 
0.888888888889 0.545454545455 0 2.0 1e-06 
0.944444444444 0.545454545455 0 2.0 1e-06 
1.0 0.545454545455 0 2.0 1e-06 
0.5 0.585858585859 0 2.0 1e-06 
0.555555555556 0.585858585859 0 2.0 1e-06 
0.611111111111 0.585858585859 0 2.0 1e-06 
0.666666666667 0.585858585859 0 2.0 1e-06 
0.722222222222 0.585858585859 0 2.0 1e-06 
0.777777777778 0.585858585859 0 2.0 1e-06 
0.833333333333 0.585858585859 0 2.0 1e-06 
0.888888888889 0.585858585859 0 2.0 1e-06 
0.944444444444 0.585858585859 0 2.0 1e-06 
1.0 0.585858585859 0 2.0 1e-06 
0.5 0.626262626263 0 2.0 1e-06 
0.555555555556 0.626262626263 0 2.0 1e-06 
0.611111111111 0.626262626263 0 2.0 1e-06 
0.666666666667 0.626262626263 0 2.0 1e-06 
0.722222222222 0.626262626263 0 2.0 1e-06 
0.777777777778 0.626262626263 0 2.0 1e-06 
0.833333333333 0.626262626263 0 2.0 1e-06 
0.888888888889 0.626262626263 0 2.0 1e-06 
0.944444444444 0.626262626263 0 2.0 1e-06 
1.0 0.626262626263 0 2.0 1e-06 
0.5 0.666666666667 0 2.0 1e-06 
0.555555555556 0.666666666667 0 2.0 1e-06 
0.611111111111 0.666666666667 0 2.0 1e-06 
0.666666666667 0.666666666667 0 2.0 1e-06 
0.722222222222 0.666666666667 0 2.0 1e-06 
0.777777777778 0.666666666667 0 2.0 1e-06 
0.833333333333 0.666666666667 0 2.0 1e-06 
0.888888888889 0.666666666667 0 2.0 1e-06 
0.944444444444 0.666666666667 0 2.0 1e-06 
1.0 0.666666666667 0 2.0 1e-06 
0.5 0.707070707071 0 2.0 1e-06 
0.555555555556 0.707070707071 0 2.0 1e-06 
0.611111111111 0.707070707071 0 2.0 1e-06 
0.666666666667 0.707070707071 0 2.0 1e-06 
0.722222222222 0.707070707071 0 2.0 1e-06 
0.777777777778 0.707070707071 0 2.0 1e-06 
0.833333333333 0.707070707071 0 2.0 1e-06 
0.888888888889 0.707070707071 0 2.0 1e-06 
0.944444444444 0.707070707071 0 2.0 1e-06 
1.0 0.707070707071 0 2.0 1e-06 
0.5 0.747474747475 0 2.0 1e-06 
0.555555555556 0.747474747475 0 2.0 1e-06 
0.611111111111 0.747474747475 0 2.0 1e-06 
0.666666666667 0.747474747475 0 2.0 1e-06 
0.722222222222 0.747474747475 0 2.0 1e-06 
0.777777777778 0.747474747475 0 2.0 1e-06 
0.833333333333 0.747474747475 0 2.0 1e-06 
0.888888888889 0.747474747475 0 2.0 1e-06 
0.944444444444 0.747474747475 0 2.0 1e-06 
1.0 0.747474747475 0 2.0 1e-06 
0.5 0.787878787879 0 2.0 1e-06 
0.555555555556 0.787878787879 0 2.0 1e-06 
0.611111111111 0.787878787879 0 2.0 1e-06 
0.666666666667 0.787878787879 0 2.0 1e-06 
0.722222222222 0.787878787879 0 2.0 1e-06 
0.777777777778 0.787878787879 0 2.0 1e-06 
0.833333333333 0.787878787879 0 2.0 1e-06 
0.888888888889 0.787878787879 0 2.0 1e-06 
0.944444444444 0.787878787879 0 2.0 1e-06 
1.0 0.787878787879 0 2.0 1e-06 
0.5 0.828282828283 0 2.0 1e-06 
0.555555555556 0.828282828283 0 2.0 1e-06 
0.611111111111 0.828282828283 0 2.0 1e-06 
0.666666666667 0.828282828283 0 2.0 1e-06 
0.722222222222 0.828282828283 0 2.0 1e-06 
0.777777777778 0.828282828283 0 2.0 1e-06 
0.833333333333 0.828282828283 0 2.0 1e-06 
0.888888888889 0.828282828283 0 2.0 1e-06 
0.944444444444 0.828282828283 0 2.0 1e-06 
1.0 0.828282828283 0 2.0 1e-06 
0.5 0.868686868687 0 2.0 1e-06 
0.555555555556 0.868686868687 0 2.0 1e-06 
0.611111111111 0.868686868687 0 2.0 1e-06 
0.666666666667 0.868686868687 0 2.0 1e-06 
0.722222222222 0.868686868687 0 2.0 1e-06 
0.777777777778 0.868686868687 0 2.0 1e-06 
0.833333333333 0.868686868687 0 2.0 1e-06 
0.888888888889 0.868686868687 0 2.0 1e-06 
0.944444444444 0.868686868687 0 2.0 1e-06 
1.0 0.868686868687 0 2.0 1e-06 
0.5 0.909090909091 0 2.0 1e-06 
0.555555555556 0.909090909091 0 2.0 1e-06 
0.611111111111 0.909090909091 0 2.0 1e-06 
0.666666666667 0.909090909091 0 2.0 1e-06 
0.722222222222 0.909090909091 0 2.0 1e-06 
0.777777777778 0.909090909091 0 2.0 1e-06 
0.833333333333 0.909090909091 0 2.0 1e-06 
0.888888888889 0.909090909091 0 2.0 1e-06 
0.944444444444 0.909090909091 0 2.0 1e-06 
1.0 0.909090909091 0 2.0 1e-06 
0.5 0.949494949495 0 2.0 1e-06 
0.555555555556 0.949494949495 0 2.0 1e-06 
0.611111111111 0.949494949495 0 2.0 1e-06 
0.666666666667 0.949494949495 0 2.0 1e-06 
0.722222222222 0.949494949495 0 2.0 1e-06 
0.777777777778 0.949494949495 0 2.0 1e-06 
0.833333333333 0.949494949495 0 2.0 1e-06 
0.888888888889 0.949494949495 0 2.0 1e-06 
0.944444444444 0.949494949495 0 2.0 1e-06 
1.0 0.949494949495 0 2.0 1e-06 
0.5 0.989898989899 0 2.0 1e-06 
0.555555555556 0.989898989899 0 2.0 1e-06 
0.611111111111 0.989898989899 0 2.0 1e-06 
0.666666666667 0.989898989899 0 2.0 1e-06 
0.722222222222 0.989898989899 0 2.0 1e-06 
0.777777777778 0.989898989899 0 2.0 1e-06 
0.833333333333 0.989898989899 0 2.0 1e-06 
0.888888888889 0.989898989899 0 2.0 1e-06 
0.944444444444 0.989898989899 0 2.0 1e-06 
1.0 0.989898989899 0 2.0 1e-06 
0.5 1.0303030303 0 2.0 1e-06 
0.555555555556 1.0303030303 0 2.0 1e-06 
0.611111111111 1.0303030303 0 2.0 1e-06 
0.666666666667 1.0303030303 0 2.0 1e-06 
0.722222222222 1.0303030303 0 2.0 1e-06 
0.777777777778 1.0303030303 0 2.0 1e-06 
0.833333333333 1.0303030303 0 2.0 1e-06 
0.888888888889 1.0303030303 0 2.0 1e-06 
0.944444444444 1.0303030303 0 2.0 1e-06 
1.0 1.0303030303 0 2.0 1e-06 
0.5 1.07070707071 0 2.0 1e-06 
0.555555555556 1.07070707071 0 2.0 1e-06 
0.611111111111 1.07070707071 0 2.0 1e-06 
0.666666666667 1.07070707071 0 2.0 1e-06 
0.722222222222 1.07070707071 0 2.0 1e-06 
0.777777777778 1.07070707071 0 2.0 1e-06 
0.833333333333 1.07070707071 0 2.0 1e-06 
0.888888888889 1.07070707071 0 2.0 1e-06 
0.944444444444 1.07070707071 0 2.0 1e-06 
1.0 1.07070707071 0 2.0 1e-06 
0.5 1.11111111111 0 2.0 1e-06 
0.555555555556 1.11111111111 0 2.0 1e-06 
0.611111111111 1.11111111111 0 2.0 1e-06 
0.666666666667 1.11111111111 0 2.0 1e-06 
0.722222222222 1.11111111111 0 2.0 1e-06 
0.777777777778 1.11111111111 0 2.0 1e-06 
0.833333333333 1.11111111111 0 2.0 1e-06 
0.888888888889 1.11111111111 0 2.0 1e-06 
0.944444444444 1.11111111111 0 2.0 1e-06 
1.0 1.11111111111 0 2.0 1e-06 
0.5 1.15151515152 0 2.0 1e-06 
0.555555555556 1.15151515152 0 2.0 1e-06 
0.611111111111 1.15151515152 0 2.0 1e-06 
0.666666666667 1.15151515152 0 2.0 1e-06 
0.722222222222 1.15151515152 0 2.0 1e-06 
0.777777777778 1.15151515152 0 2.0 1e-06 
0.833333333333 1.15151515152 0 2.0 1e-06 
0.888888888889 1.15151515152 0 2.0 1e-06 
0.944444444444 1.15151515152 0 2.0 1e-06 
1.0 1.15151515152 0 2.0 1e-06 
0.5 1.19191919192 0 2.0 1e-06 
0.555555555556 1.19191919192 0 2.0 1e-06 
0.611111111111 1.19191919192 0 2.0 1e-06 
0.666666666667 1.19191919192 0 2.0 1e-06 
0.722222222222 1.19191919192 0 2.0 1e-06 
0.777777777778 1.19191919192 0 2.0 1e-06 
0.833333333333 1.19191919192 0 2.0 1e-06 
0.888888888889 1.19191919192 0 2.0 1e-06 
0.944444444444 1.19191919192 0 2.0 1e-06 
1.0 1.19191919192 0 2.0 1e-06 
0.5 1.23232323232 0 2.0 1e-06 
0.555555555556 1.23232323232 0 2.0 1e-06 
0.611111111111 1.23232323232 0 2.0 1e-06 
0.666666666667 1.23232323232 0 2.0 1e-06 
0.722222222222 1.23232323232 0 2.0 1e-06 
0.777777777778 1.23232323232 0 2.0 1e-06 
0.833333333333 1.23232323232 0 2.0 1e-06 
0.888888888889 1.23232323232 0 2.0 1e-06 
0.944444444444 1.23232323232 0 2.0 1e-06 
1.0 1.23232323232 0 2.0 1e-06 
0.5 1.27272727273 0 2.0 1e-06 
0.555555555556 1.27272727273 0 2.0 1e-06 
0.611111111111 1.27272727273 0 2.0 1e-06 
0.666666666667 1.27272727273 0 2.0 1e-06 
0.722222222222 1.27272727273 0 2.0 1e-06 
0.777777777778 1.27272727273 0 2.0 1e-06 
0.833333333333 1.27272727273 0 2.0 1e-06 
0.888888888889 1.27272727273 0 2.0 1e-06 
0.944444444444 1.27272727273 0 2.0 1e-06 
1.0 1.27272727273 0 2.0 1e-06 
0.5 1.31313131313 0 2.0 1e-06 
0.555555555556 1.31313131313 0 2.0 1e-06 
0.611111111111 1.31313131313 0 2.0 1e-06 
0.666666666667 1.31313131313 0 2.0 1e-06 
0.722222222222 1.31313131313 0 2.0 1e-06 
0.777777777778 1.31313131313 0 2.0 1e-06 
0.833333333333 1.31313131313 0 2.0 1e-06 
0.888888888889 1.31313131313 0 2.0 1e-06 
0.944444444444 1.31313131313 0 2.0 1e-06 
1.0 1.31313131313 0 2.0 1e-06 
0.5 1.35353535354 0 2.0 1e-06 
0.555555555556 1.35353535354 0 2.0 1e-06 
0.611111111111 1.35353535354 0 2.0 1e-06 
0.666666666667 1.35353535354 0 2.0 1e-06 
0.722222222222 1.35353535354 0 2.0 1e-06 
0.777777777778 1.35353535354 0 2.0 1e-06 
0.833333333333 1.35353535354 0 2.0 1e-06 
0.888888888889 1.35353535354 0 2.0 1e-06 
0.944444444444 1.35353535354 0 2.0 1e-06 
1.0 1.35353535354 0 2.0 1e-06 
0.5 1.39393939394 0 2.0 1e-06 
0.555555555556 1.39393939394 0 2.0 1e-06 
0.611111111111 1.39393939394 0 2.0 1e-06 
0.666666666667 1.39393939394 0 2.0 1e-06 
0.722222222222 1.39393939394 0 2.0 1e-06 
0.777777777778 1.39393939394 0 2.0 1e-06 
0.833333333333 1.39393939394 0 2.0 1e-06 
0.888888888889 1.39393939394 0 2.0 1e-06 
0.944444444444 1.39393939394 0 2.0 1e-06 
1.0 1.39393939394 0 2.0 1e-06 
0.5 1.43434343434 0 2.0 1e-06 
0.555555555556 1.43434343434 0 2.0 1e-06 
0.611111111111 1.43434343434 0 2.0 1e-06 
0.666666666667 1.43434343434 0 2.0 1e-06 
0.722222222222 1.43434343434 0 2.0 1e-06 
0.777777777778 1.43434343434 0 2.0 1e-06 
0.833333333333 1.43434343434 0 2.0 1e-06 
0.888888888889 1.43434343434 0 2.0 1e-06 
0.944444444444 1.43434343434 0 2.0 1e-06 
1.0 1.43434343434 0 2.0 1e-06 
0.5 1.47474747475 0 2.0 1e-06 
0.555555555556 1.47474747475 0 2.0 1e-06 
0.611111111111 1.47474747475 0 2.0 1e-06 
0.666666666667 1.47474747475 0 2.0 1e-06 
0.722222222222 1.47474747475 0 2.0 1e-06 
0.777777777778 1.47474747475 0 2.0 1e-06 
0.833333333333 1.47474747475 0 2.0 1e-06 
0.888888888889 1.47474747475 0 2.0 1e-06 
0.944444444444 1.47474747475 0 2.0 1e-06 
1.0 1.47474747475 0 2.0 1e-06 
0.5 1.51515151515 0 2.0 1e-06 
0.555555555556 1.51515151515 0 2.0 1e-06 
0.611111111111 1.51515151515 0 2.0 1e-06 
0.666666666667 1.51515151515 0 2.0 1e-06 
0.722222222222 1.51515151515 0 2.0 1e-06 
0.777777777778 1.51515151515 0 2.0 1e-06 
0.833333333333 1.51515151515 0 2.0 1e-06 
0.888888888889 1.51515151515 0 2.0 1e-06 
0.944444444444 1.51515151515 0 2.0 1e-06 
1.0 1.51515151515 0 2.0 1e-06 
0.5 1.55555555556 0 2.0 1e-06 
0.555555555556 1.55555555556 0 2.0 1e-06 
0.611111111111 1.55555555556 0 2.0 1e-06 
0.666666666667 1.55555555556 0 2.0 1e-06 
0.722222222222 1.55555555556 0 2.0 1e-06 
0.777777777778 1.55555555556 0 2.0 1e-06 
0.833333333333 1.55555555556 0 2.0 1e-06 
0.888888888889 1.55555555556 0 2.0 1e-06 
0.944444444444 1.55555555556 0 2.0 1e-06 
1.0 1.55555555556 0 2.0 1e-06 
0.5 1.59595959596 0 2.0 1e-06 
0.555555555556 1.59595959596 0 2.0 1e-06 
0.611111111111 1.59595959596 0 2.0 1e-06 
0.666666666667 1.59595959596 0 2.0 1e-06 
0.722222222222 1.59595959596 0 2.0 1e-06 
0.777777777778 1.59595959596 0 2.0 1e-06 
0.833333333333 1.59595959596 0 2.0 1e-06 
0.888888888889 1.59595959596 0 2.0 1e-06 
0.944444444444 1.59595959596 0 2.0 1e-06 
1.0 1.59595959596 0 2.0 1e-06 
0.5 1.63636363636 0 2.0 1e-06 
0.555555555556 1.63636363636 0 2.0 1e-06 
0.611111111111 1.63636363636 0 2.0 1e-06 
0.666666666667 1.63636363636 0 2.0 1e-06 
0.722222222222 1.63636363636 0 2.0 1e-06 
0.777777777778 1.63636363636 0 2.0 1e-06 
0.833333333333 1.63636363636 0 2.0 1e-06 
0.888888888889 1.63636363636 0 2.0 1e-06 
0.944444444444 1.63636363636 0 2.0 1e-06 
1.0 1.63636363636 0 2.0 1e-06 
0.5 1.67676767677 0 2.0 1e-06 
0.555555555556 1.67676767677 0 2.0 1e-06 
0.611111111111 1.67676767677 0 2.0 1e-06 
0.666666666667 1.67676767677 0 2.0 1e-06 
0.722222222222 1.67676767677 0 2.0 1e-06 
0.777777777778 1.67676767677 0 2.0 1e-06 
0.833333333333 1.67676767677 0 2.0 1e-06 
0.888888888889 1.67676767677 0 2.0 1e-06 
0.944444444444 1.67676767677 0 2.0 1e-06 
1.0 1.67676767677 0 2.0 1e-06 
0.5 1.71717171717 0 2.0 1e-06 
0.555555555556 1.71717171717 0 2.0 1e-06 
0.611111111111 1.71717171717 0 2.0 1e-06 
0.666666666667 1.71717171717 0 2.0 1e-06 
0.722222222222 1.71717171717 0 2.0 1e-06 
0.777777777778 1.71717171717 0 2.0 1e-06 
0.833333333333 1.71717171717 0 2.0 1e-06 
0.888888888889 1.71717171717 0 2.0 1e-06 
0.944444444444 1.71717171717 0 2.0 1e-06 
1.0 1.71717171717 0 2.0 1e-06 
0.5 1.75757575758 0 2.0 1e-06 
0.555555555556 1.75757575758 0 2.0 1e-06 
0.611111111111 1.75757575758 0 2.0 1e-06 
0.666666666667 1.75757575758 0 2.0 1e-06 
0.722222222222 1.75757575758 0 2.0 1e-06 
0.777777777778 1.75757575758 0 2.0 1e-06 
0.833333333333 1.75757575758 0 2.0 1e-06 
0.888888888889 1.75757575758 0 2.0 1e-06 
0.944444444444 1.75757575758 0 2.0 1e-06 
1.0 1.75757575758 0 2.0 1e-06 
0.5 1.79797979798 0 2.0 1e-06 
0.555555555556 1.79797979798 0 2.0 1e-06 
0.611111111111 1.79797979798 0 2.0 1e-06 
0.666666666667 1.79797979798 0 2.0 1e-06 
0.722222222222 1.79797979798 0 2.0 1e-06 
0.777777777778 1.79797979798 0 2.0 1e-06 
0.833333333333 1.79797979798 0 2.0 1e-06 
0.888888888889 1.79797979798 0 2.0 1e-06 
0.944444444444 1.79797979798 0 2.0 1e-06 
1.0 1.79797979798 0 2.0 1e-06 
0.5 1.83838383838 0 2.0 1e-06 
0.555555555556 1.83838383838 0 2.0 1e-06 
0.611111111111 1.83838383838 0 2.0 1e-06 
0.666666666667 1.83838383838 0 2.0 1e-06 
0.722222222222 1.83838383838 0 2.0 1e-06 
0.777777777778 1.83838383838 0 2.0 1e-06 
0.833333333333 1.83838383838 0 2.0 1e-06 
0.888888888889 1.83838383838 0 2.0 1e-06 
0.944444444444 1.83838383838 0 2.0 1e-06 
1.0 1.83838383838 0 2.0 1e-06 
0.5 1.87878787879 0 2.0 1e-06 
0.555555555556 1.87878787879 0 2.0 1e-06 
0.611111111111 1.87878787879 0 2.0 1e-06 
0.666666666667 1.87878787879 0 2.0 1e-06 
0.722222222222 1.87878787879 0 2.0 1e-06 
0.777777777778 1.87878787879 0 2.0 1e-06 
0.833333333333 1.87878787879 0 2.0 1e-06 
0.888888888889 1.87878787879 0 2.0 1e-06 
0.944444444444 1.87878787879 0 2.0 1e-06 
1.0 1.87878787879 0 2.0 1e-06 
0.5 1.91919191919 0 2.0 1e-06 
0.555555555556 1.91919191919 0 2.0 1e-06 
0.611111111111 1.91919191919 0 2.0 1e-06 
0.666666666667 1.91919191919 0 2.0 1e-06 
0.722222222222 1.91919191919 0 2.0 1e-06 
0.777777777778 1.91919191919 0 2.0 1e-06 
0.833333333333 1.91919191919 0 2.0 1e-06 
0.888888888889 1.91919191919 0 2.0 1e-06 
0.944444444444 1.91919191919 0 2.0 1e-06 
1.0 1.91919191919 0 2.0 1e-06 
0.5 1.9595959596 0 2.0 1e-06 
0.555555555556 1.9595959596 0 2.0 1e-06 
0.611111111111 1.9595959596 0 2.0 1e-06 
0.666666666667 1.9595959596 0 2.0 1e-06 
0.722222222222 1.9595959596 0 2.0 1e-06 
0.777777777778 1.9595959596 0 2.0 1e-06 
0.833333333333 1.9595959596 0 2.0 1e-06 
0.888888888889 1.9595959596 0 2.0 1e-06 
0.944444444444 1.9595959596 0 2.0 1e-06 
1.0 1.9595959596 0 2.0 1e-06 
0.5 2.0 0 2.0 1e-06 
0.555555555556 2.0 0 2.0 1e-06 
0.611111111111 2.0 0 2.0 1e-06 
0.666666666667 2.0 0 2.0 1e-06 
0.722222222222 2.0 0 2.0 1e-06 
0.777777777778 2.0 0 2.0 1e-06 
0.833333333333 2.0 0 2.0 1e-06 
0.888888888889 2.0 0 2.0 1e-06 
0.944444444444 2.0 0 2.0 1e-06 
1.0 2.0 0 2.0 1e-06 
.ENDDATA 
.dc sweep DATA = datadc 
.print dc X1:IDS X1:QFG 
.end