*script to generate hspice simulation using cmdp, Juan Duarte 
*Date: 07/21/2015, time: 07:55:49

.option abstol=1e-6 reltol=1e-6 post ingold 
.option measform=1 
.temp 27 

.hdl "/users/jpduarte/research/BSIMCMG/workingcode/bsimcmg.va" 
.include "/users/jpduarte/research/userjp/ncfet/modelcards/modelcard.nmos" 

.PARAM Vd_value = 0 
.PARAM Vg_value = 0 
.PARAM Vs_value = 0 
.PARAM Vb_value = 0 
.PARAM L_value = 1e-06 

Vd Vd 0.0 dc = Vd_value 
Vg Vg 0.0 dc = Vg_value 
Vs Vs 0.0 dc = Vs_value 
Vb Vb 0.0 dc = Vb_value 

X1 Vd Vg Vs Vb nmos1 L = 'L_value'

.DATA datadc Vd_value Vg_value Vs_value Vb_value L_value 
0.05 0.0 0 0 1e-06 
0.3 0.0 0 0 1e-06 
0.05 0.0030303030303 0 0 1e-06 
0.3 0.0030303030303 0 0 1e-06 
0.05 0.00606060606061 0 0 1e-06 
0.3 0.00606060606061 0 0 1e-06 
0.05 0.00909090909091 0 0 1e-06 
0.3 0.00909090909091 0 0 1e-06 
0.05 0.0121212121212 0 0 1e-06 
0.3 0.0121212121212 0 0 1e-06 
0.05 0.0151515151515 0 0 1e-06 
0.3 0.0151515151515 0 0 1e-06 
0.05 0.0181818181818 0 0 1e-06 
0.3 0.0181818181818 0 0 1e-06 
0.05 0.0212121212121 0 0 1e-06 
0.3 0.0212121212121 0 0 1e-06 
0.05 0.0242424242424 0 0 1e-06 
0.3 0.0242424242424 0 0 1e-06 
0.05 0.0272727272727 0 0 1e-06 
0.3 0.0272727272727 0 0 1e-06 
0.05 0.030303030303 0 0 1e-06 
0.3 0.030303030303 0 0 1e-06 
0.05 0.0333333333333 0 0 1e-06 
0.3 0.0333333333333 0 0 1e-06 
0.05 0.0363636363636 0 0 1e-06 
0.3 0.0363636363636 0 0 1e-06 
0.05 0.0393939393939 0 0 1e-06 
0.3 0.0393939393939 0 0 1e-06 
0.05 0.0424242424242 0 0 1e-06 
0.3 0.0424242424242 0 0 1e-06 
0.05 0.0454545454545 0 0 1e-06 
0.3 0.0454545454545 0 0 1e-06 
0.05 0.0484848484848 0 0 1e-06 
0.3 0.0484848484848 0 0 1e-06 
0.05 0.0515151515152 0 0 1e-06 
0.3 0.0515151515152 0 0 1e-06 
0.05 0.0545454545455 0 0 1e-06 
0.3 0.0545454545455 0 0 1e-06 
0.05 0.0575757575758 0 0 1e-06 
0.3 0.0575757575758 0 0 1e-06 
0.05 0.0606060606061 0 0 1e-06 
0.3 0.0606060606061 0 0 1e-06 
0.05 0.0636363636364 0 0 1e-06 
0.3 0.0636363636364 0 0 1e-06 
0.05 0.0666666666667 0 0 1e-06 
0.3 0.0666666666667 0 0 1e-06 
0.05 0.069696969697 0 0 1e-06 
0.3 0.069696969697 0 0 1e-06 
0.05 0.0727272727273 0 0 1e-06 
0.3 0.0727272727273 0 0 1e-06 
0.05 0.0757575757576 0 0 1e-06 
0.3 0.0757575757576 0 0 1e-06 
0.05 0.0787878787879 0 0 1e-06 
0.3 0.0787878787879 0 0 1e-06 
0.05 0.0818181818182 0 0 1e-06 
0.3 0.0818181818182 0 0 1e-06 
0.05 0.0848484848485 0 0 1e-06 
0.3 0.0848484848485 0 0 1e-06 
0.05 0.0878787878788 0 0 1e-06 
0.3 0.0878787878788 0 0 1e-06 
0.05 0.0909090909091 0 0 1e-06 
0.3 0.0909090909091 0 0 1e-06 
0.05 0.0939393939394 0 0 1e-06 
0.3 0.0939393939394 0 0 1e-06 
0.05 0.0969696969697 0 0 1e-06 
0.3 0.0969696969697 0 0 1e-06 
0.05 0.1 0 0 1e-06 
0.3 0.1 0 0 1e-06 
0.05 0.10303030303 0 0 1e-06 
0.3 0.10303030303 0 0 1e-06 
0.05 0.106060606061 0 0 1e-06 
0.3 0.106060606061 0 0 1e-06 
0.05 0.109090909091 0 0 1e-06 
0.3 0.109090909091 0 0 1e-06 
0.05 0.112121212121 0 0 1e-06 
0.3 0.112121212121 0 0 1e-06 
0.05 0.115151515152 0 0 1e-06 
0.3 0.115151515152 0 0 1e-06 
0.05 0.118181818182 0 0 1e-06 
0.3 0.118181818182 0 0 1e-06 
0.05 0.121212121212 0 0 1e-06 
0.3 0.121212121212 0 0 1e-06 
0.05 0.124242424242 0 0 1e-06 
0.3 0.124242424242 0 0 1e-06 
0.05 0.127272727273 0 0 1e-06 
0.3 0.127272727273 0 0 1e-06 
0.05 0.130303030303 0 0 1e-06 
0.3 0.130303030303 0 0 1e-06 
0.05 0.133333333333 0 0 1e-06 
0.3 0.133333333333 0 0 1e-06 
0.05 0.136363636364 0 0 1e-06 
0.3 0.136363636364 0 0 1e-06 
0.05 0.139393939394 0 0 1e-06 
0.3 0.139393939394 0 0 1e-06 
0.05 0.142424242424 0 0 1e-06 
0.3 0.142424242424 0 0 1e-06 
0.05 0.145454545455 0 0 1e-06 
0.3 0.145454545455 0 0 1e-06 
0.05 0.148484848485 0 0 1e-06 
0.3 0.148484848485 0 0 1e-06 
0.05 0.151515151515 0 0 1e-06 
0.3 0.151515151515 0 0 1e-06 
0.05 0.154545454545 0 0 1e-06 
0.3 0.154545454545 0 0 1e-06 
0.05 0.157575757576 0 0 1e-06 
0.3 0.157575757576 0 0 1e-06 
0.05 0.160606060606 0 0 1e-06 
0.3 0.160606060606 0 0 1e-06 
0.05 0.163636363636 0 0 1e-06 
0.3 0.163636363636 0 0 1e-06 
0.05 0.166666666667 0 0 1e-06 
0.3 0.166666666667 0 0 1e-06 
0.05 0.169696969697 0 0 1e-06 
0.3 0.169696969697 0 0 1e-06 
0.05 0.172727272727 0 0 1e-06 
0.3 0.172727272727 0 0 1e-06 
0.05 0.175757575758 0 0 1e-06 
0.3 0.175757575758 0 0 1e-06 
0.05 0.178787878788 0 0 1e-06 
0.3 0.178787878788 0 0 1e-06 
0.05 0.181818181818 0 0 1e-06 
0.3 0.181818181818 0 0 1e-06 
0.05 0.184848484848 0 0 1e-06 
0.3 0.184848484848 0 0 1e-06 
0.05 0.187878787879 0 0 1e-06 
0.3 0.187878787879 0 0 1e-06 
0.05 0.190909090909 0 0 1e-06 
0.3 0.190909090909 0 0 1e-06 
0.05 0.193939393939 0 0 1e-06 
0.3 0.193939393939 0 0 1e-06 
0.05 0.19696969697 0 0 1e-06 
0.3 0.19696969697 0 0 1e-06 
0.05 0.2 0 0 1e-06 
0.3 0.2 0 0 1e-06 
0.05 0.20303030303 0 0 1e-06 
0.3 0.20303030303 0 0 1e-06 
0.05 0.206060606061 0 0 1e-06 
0.3 0.206060606061 0 0 1e-06 
0.05 0.209090909091 0 0 1e-06 
0.3 0.209090909091 0 0 1e-06 
0.05 0.212121212121 0 0 1e-06 
0.3 0.212121212121 0 0 1e-06 
0.05 0.215151515152 0 0 1e-06 
0.3 0.215151515152 0 0 1e-06 
0.05 0.218181818182 0 0 1e-06 
0.3 0.218181818182 0 0 1e-06 
0.05 0.221212121212 0 0 1e-06 
0.3 0.221212121212 0 0 1e-06 
0.05 0.224242424242 0 0 1e-06 
0.3 0.224242424242 0 0 1e-06 
0.05 0.227272727273 0 0 1e-06 
0.3 0.227272727273 0 0 1e-06 
0.05 0.230303030303 0 0 1e-06 
0.3 0.230303030303 0 0 1e-06 
0.05 0.233333333333 0 0 1e-06 
0.3 0.233333333333 0 0 1e-06 
0.05 0.236363636364 0 0 1e-06 
0.3 0.236363636364 0 0 1e-06 
0.05 0.239393939394 0 0 1e-06 
0.3 0.239393939394 0 0 1e-06 
0.05 0.242424242424 0 0 1e-06 
0.3 0.242424242424 0 0 1e-06 
0.05 0.245454545455 0 0 1e-06 
0.3 0.245454545455 0 0 1e-06 
0.05 0.248484848485 0 0 1e-06 
0.3 0.248484848485 0 0 1e-06 
0.05 0.251515151515 0 0 1e-06 
0.3 0.251515151515 0 0 1e-06 
0.05 0.254545454545 0 0 1e-06 
0.3 0.254545454545 0 0 1e-06 
0.05 0.257575757576 0 0 1e-06 
0.3 0.257575757576 0 0 1e-06 
0.05 0.260606060606 0 0 1e-06 
0.3 0.260606060606 0 0 1e-06 
0.05 0.263636363636 0 0 1e-06 
0.3 0.263636363636 0 0 1e-06 
0.05 0.266666666667 0 0 1e-06 
0.3 0.266666666667 0 0 1e-06 
0.05 0.269696969697 0 0 1e-06 
0.3 0.269696969697 0 0 1e-06 
0.05 0.272727272727 0 0 1e-06 
0.3 0.272727272727 0 0 1e-06 
0.05 0.275757575758 0 0 1e-06 
0.3 0.275757575758 0 0 1e-06 
0.05 0.278787878788 0 0 1e-06 
0.3 0.278787878788 0 0 1e-06 
0.05 0.281818181818 0 0 1e-06 
0.3 0.281818181818 0 0 1e-06 
0.05 0.284848484848 0 0 1e-06 
0.3 0.284848484848 0 0 1e-06 
0.05 0.287878787879 0 0 1e-06 
0.3 0.287878787879 0 0 1e-06 
0.05 0.290909090909 0 0 1e-06 
0.3 0.290909090909 0 0 1e-06 
0.05 0.293939393939 0 0 1e-06 
0.3 0.293939393939 0 0 1e-06 
0.05 0.29696969697 0 0 1e-06 
0.3 0.29696969697 0 0 1e-06 
0.05 0.3 0 0 1e-06 
0.3 0.3 0 0 1e-06 
.ENDDATA 
.dc sweep DATA = datadc 
.print dc X1:Ids X1:Qg X1:E_FE X1:V_FE 
.end