*script to generate hspice simulation using cmdp, Juan Duarte 
*Date: 04/25/2015, time: 13:59:53

.option abstol=1e-6 reltol=1e-6 post ingold 
.option measform=1 
.temp 27 

.hdl "/users/jpduarte/BSIM_CM_Matlab/BSIM_model_development_v2/DM_Verilog_Hspice/Models_Verilog/BSIMIMGref/code/bsimimg.va" 
.include "/users/jpduarte/BSIM_CM_Matlab/BSIM_model_development_v2/DM_Verilog_Hspice/Models_Verilog/BSIMIMG/benchmark_tests/modelcard.nmos" 

.PARAM Vd_value = 0 
.PARAM Vgf_value = 0 
.PARAM Vs_value = 0 
.PARAM Vgb_value = 0 
.PARAM L_value = 5e-08 

Vd Vd 0.0 dc = Vd_value 
Vgf Vgf 0.0 dc = Vgf_value 
Vs Vs 0.0 dc = Vs_value 
Vgb Vgb 0.0 dc = Vgb_value 

X1 Vd Vgf Vs Vgb nmos1 L = 'L_value'

.DATA datadc Vd_value Vgf_value Vs_value Vgb_value L_value 
0.05 0.0 0 0 5e-08 
0.145 0.0 0 0 5e-08 
0.24 0.0 0 0 5e-08 
0.335 0.0 0 0 5e-08 
0.43 0.0 0 0 5e-08 
0.525 0.0 0 0 5e-08 
0.62 0.0 0 0 5e-08 
0.715 0.0 0 0 5e-08 
0.81 0.0 0 0 5e-08 
0.905 0.0 0 0 5e-08 
1.0 0.0 0 0 5e-08 
0.05 0.0344827586207 0 0 5e-08 
0.145 0.0344827586207 0 0 5e-08 
0.24 0.0344827586207 0 0 5e-08 
0.335 0.0344827586207 0 0 5e-08 
0.43 0.0344827586207 0 0 5e-08 
0.525 0.0344827586207 0 0 5e-08 
0.62 0.0344827586207 0 0 5e-08 
0.715 0.0344827586207 0 0 5e-08 
0.81 0.0344827586207 0 0 5e-08 
0.905 0.0344827586207 0 0 5e-08 
1.0 0.0344827586207 0 0 5e-08 
0.05 0.0689655172414 0 0 5e-08 
0.145 0.0689655172414 0 0 5e-08 
0.24 0.0689655172414 0 0 5e-08 
0.335 0.0689655172414 0 0 5e-08 
0.43 0.0689655172414 0 0 5e-08 
0.525 0.0689655172414 0 0 5e-08 
0.62 0.0689655172414 0 0 5e-08 
0.715 0.0689655172414 0 0 5e-08 
0.81 0.0689655172414 0 0 5e-08 
0.905 0.0689655172414 0 0 5e-08 
1.0 0.0689655172414 0 0 5e-08 
0.05 0.103448275862 0 0 5e-08 
0.145 0.103448275862 0 0 5e-08 
0.24 0.103448275862 0 0 5e-08 
0.335 0.103448275862 0 0 5e-08 
0.43 0.103448275862 0 0 5e-08 
0.525 0.103448275862 0 0 5e-08 
0.62 0.103448275862 0 0 5e-08 
0.715 0.103448275862 0 0 5e-08 
0.81 0.103448275862 0 0 5e-08 
0.905 0.103448275862 0 0 5e-08 
1.0 0.103448275862 0 0 5e-08 
0.05 0.137931034483 0 0 5e-08 
0.145 0.137931034483 0 0 5e-08 
0.24 0.137931034483 0 0 5e-08 
0.335 0.137931034483 0 0 5e-08 
0.43 0.137931034483 0 0 5e-08 
0.525 0.137931034483 0 0 5e-08 
0.62 0.137931034483 0 0 5e-08 
0.715 0.137931034483 0 0 5e-08 
0.81 0.137931034483 0 0 5e-08 
0.905 0.137931034483 0 0 5e-08 
1.0 0.137931034483 0 0 5e-08 
0.05 0.172413793103 0 0 5e-08 
0.145 0.172413793103 0 0 5e-08 
0.24 0.172413793103 0 0 5e-08 
0.335 0.172413793103 0 0 5e-08 
0.43 0.172413793103 0 0 5e-08 
0.525 0.172413793103 0 0 5e-08 
0.62 0.172413793103 0 0 5e-08 
0.715 0.172413793103 0 0 5e-08 
0.81 0.172413793103 0 0 5e-08 
0.905 0.172413793103 0 0 5e-08 
1.0 0.172413793103 0 0 5e-08 
0.05 0.206896551724 0 0 5e-08 
0.145 0.206896551724 0 0 5e-08 
0.24 0.206896551724 0 0 5e-08 
0.335 0.206896551724 0 0 5e-08 
0.43 0.206896551724 0 0 5e-08 
0.525 0.206896551724 0 0 5e-08 
0.62 0.206896551724 0 0 5e-08 
0.715 0.206896551724 0 0 5e-08 
0.81 0.206896551724 0 0 5e-08 
0.905 0.206896551724 0 0 5e-08 
1.0 0.206896551724 0 0 5e-08 
0.05 0.241379310345 0 0 5e-08 
0.145 0.241379310345 0 0 5e-08 
0.24 0.241379310345 0 0 5e-08 
0.335 0.241379310345 0 0 5e-08 
0.43 0.241379310345 0 0 5e-08 
0.525 0.241379310345 0 0 5e-08 
0.62 0.241379310345 0 0 5e-08 
0.715 0.241379310345 0 0 5e-08 
0.81 0.241379310345 0 0 5e-08 
0.905 0.241379310345 0 0 5e-08 
1.0 0.241379310345 0 0 5e-08 
0.05 0.275862068966 0 0 5e-08 
0.145 0.275862068966 0 0 5e-08 
0.24 0.275862068966 0 0 5e-08 
0.335 0.275862068966 0 0 5e-08 
0.43 0.275862068966 0 0 5e-08 
0.525 0.275862068966 0 0 5e-08 
0.62 0.275862068966 0 0 5e-08 
0.715 0.275862068966 0 0 5e-08 
0.81 0.275862068966 0 0 5e-08 
0.905 0.275862068966 0 0 5e-08 
1.0 0.275862068966 0 0 5e-08 
0.05 0.310344827586 0 0 5e-08 
0.145 0.310344827586 0 0 5e-08 
0.24 0.310344827586 0 0 5e-08 
0.335 0.310344827586 0 0 5e-08 
0.43 0.310344827586 0 0 5e-08 
0.525 0.310344827586 0 0 5e-08 
0.62 0.310344827586 0 0 5e-08 
0.715 0.310344827586 0 0 5e-08 
0.81 0.310344827586 0 0 5e-08 
0.905 0.310344827586 0 0 5e-08 
1.0 0.310344827586 0 0 5e-08 
0.05 0.344827586207 0 0 5e-08 
0.145 0.344827586207 0 0 5e-08 
0.24 0.344827586207 0 0 5e-08 
0.335 0.344827586207 0 0 5e-08 
0.43 0.344827586207 0 0 5e-08 
0.525 0.344827586207 0 0 5e-08 
0.62 0.344827586207 0 0 5e-08 
0.715 0.344827586207 0 0 5e-08 
0.81 0.344827586207 0 0 5e-08 
0.905 0.344827586207 0 0 5e-08 
1.0 0.344827586207 0 0 5e-08 
0.05 0.379310344828 0 0 5e-08 
0.145 0.379310344828 0 0 5e-08 
0.24 0.379310344828 0 0 5e-08 
0.335 0.379310344828 0 0 5e-08 
0.43 0.379310344828 0 0 5e-08 
0.525 0.379310344828 0 0 5e-08 
0.62 0.379310344828 0 0 5e-08 
0.715 0.379310344828 0 0 5e-08 
0.81 0.379310344828 0 0 5e-08 
0.905 0.379310344828 0 0 5e-08 
1.0 0.379310344828 0 0 5e-08 
0.05 0.413793103448 0 0 5e-08 
0.145 0.413793103448 0 0 5e-08 
0.24 0.413793103448 0 0 5e-08 
0.335 0.413793103448 0 0 5e-08 
0.43 0.413793103448 0 0 5e-08 
0.525 0.413793103448 0 0 5e-08 
0.62 0.413793103448 0 0 5e-08 
0.715 0.413793103448 0 0 5e-08 
0.81 0.413793103448 0 0 5e-08 
0.905 0.413793103448 0 0 5e-08 
1.0 0.413793103448 0 0 5e-08 
0.05 0.448275862069 0 0 5e-08 
0.145 0.448275862069 0 0 5e-08 
0.24 0.448275862069 0 0 5e-08 
0.335 0.448275862069 0 0 5e-08 
0.43 0.448275862069 0 0 5e-08 
0.525 0.448275862069 0 0 5e-08 
0.62 0.448275862069 0 0 5e-08 
0.715 0.448275862069 0 0 5e-08 
0.81 0.448275862069 0 0 5e-08 
0.905 0.448275862069 0 0 5e-08 
1.0 0.448275862069 0 0 5e-08 
0.05 0.48275862069 0 0 5e-08 
0.145 0.48275862069 0 0 5e-08 
0.24 0.48275862069 0 0 5e-08 
0.335 0.48275862069 0 0 5e-08 
0.43 0.48275862069 0 0 5e-08 
0.525 0.48275862069 0 0 5e-08 
0.62 0.48275862069 0 0 5e-08 
0.715 0.48275862069 0 0 5e-08 
0.81 0.48275862069 0 0 5e-08 
0.905 0.48275862069 0 0 5e-08 
1.0 0.48275862069 0 0 5e-08 
0.05 0.51724137931 0 0 5e-08 
0.145 0.51724137931 0 0 5e-08 
0.24 0.51724137931 0 0 5e-08 
0.335 0.51724137931 0 0 5e-08 
0.43 0.51724137931 0 0 5e-08 
0.525 0.51724137931 0 0 5e-08 
0.62 0.51724137931 0 0 5e-08 
0.715 0.51724137931 0 0 5e-08 
0.81 0.51724137931 0 0 5e-08 
0.905 0.51724137931 0 0 5e-08 
1.0 0.51724137931 0 0 5e-08 
0.05 0.551724137931 0 0 5e-08 
0.145 0.551724137931 0 0 5e-08 
0.24 0.551724137931 0 0 5e-08 
0.335 0.551724137931 0 0 5e-08 
0.43 0.551724137931 0 0 5e-08 
0.525 0.551724137931 0 0 5e-08 
0.62 0.551724137931 0 0 5e-08 
0.715 0.551724137931 0 0 5e-08 
0.81 0.551724137931 0 0 5e-08 
0.905 0.551724137931 0 0 5e-08 
1.0 0.551724137931 0 0 5e-08 
0.05 0.586206896552 0 0 5e-08 
0.145 0.586206896552 0 0 5e-08 
0.24 0.586206896552 0 0 5e-08 
0.335 0.586206896552 0 0 5e-08 
0.43 0.586206896552 0 0 5e-08 
0.525 0.586206896552 0 0 5e-08 
0.62 0.586206896552 0 0 5e-08 
0.715 0.586206896552 0 0 5e-08 
0.81 0.586206896552 0 0 5e-08 
0.905 0.586206896552 0 0 5e-08 
1.0 0.586206896552 0 0 5e-08 
0.05 0.620689655172 0 0 5e-08 
0.145 0.620689655172 0 0 5e-08 
0.24 0.620689655172 0 0 5e-08 
0.335 0.620689655172 0 0 5e-08 
0.43 0.620689655172 0 0 5e-08 
0.525 0.620689655172 0 0 5e-08 
0.62 0.620689655172 0 0 5e-08 
0.715 0.620689655172 0 0 5e-08 
0.81 0.620689655172 0 0 5e-08 
0.905 0.620689655172 0 0 5e-08 
1.0 0.620689655172 0 0 5e-08 
0.05 0.655172413793 0 0 5e-08 
0.145 0.655172413793 0 0 5e-08 
0.24 0.655172413793 0 0 5e-08 
0.335 0.655172413793 0 0 5e-08 
0.43 0.655172413793 0 0 5e-08 
0.525 0.655172413793 0 0 5e-08 
0.62 0.655172413793 0 0 5e-08 
0.715 0.655172413793 0 0 5e-08 
0.81 0.655172413793 0 0 5e-08 
0.905 0.655172413793 0 0 5e-08 
1.0 0.655172413793 0 0 5e-08 
0.05 0.689655172414 0 0 5e-08 
0.145 0.689655172414 0 0 5e-08 
0.24 0.689655172414 0 0 5e-08 
0.335 0.689655172414 0 0 5e-08 
0.43 0.689655172414 0 0 5e-08 
0.525 0.689655172414 0 0 5e-08 
0.62 0.689655172414 0 0 5e-08 
0.715 0.689655172414 0 0 5e-08 
0.81 0.689655172414 0 0 5e-08 
0.905 0.689655172414 0 0 5e-08 
1.0 0.689655172414 0 0 5e-08 
0.05 0.724137931034 0 0 5e-08 
0.145 0.724137931034 0 0 5e-08 
0.24 0.724137931034 0 0 5e-08 
0.335 0.724137931034 0 0 5e-08 
0.43 0.724137931034 0 0 5e-08 
0.525 0.724137931034 0 0 5e-08 
0.62 0.724137931034 0 0 5e-08 
0.715 0.724137931034 0 0 5e-08 
0.81 0.724137931034 0 0 5e-08 
0.905 0.724137931034 0 0 5e-08 
1.0 0.724137931034 0 0 5e-08 
0.05 0.758620689655 0 0 5e-08 
0.145 0.758620689655 0 0 5e-08 
0.24 0.758620689655 0 0 5e-08 
0.335 0.758620689655 0 0 5e-08 
0.43 0.758620689655 0 0 5e-08 
0.525 0.758620689655 0 0 5e-08 
0.62 0.758620689655 0 0 5e-08 
0.715 0.758620689655 0 0 5e-08 
0.81 0.758620689655 0 0 5e-08 
0.905 0.758620689655 0 0 5e-08 
1.0 0.758620689655 0 0 5e-08 
0.05 0.793103448276 0 0 5e-08 
0.145 0.793103448276 0 0 5e-08 
0.24 0.793103448276 0 0 5e-08 
0.335 0.793103448276 0 0 5e-08 
0.43 0.793103448276 0 0 5e-08 
0.525 0.793103448276 0 0 5e-08 
0.62 0.793103448276 0 0 5e-08 
0.715 0.793103448276 0 0 5e-08 
0.81 0.793103448276 0 0 5e-08 
0.905 0.793103448276 0 0 5e-08 
1.0 0.793103448276 0 0 5e-08 
0.05 0.827586206897 0 0 5e-08 
0.145 0.827586206897 0 0 5e-08 
0.24 0.827586206897 0 0 5e-08 
0.335 0.827586206897 0 0 5e-08 
0.43 0.827586206897 0 0 5e-08 
0.525 0.827586206897 0 0 5e-08 
0.62 0.827586206897 0 0 5e-08 
0.715 0.827586206897 0 0 5e-08 
0.81 0.827586206897 0 0 5e-08 
0.905 0.827586206897 0 0 5e-08 
1.0 0.827586206897 0 0 5e-08 
0.05 0.862068965517 0 0 5e-08 
0.145 0.862068965517 0 0 5e-08 
0.24 0.862068965517 0 0 5e-08 
0.335 0.862068965517 0 0 5e-08 
0.43 0.862068965517 0 0 5e-08 
0.525 0.862068965517 0 0 5e-08 
0.62 0.862068965517 0 0 5e-08 
0.715 0.862068965517 0 0 5e-08 
0.81 0.862068965517 0 0 5e-08 
0.905 0.862068965517 0 0 5e-08 
1.0 0.862068965517 0 0 5e-08 
0.05 0.896551724138 0 0 5e-08 
0.145 0.896551724138 0 0 5e-08 
0.24 0.896551724138 0 0 5e-08 
0.335 0.896551724138 0 0 5e-08 
0.43 0.896551724138 0 0 5e-08 
0.525 0.896551724138 0 0 5e-08 
0.62 0.896551724138 0 0 5e-08 
0.715 0.896551724138 0 0 5e-08 
0.81 0.896551724138 0 0 5e-08 
0.905 0.896551724138 0 0 5e-08 
1.0 0.896551724138 0 0 5e-08 
0.05 0.931034482759 0 0 5e-08 
0.145 0.931034482759 0 0 5e-08 
0.24 0.931034482759 0 0 5e-08 
0.335 0.931034482759 0 0 5e-08 
0.43 0.931034482759 0 0 5e-08 
0.525 0.931034482759 0 0 5e-08 
0.62 0.931034482759 0 0 5e-08 
0.715 0.931034482759 0 0 5e-08 
0.81 0.931034482759 0 0 5e-08 
0.905 0.931034482759 0 0 5e-08 
1.0 0.931034482759 0 0 5e-08 
0.05 0.965517241379 0 0 5e-08 
0.145 0.965517241379 0 0 5e-08 
0.24 0.965517241379 0 0 5e-08 
0.335 0.965517241379 0 0 5e-08 
0.43 0.965517241379 0 0 5e-08 
0.525 0.965517241379 0 0 5e-08 
0.62 0.965517241379 0 0 5e-08 
0.715 0.965517241379 0 0 5e-08 
0.81 0.965517241379 0 0 5e-08 
0.905 0.965517241379 0 0 5e-08 
1.0 0.965517241379 0 0 5e-08 
0.05 1.0 0 0 5e-08 
0.145 1.0 0 0 5e-08 
0.24 1.0 0 0 5e-08 
0.335 1.0 0 0 5e-08 
0.43 1.0 0 0 5e-08 
0.525 1.0 0 0 5e-08 
0.62 1.0 0 0 5e-08 
0.715 1.0 0 0 5e-08 
0.81 1.0 0 0 5e-08 
0.905 1.0 0 0 5e-08 
1.0 1.0 0 0 5e-08 
.ENDDATA 
.dc sweep DATA = datadc 
.print dc X1:IDS X1:CDFGI X1:CDSI X1:vbgs 
.end